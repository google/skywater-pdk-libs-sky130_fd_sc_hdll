* File: sky130_fd_sc_hdll__nor3_4.pex.spice
* Created: Thu Aug 27 19:16:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR3_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 38 39
r72 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r73 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=1.75 $Y=1.202
+ $X2=1.925 $Y2=1.202
r74 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.75
+ $Y=1.16 $X2=1.75 $Y2=1.16
r75 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.75 $Y2=1.202
r76 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r77 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.43 $Y2=1.202
r78 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r79 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=0.58 $Y=1.202
+ $X2=0.96 $Y2=1.202
r80 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.16 $X2=0.58 $Y2=1.16
r81 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.58 $Y2=1.202
r82 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r83 25 38 55.7186 $w=2.08e-07 $l=1.055e-06 $layer=LI1_cond $X=0.695 $Y=1.18
+ $X2=1.75 $Y2=1.18
r84 25 31 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=0.695 $Y=1.18
+ $X2=0.58 $Y2=1.18
r85 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r86 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r87 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r88 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r89 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r90 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r91 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r92 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r93 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r94 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r95 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r96 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=0.56
r97 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r98 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r99 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r100 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 26 27 28 30 31 35 38 47 53
r126 47 48 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=3.335 $Y=1.202
+ $X2=3.36 $Y2=1.202
r127 46 47 60.5722 $w=3.74e-07 $l=4.7e-07 $layer=POLY_cond $X=2.865 $Y=1.202
+ $X2=3.335 $Y2=1.202
r128 45 53 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.85 $Y=1.18
+ $X2=2.965 $Y2=1.18
r129 44 46 1.93316 $w=3.74e-07 $l=1.5e-08 $layer=POLY_cond $X=2.85 $Y=1.202
+ $X2=2.865 $Y2=1.202
r130 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.85
+ $Y=1.16 $X2=2.85 $Y2=1.16
r131 42 44 1.28877 $w=3.74e-07 $l=1e-08 $layer=POLY_cond $X=2.84 $Y=1.202
+ $X2=2.85 $Y2=1.202
r132 41 42 57.3503 $w=3.74e-07 $l=4.45e-07 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.84 $Y2=1.202
r133 40 41 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=2.37 $Y=1.202
+ $X2=2.395 $Y2=1.202
r134 38 53 1.05628 $w=2.08e-07 $l=2e-08 $layer=LI1_cond $X=2.985 $Y=1.18
+ $X2=2.965 $Y2=1.18
r135 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.71
+ $Y=1.16 $X2=5.71 $Y2=1.16
r136 32 35 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=5.63 $Y=1.18 $X2=5.71
+ $Y2=1.18
r137 31 38 49.1169 $w=2.08e-07 $l=9.3e-07 $layer=LI1_cond $X=3.915 $Y=1.18
+ $X2=2.985 $Y2=1.18
r138 29 32 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.63 $Y=1.285
+ $X2=5.63 $Y2=1.18
r139 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.63 $Y=1.285
+ $X2=5.63 $Y2=1.445
r140 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.545 $Y=1.53
+ $X2=5.63 $Y2=1.445
r141 27 28 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=5.545 $Y=1.53
+ $X2=4.085 $Y2=1.53
r142 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4 $Y=1.445
+ $X2=4.085 $Y2=1.53
r143 25 31 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=4 $Y=1.285
+ $X2=3.915 $Y2=1.18
r144 25 26 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4 $Y=1.285 $X2=4
+ $Y2=1.445
r145 22 36 38.7084 $w=3.43e-07 $l=1.77059e-07 $layer=POLY_cond $X=5.71 $Y=0.995
+ $X2=5.735 $Y2=1.16
r146 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.71 $Y=0.995
+ $X2=5.71 $Y2=0.56
r147 19 36 45.964 $w=3.43e-07 $l=2.73861e-07 $layer=POLY_cond $X=5.685 $Y=1.41
+ $X2=5.735 $Y2=1.16
r148 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.685 $Y=1.41
+ $X2=5.685 $Y2=1.985
r149 16 48 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=1.202
r150 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=0.56
r151 13 47 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.202
r152 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.985
r153 10 46 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.202
r154 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.985
r155 7 42 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=1.202
r156 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=0.56
r157 4 41 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.202
r158 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r159 1 40 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=1.202
r160 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_4%C 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 35 36
r89 36 37 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.215 $Y=1.202
+ $X2=5.24 $Y2=1.202
r90 34 36 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=5.04 $Y=1.202
+ $X2=5.215 $Y2=1.202
r91 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.04
+ $Y=1.16 $X2=5.04 $Y2=1.16
r92 32 34 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=4.745 $Y=1.202
+ $X2=5.04 $Y2=1.202
r93 31 32 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.72 $Y=1.202
+ $X2=4.745 $Y2=1.202
r94 30 31 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.275 $Y=1.202
+ $X2=4.72 $Y2=1.202
r95 29 30 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.25 $Y=1.202
+ $X2=4.275 $Y2=1.202
r96 28 29 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=3.805 $Y=1.202
+ $X2=4.25 $Y2=1.202
r97 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.78 $Y=1.202
+ $X2=3.805 $Y2=1.202
r98 25 35 0.345283 $w=1.058e-06 $l=3e-08 $layer=LI1_cond $X=4.785 $Y=1.19
+ $X2=4.785 $Y2=1.16
r99 22 37 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=1.202
r100 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=0.56
r101 19 36 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.202
r102 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.985
r103 16 32 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.202
r104 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.985
r105 13 31 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.72 $Y=0.995
+ $X2=4.72 $Y2=1.202
r106 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.72 $Y=0.995
+ $X2=4.72 $Y2=0.56
r107 10 30 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.202
r108 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.985
r109 7 29 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.25 $Y=0.995
+ $X2=4.25 $Y2=1.202
r110 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.25 $Y=0.995
+ $X2=4.25 $Y2=0.56
r111 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.202
r112 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.985
r113 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.78 $Y=0.995
+ $X2=3.78 $Y2=1.202
r114 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.78 $Y=0.995
+ $X2=3.78 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 32 37 43 52 54 55 56
r92 54 56 0.140654 $w=2.7e-07 $l=1.95e-07 $layer=MET1_cond $X=5.89 $Y=2.2
+ $X2=5.695 $Y2=2.2
r93 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.89 $Y=2.21
+ $X2=5.89 $Y2=2.21
r94 52 56 3.36014 $w=1.4e-07 $l=2.715e-06 $layer=MET1_cond $X=2.98 $Y=2.21
+ $X2=5.695 $Y2=2.21
r95 49 52 0.143387 $w=2.7e-07 $l=2e-07 $layer=MET1_cond $X=2.78 $Y=2.2 $X2=2.98
+ $Y2=2.2
r96 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.78 $Y=2.21
+ $X2=2.78 $Y2=2.21
r97 43 50 5.91385 $w=3.78e-07 $l=1.95e-07 $layer=LI1_cond $X=2.975 $Y=2.275
+ $X2=2.78 $Y2=2.275
r98 43 45 2.85751 $w=3.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.975 $Y=2.275
+ $X2=3.1 $Y2=2.275
r99 40 50 15.0121 $w=3.78e-07 $l=4.95e-07 $layer=LI1_cond $X=2.285 $Y=2.275
+ $X2=2.78 $Y2=2.275
r100 40 42 2.85751 $w=3.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=2.275
+ $X2=2.16 $Y2=2.275
r101 30 45 4.34342 $w=2.5e-07 $l=1.9e-07 $layer=LI1_cond $X=3.1 $Y=2.085 $X2=3.1
+ $Y2=2.275
r102 30 32 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.1 $Y=2.085
+ $X2=3.1 $Y2=1.96
r103 29 42 4.34342 $w=2.5e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=2.085
+ $X2=2.16 $Y2=2.275
r104 28 39 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=1.625
+ $X2=2.16 $Y2=1.54
r105 28 29 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.16 $Y=1.625
+ $X2=2.16 $Y2=2.085
r106 27 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=1.54
+ $X2=1.22 $Y2=1.54
r107 26 39 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=2.16 $Y2=1.54
r108 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=1.345 $Y2=1.54
r109 22 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=1.54
r110 22 24 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=2.3
r111 21 35 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.277 $Y2=1.54
r112 20 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=1.22 $Y2=1.54
r113 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=0.405 $Y2=1.54
r114 16 35 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=1.54
r115 16 18 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=2.3
r116 5 55 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.775
+ $Y=1.485 $X2=5.92 $Y2=2.3
r117 4 45 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=2.3
r118 4 32 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=1.96
r119 3 42 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.3
r120 3 39 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.62
r121 2 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r122 2 24 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r123 1 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r124 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_4%VPWR 1 2 11 13 17 19 26 27 30 33 36
r80 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r81 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r82 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r83 26 27 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r84 24 27 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=2.07 $Y=2.72 $X2=6.21
+ $Y2=2.72
r85 24 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r86 23 26 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=6.21 $Y2=2.72
r87 23 24 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r88 21 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.69 $Y2=2.72
r89 21 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=2.07 $Y2=2.72
r90 19 31 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r91 19 36 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r92 15 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=2.72
r93 15 17 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=1.96
r94 14 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r95 13 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=1.69 $Y2=2.72
r96 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=0.875 $Y2=2.72
r97 9 30 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r98 9 11 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r99 2 17 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.96
r100 1 11 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_4%A_497_297# 1 2 3 4 15 17 18 19 21 24 30 35
r66 35 37 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=5.45 $Y=2.3 $X2=5.45
+ $Y2=2.38
r67 30 32 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.51 $Y=2.3 $X2=4.51
+ $Y2=2.38
r68 22 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.635 $Y=2.38
+ $X2=4.51 $Y2=2.38
r69 21 37 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.325 $Y=2.38
+ $X2=5.45 $Y2=2.38
r70 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.325 $Y=2.38
+ $X2=4.635 $Y2=2.38
r71 20 28 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.695 $Y=2.38
+ $X2=3.57 $Y2=2.38
r72 19 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.385 $Y=2.38
+ $X2=4.51 $Y2=2.38
r73 19 20 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.385 $Y=2.38
+ $X2=3.695 $Y2=2.38
r74 18 28 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=2.295
+ $X2=3.57 $Y2=2.38
r75 17 26 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=1.625
+ $X2=3.57 $Y2=1.54
r76 17 18 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.57 $Y=1.625
+ $X2=3.57 $Y2=2.295
r77 16 24 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=1.54
+ $X2=2.63 $Y2=1.54
r78 15 26 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.445 $Y=1.54
+ $X2=3.57 $Y2=1.54
r79 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.445 $Y=1.54
+ $X2=2.755 $Y2=1.54
r80 4 35 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.305
+ $Y=1.485 $X2=5.45 $Y2=2.3
r81 3 30 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.365
+ $Y=1.485 $X2=4.51 $Y2=2.3
r82 2 28 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=2.3
r83 2 26 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=1.62
r84 1 24 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_4%Y 1 2 3 4 5 6 7 8 27 29 30 33 35 39 41 45
+ 47 49 53 55 57 61 63 65 66 67 68 73 74 80 83
r182 82 83 10.1336 $w=2.88e-07 $l=2.55e-07 $layer=LI1_cond $X=6.2 $Y=1.785
+ $X2=6.2 $Y2=1.53
r183 81 83 24.8371 $w=2.88e-07 $l=6.25e-07 $layer=LI1_cond $X=6.2 $Y=0.905
+ $X2=6.2 $Y2=1.53
r184 76 78 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=1.875
+ $X2=4.98 $Y2=1.96
r185 74 76 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.98 $Y=1.87
+ $X2=4.98 $Y2=1.875
r186 68 71 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=1.875
+ $X2=4.04 $Y2=1.96
r187 64 80 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.615 $Y=0.815
+ $X2=5.425 $Y2=0.815
r188 63 81 7.31368 $w=1.8e-07 $l=1.84594e-07 $layer=LI1_cond $X=6.055 $Y=0.815
+ $X2=6.2 $Y2=0.905
r189 63 64 27.1111 $w=1.78e-07 $l=4.4e-07 $layer=LI1_cond $X=6.055 $Y=0.815
+ $X2=5.615 $Y2=0.815
r190 59 80 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.425 $Y=0.725
+ $X2=5.425 $Y2=0.815
r191 59 61 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.425 $Y=0.725
+ $X2=5.425 $Y2=0.39
r192 58 74 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.105 $Y=1.87
+ $X2=4.98 $Y2=1.87
r193 57 82 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=6.055 $Y=1.87
+ $X2=6.2 $Y2=1.785
r194 57 58 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=6.055 $Y=1.87
+ $X2=5.105 $Y2=1.87
r195 56 73 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.675 $Y=0.815
+ $X2=4.485 $Y2=0.815
r196 55 80 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.235 $Y=0.815
+ $X2=5.425 $Y2=0.815
r197 55 56 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.235 $Y=0.815
+ $X2=4.675 $Y2=0.815
r198 51 73 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.485 $Y=0.725
+ $X2=4.485 $Y2=0.815
r199 51 53 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.485 $Y=0.725
+ $X2=4.485 $Y2=0.39
r200 50 68 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.165 $Y=1.875
+ $X2=4.04 $Y2=1.875
r201 49 76 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=1.875
+ $X2=4.98 $Y2=1.875
r202 49 50 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=4.855 $Y=1.875
+ $X2=4.165 $Y2=1.875
r203 48 67 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.735 $Y=0.815
+ $X2=3.545 $Y2=0.815
r204 47 73 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.295 $Y=0.815
+ $X2=4.485 $Y2=0.815
r205 47 48 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.295 $Y=0.815
+ $X2=3.735 $Y2=0.815
r206 43 67 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.545 $Y2=0.815
r207 43 45 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.545 $Y2=0.39
r208 42 66 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.795 $Y=0.815
+ $X2=2.605 $Y2=0.815
r209 41 67 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=3.545 $Y2=0.815
r210 41 42 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=2.795 $Y2=0.815
r211 37 66 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.605 $Y2=0.815
r212 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.605 $Y2=0.39
r213 36 65 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=0.815
+ $X2=1.665 $Y2=0.815
r214 35 66 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=2.605 $Y2=0.815
r215 35 36 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=1.855 $Y2=0.815
r216 31 65 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.815
r217 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.39
r218 29 65 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=1.665 $Y2=0.815
r219 29 30 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=0.915 $Y2=0.815
r220 25 30 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.815
r221 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r222 8 78 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=4.835
+ $Y=1.485 $X2=4.98 $Y2=1.96
r223 7 71 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.485 $X2=4.04 $Y2=1.96
r224 6 61 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.315
+ $Y=0.235 $X2=5.45 $Y2=0.39
r225 5 53 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.325
+ $Y=0.235 $X2=4.51 $Y2=0.39
r226 4 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.435
+ $Y=0.235 $X2=3.57 $Y2=0.39
r227 3 39 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.235 $X2=2.63 $Y2=0.39
r228 2 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r229 1 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_4%VGND 1 2 3 4 5 6 7 22 24 26 30 34 38 42 46
+ 50 53 54 56 57 59 60 62 63 65 66 67 86 87 93
r114 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r115 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r116 84 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r117 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r118 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r119 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r120 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r121 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r122 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r123 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r124 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r125 72 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r126 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r127 69 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r128 69 71 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=2.07 $Y2=0
r129 67 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r130 67 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r131 65 83 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.75
+ $Y2=0
r132 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.92
+ $Y2=0
r133 64 86 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.005 $Y=0
+ $X2=6.21 $Y2=0
r134 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0 $X2=5.92
+ $Y2=0
r135 62 80 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.83
+ $Y2=0
r136 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.98
+ $Y2=0
r137 61 83 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.065 $Y=0
+ $X2=5.75 $Y2=0
r138 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=4.98
+ $Y2=0
r139 59 77 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.955 $Y=0 $X2=3.91
+ $Y2=0
r140 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0 $X2=4.04
+ $Y2=0
r141 58 80 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.125 $Y=0
+ $X2=4.83 $Y2=0
r142 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0 $X2=4.04
+ $Y2=0
r143 56 74 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=2.99
+ $Y2=0
r144 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.1
+ $Y2=0
r145 55 77 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=3.91 $Y2=0
r146 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.1
+ $Y2=0
r147 53 71 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r148 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.16
+ $Y2=0
r149 52 74 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.99 $Y2=0
r150 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r151 48 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r152 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.39
r153 44 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r154 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.39
r155 40 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r156 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.39
r157 36 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0
r158 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0.39
r159 32 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r160 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.39
r161 28 93 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r162 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r163 27 90 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r164 26 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r165 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=0.365 $Y2=0
r166 22 90 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r167 22 24 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r168 7 50 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.785
+ $Y=0.235 $X2=5.92 $Y2=0.39
r169 6 46 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.795
+ $Y=0.235 $X2=4.98 $Y2=0.39
r170 5 42 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.235 $X2=4.04 $Y2=0.39
r171 4 38 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.39
r172 3 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r173 2 30 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
r174 1 24 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

