* File: sky130_fd_sc_hdll__and3b_1.pex.spice
* Created: Thu Aug 27 18:58:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND3B_1%A_N 2 3 5 8 9 10 11 16 18
r25 16 19 77.9987 $w=4.85e-07 $l=5.35e-07 $layer=POLY_cond $X=0.352 $Y=1.16
+ $X2=0.352 $Y2=1.695
r26 16 18 46.1122 $w=4.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.352 $Y=1.16
+ $X2=0.352 $Y2=0.995
r27 10 11 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.255 $Y=1.53
+ $X2=0.255 $Y2=1.87
r28 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.16
+ $X2=0.255 $Y2=1.53
r29 9 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.26 $Y=1.16
+ $X2=0.26 $Y2=1.16
r30 8 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.52 $Y=0.675
+ $X2=0.52 $Y2=0.995
r31 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r32 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r33 2 19 64.6575 $w=2e-07 $l=1.95e-07 $layer=POLY_cond $X=0.495 $Y=1.89
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_1%A_117_413# 1 2 7 9 12 14 16 20
c41 20 0 2.08002e-19 $X=1.35 $Y=1.16
r42 24 25 14.4424 $w=3.21e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0.74
+ $X2=0.705 $Y2=1.12
r43 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.35
+ $Y=1.16 $X2=1.35 $Y2=1.16
r44 18 25 2.20369 $w=2.5e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.12
+ $X2=0.705 $Y2=1.12
r45 18 20 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=0.895 $Y=1.12
+ $X2=1.35 $Y2=1.12
r46 14 25 7.43575 $w=3.21e-07 $l=1.36931e-07 $layer=LI1_cond $X=0.73 $Y=1.245
+ $X2=0.705 $Y2=1.12
r47 14 16 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=0.73 $Y=1.245
+ $X2=0.73 $Y2=2.26
r48 10 21 38.5363 $w=3.15e-07 $l=2.13014e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.4 $Y2=1.16
r49 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.475
r50 7 21 57.7442 $w=3.15e-07 $l=3.6e-07 $layer=POLY_cond $X=1.485 $Y=1.48
+ $X2=1.4 $Y2=1.16
r51 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.485 $Y=1.48
+ $X2=1.485 $Y2=1.765
r52 2 16 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.26
r53 1 24 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.465 $X2=0.73 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_1%B 1 2 4 7 10 18
c39 7 0 1.69741e-19 $X=1.98 $Y=0.475
c40 1 0 3.82617e-20 $X=1.955 $Y=1.48
r41 14 18 3.22006 $w=3.38e-07 $l=9.5e-08 $layer=LI1_cond $X=2.005 $Y=2.295
+ $X2=2.1 $Y2=2.295
r42 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.005
+ $Y=2.3 $X2=2.005 $Y2=2.3
r43 10 18 5.08431 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=2.25 $Y=2.295
+ $X2=2.1 $Y2=2.295
r44 7 9 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=1.98 $Y=0.475
+ $X2=1.98 $Y2=1.2
r45 2 13 38.4563 $w=3.24e-07 $l=2.26031e-07 $layer=POLY_cond $X=1.955 $Y=2.105
+ $X2=2.022 $Y2=2.3
r46 2 4 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.955 $Y=2.105
+ $X2=1.955 $Y2=1.765
r47 1 9 110.989 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=1.955 $Y=1.48
+ $X2=1.955 $Y2=1.2
r48 1 4 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.955 $Y=1.48
+ $X2=1.955 $Y2=1.765
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_1%C 3 5 7 8 9
c32 3 0 5.85457e-20 $X=2.385 $Y=0.475
r33 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.445
+ $Y=1.16 $X2=2.445 $Y2=1.16
r34 9 14 9.78787 $w=3.63e-07 $l=3.1e-07 $layer=LI1_cond $X=2.462 $Y=0.85
+ $X2=2.462 $Y2=1.16
r35 8 9 10.7351 $w=3.63e-07 $l=3.4e-07 $layer=LI1_cond $X=2.462 $Y=0.51
+ $X2=2.462 $Y2=0.85
r36 5 13 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.48 $Y=1.41
+ $X2=2.445 $Y2=1.16
r37 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.48 $Y=1.41 $X2=2.48
+ $Y2=1.695
r38 1 13 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.385 $Y=0.995
+ $X2=2.445 $Y2=1.16
r39 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.385 $Y=0.995
+ $X2=2.385 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_1%A_225_311# 1 2 3 10 12 13 15 18 20 24 25
+ 27 30 31 34 37 40
c81 34 0 5.85457e-20 $X=3.1 $Y=1.16
r82 39 40 7.25089 $w=4.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=1.657
+ $X2=2.155 $Y2=1.657
r83 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=1.16 $X2=3.1 $Y2=1.16
r84 32 34 13.8817 $w=2.18e-07 $l=2.65e-07 $layer=LI1_cond $X=3.075 $Y=1.425
+ $X2=3.075 $Y2=1.16
r85 31 39 3.78115 $w=4.63e-07 $l=1.47e-07 $layer=LI1_cond $X=2.387 $Y=1.657
+ $X2=2.24 $Y2=1.657
r86 30 32 6.49156 $w=4.22e-07 $l=2.81681e-07 $layer=LI1_cond $X=2.965 $Y=1.657
+ $X2=3.075 $Y2=1.425
r87 30 31 14.8674 $w=4.63e-07 $l=5.78e-07 $layer=LI1_cond $X=2.965 $Y=1.657
+ $X2=2.387 $Y2=1.657
r88 29 37 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.945 $Y=1.51
+ $X2=1.817 $Y2=1.51
r89 29 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.945 $Y=1.51
+ $X2=2.155 $Y2=1.51
r90 27 37 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.817 $Y=1.425
+ $X2=1.817 $Y2=1.51
r91 26 27 39.5446 $w=2.53e-07 $l=8.75e-07 $layer=LI1_cond $X=1.817 $Y=0.55
+ $X2=1.817 $Y2=1.425
r92 24 37 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.69 $Y=1.51
+ $X2=1.817 $Y2=1.51
r93 24 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.69 $Y=1.51
+ $X2=1.335 $Y2=1.51
r94 20 26 6.81977 $w=2.65e-07 $l=1.85957e-07 $layer=LI1_cond $X=1.69 $Y=0.417
+ $X2=1.817 $Y2=0.55
r95 20 22 18.0477 $w=2.63e-07 $l=4.15e-07 $layer=LI1_cond $X=1.69 $Y=0.417
+ $X2=1.275 $Y2=0.417
r96 16 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.21 $Y=1.595
+ $X2=1.335 $Y2=1.51
r97 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=1.595
+ $X2=1.21 $Y2=1.76
r98 13 35 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.16 $Y=0.995
+ $X2=3.1 $Y2=1.16
r99 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.16 $Y=0.995
+ $X2=3.16 $Y2=0.56
r100 10 35 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.135 $Y=1.41
+ $X2=3.1 $Y2=1.16
r101 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.135 $Y=1.41
+ $X2=3.135 $Y2=1.985
r102 3 39 600 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.555 $X2=2.24 $Y2=1.725
r103 2 18 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.555 $X2=1.25 $Y2=1.76
r104 1 22 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.15
+ $Y=0.265 $X2=1.275 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_1%VPWR 1 2 3 10 12 14 20 25 28 29 30 37 38
+ 44
r55 46 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r57 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 35 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r60 32 34 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.75 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 30 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 30 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 28 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.53 $Y2=2.72
r64 28 29 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.902 $Y2=2.72
r65 27 37 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.01 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 27 29 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=3.01 $Y=2.72
+ $X2=2.902 $Y2=2.72
r67 18 29 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.902 $Y=2.635
+ $X2=2.902 $Y2=2.72
r68 18 20 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=2.902 $Y=2.635
+ $X2=2.902 $Y2=2.34
r69 16 25 5.42871 $w=1.88e-07 $l=9.3e-08 $layer=LI1_cond $X=1.627 $Y=1.86
+ $X2=1.72 $Y2=1.86
r70 16 44 8.23174 $w=2.43e-07 $l=1.75e-07 $layer=LI1_cond $X=1.627 $Y=1.955
+ $X2=1.627 $Y2=2.13
r71 15 41 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r72 14 32 8.98481 $w=1.7e-07 $l=3.33e-07 $layer=LI1_cond $X=1.417 $Y=2.72
+ $X2=1.75 $Y2=2.72
r73 14 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r74 14 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 14 44 15.623 $w=6.63e-07 $l=5.9e-07 $layer=LI1_cond $X=1.417 $Y=2.72
+ $X2=1.417 $Y2=2.13
r76 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.085 $Y=2.72
+ $X2=0.345 $Y2=2.72
r77 10 41 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r78 10 12 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.29
r79 3 20 600 $w=1.7e-07 $l=1.00657e-06 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=1.485 $X2=2.9 $Y2=2.34
r80 2 25 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.555 $X2=1.72 $Y2=1.85
r81 1 12 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_1%X 1 2 9 10 12 13 14 22
r16 14 22 12.1768 $w=2.63e-07 $l=2.8e-07 $layer=LI1_cond $X=3.402 $Y=2.21
+ $X2=3.402 $Y2=1.93
r17 11 13 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=3.405 $Y=0.605
+ $X2=3.405 $Y2=0.51
r18 11 12 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.405 $Y=0.605
+ $X2=3.405 $Y2=0.735
r19 10 12 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.45 $Y=1.765
+ $X2=3.45 $Y2=0.735
r20 9 22 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=3.402 $Y=1.897
+ $X2=3.402 $Y2=1.93
r21 9 10 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=3.402 $Y=1.897
+ $X2=3.402 $Y2=1.765
r22 2 22 300 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_PDIFF $count=2 $X=3.225
+ $Y=1.485 $X2=3.37 $Y2=1.93
r23 1 13 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=3.235
+ $Y=0.235 $X2=3.37 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_1%VGND 1 2 7 9 13 15 17 27 28 34
r36 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r37 28 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r38 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r39 25 34 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=2.96
+ $Y2=0
r40 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.45
+ $Y2=0
r41 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r42 23 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r43 21 24 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r44 20 23 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r45 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r46 18 31 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r47 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r48 17 34 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.96
+ $Y2=0
r49 17 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.53
+ $Y2=0
r50 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r51 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r52 11 34 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.96 $Y=0.085
+ $X2=2.96 $Y2=0
r53 11 13 14.9023 $w=2.88e-07 $l=3.75e-07 $layer=LI1_cond $X=2.96 $Y=0.085
+ $X2=2.96 $Y2=0.46
r54 7 31 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r55 7 9 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.73
r56 2 13 182 $w=1.7e-07 $l=5.6921e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.265 $X2=2.94 $Y2=0.46
r57 1 9 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.73
.ends

