* File: sky130_fd_sc_hdll__clkinv_2.spice
* Created: Wed Sep  2 08:26:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkinv_2.pex.spice"
.subckt sky130_fd_sc_hdll__clkinv_2  VNB VPB A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.1323
+ AS=0.0693 PD=1.47 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.1092
+ AS=0.0693 PD=1.36 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.275
+ AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.1575
+ AS=0.15 PD=1.315 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1004 N_Y_M1002_d N_A_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1 AD=0.1575
+ AS=0.275 PD=1.315 PS=2.55 NRD=4.9053 NRS=1.9503 M=1 R=5.55556 SA=90001.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX5_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hdll__clkinv_2.pxi.spice"
*
.ends
*
*
