* File: sky130_fd_sc_hdll__isobufsrc_2.pxi.spice
* Created: Thu Aug 27 19:09:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%SLEEP N_SLEEP_c_65_n N_SLEEP_M1004_g
+ N_SLEEP_c_68_n N_SLEEP_M1000_g N_SLEEP_c_69_n N_SLEEP_M1007_g N_SLEEP_c_66_n
+ N_SLEEP_M1009_g SLEEP N_SLEEP_c_67_n SLEEP
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%SLEEP
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%A_271_21# N_A_271_21#_M1001_s
+ N_A_271_21#_M1006_s N_A_271_21#_c_101_n N_A_271_21#_M1005_g
+ N_A_271_21#_c_111_n N_A_271_21#_M1002_g N_A_271_21#_c_112_n
+ N_A_271_21#_M1003_g N_A_271_21#_c_102_n N_A_271_21#_M1008_g
+ N_A_271_21#_c_103_n N_A_271_21#_c_104_n N_A_271_21#_c_105_n
+ N_A_271_21#_c_106_n N_A_271_21#_c_107_n N_A_271_21#_c_108_n
+ N_A_271_21#_c_116_n N_A_271_21#_c_109_n N_A_271_21#_c_110_n
+ N_A_271_21#_c_117_n PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%A_271_21#
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%A N_A_M1001_g N_A_c_186_n N_A_c_187_n
+ N_A_M1006_g A A A N_A_c_184_n N_A_c_185_n A
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%A
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%A_27_297# N_A_27_297#_M1000_s
+ N_A_27_297#_M1007_s N_A_27_297#_M1003_d N_A_27_297#_c_217_n
+ N_A_27_297#_c_218_n N_A_27_297#_c_219_n N_A_27_297#_c_220_n
+ N_A_27_297#_c_243_p N_A_27_297#_c_229_n N_A_27_297#_c_221_n
+ N_A_27_297#_c_222_n N_A_27_297#_c_223_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%VPWR N_VPWR_M1000_d N_VPWR_M1006_d
+ N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_264_n N_VPWR_c_265_n VPWR
+ N_VPWR_c_266_n N_VPWR_c_261_n N_VPWR_c_268_n VPWR
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%VPWR
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%X N_X_M1004_d N_X_M1005_s N_X_M1002_s
+ N_X_c_306_n N_X_c_301_n N_X_c_302_n N_X_c_303_n N_X_c_304_n X N_X_c_315_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%X
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%VGND N_VGND_M1004_s N_VGND_M1009_s
+ N_VGND_M1008_d N_VGND_M1001_d N_VGND_c_347_n N_VGND_c_348_n N_VGND_c_349_n
+ N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n N_VGND_c_354_n
+ N_VGND_c_355_n N_VGND_c_356_n VGND N_VGND_c_357_n N_VGND_c_358_n
+ N_VGND_c_359_n PM_SKY130_FD_SC_HDLL__ISOBUFSRC_2%VGND
cc_1 VNB N_SLEEP_c_65_n 0.0225874f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_SLEEP_c_66_n 0.0170154f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_3 VNB N_SLEEP_c_67_n 0.0495494f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_4 VNB N_A_271_21#_c_101_n 0.0169786f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_5 VNB N_A_271_21#_c_102_n 0.020486f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_6 VNB N_A_271_21#_c_103_n 0.033547f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_7 VNB N_A_271_21#_c_104_n 6.18364e-19 $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_8 VNB N_A_271_21#_c_105_n 0.0335288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_271_21#_c_106_n 0.00446681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_271_21#_c_107_n 0.00111853f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_271_21#_c_108_n 0.00210521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_271_21#_c_109_n 0.00656081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_271_21#_c_110_n 0.00296896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB A 0.0316127f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_15 VNB A 0.00154447f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_16 VNB N_A_c_184_n 0.0337543f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_17 VNB N_A_c_185_n 0.0405294f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_18 VNB N_VPWR_c_261_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_301_n 0.00446631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_302_n 0.00262656f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_21 VNB N_X_c_303_n 0.00186872f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_22 VNB N_X_c_304_n 0.0024364f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_23 VNB N_VGND_c_347_n 0.0102948f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.105
cc_24 VNB N_VGND_c_348_n 0.0350705f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_25 VNB N_VGND_c_349_n 0.0199314f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.202
cc_26 VNB N_VGND_c_350_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_27 VNB N_VGND_c_351_n 0.00593538f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=1.17
cc_28 VNB N_VGND_c_352_n 0.0314987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_353_n 0.0201171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_354_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_355_n 0.0229836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_356_n 0.00490486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_357_n 0.0148721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_358_n 0.22467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_359_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_SLEEP_c_68_n 0.0201091f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_37 VPB N_SLEEP_c_69_n 0.0160034f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_38 VPB N_SLEEP_c_67_n 0.0226576f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_39 VPB N_A_271_21#_c_111_n 0.0161046f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_40 VPB N_A_271_21#_c_112_n 0.0192931f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.105
cc_41 VPB N_A_271_21#_c_103_n 0.0218611f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_42 VPB N_A_271_21#_c_105_n 0.0129763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_271_21#_c_107_n 0.00372552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_271_21#_c_116_n 0.0113542f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_271_21#_c_117_n 0.0119803f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_c_186_n 0.0387601f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_47 VPB N_A_c_187_n 0.0321357f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_48 VPB A 0.0386618f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_49 VPB N_A_c_184_n 0.00856578f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_50 VPB N_A_27_297#_c_217_n 0.0151236f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_51 VPB N_A_27_297#_c_218_n 0.0318598f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_52 VPB N_A_27_297#_c_219_n 0.00234749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_297#_c_220_n 0.00428099f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_54 VPB N_A_27_297#_c_221_n 0.00613585f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.17
cc_55 VPB N_A_27_297#_c_222_n 0.00186297f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_56 VPB N_A_27_297#_c_223_n 0.00458309f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=1.17
cc_57 VPB N_VPWR_c_262_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_58 VPB N_VPWR_c_263_n 0.00518f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_59 VPB N_VPWR_c_264_n 0.0549315f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_60 VPB N_VPWR_c_265_n 0.00478203f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_61 VPB N_VPWR_c_266_n 0.0142849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_261_n 0.0602703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_268_n 0.0238232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_X_c_303_n 0.00137251f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_65 N_SLEEP_c_66_n N_A_271_21#_c_101_n 0.0241348f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_66 N_SLEEP_c_69_n N_A_271_21#_c_111_n 0.00941998f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_67 SLEEP N_A_271_21#_c_103_n 8.22187e-19 $X=0.615 $Y=1.105 $X2=0 $Y2=0
cc_68 N_SLEEP_c_67_n N_A_271_21#_c_103_n 0.0241348f $X=0.985 $Y=1.202 $X2=0
+ $Y2=0
cc_69 N_SLEEP_c_68_n N_A_27_297#_c_219_n 0.0191894f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_70 N_SLEEP_c_69_n N_A_27_297#_c_219_n 0.0183679f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_71 SLEEP N_A_27_297#_c_219_n 0.0354252f $X=0.615 $Y=1.105 $X2=0 $Y2=0
cc_72 N_SLEEP_c_67_n N_A_27_297#_c_219_n 0.00826156f $X=0.985 $Y=1.202 $X2=0
+ $Y2=0
cc_73 N_SLEEP_c_68_n N_VPWR_c_262_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_74 N_SLEEP_c_69_n N_VPWR_c_262_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_75 N_SLEEP_c_69_n N_VPWR_c_264_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_76 N_SLEEP_c_68_n N_VPWR_c_261_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_77 N_SLEEP_c_69_n N_VPWR_c_261_n 0.0124344f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_78 N_SLEEP_c_68_n N_VPWR_c_268_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_79 N_SLEEP_c_65_n N_X_c_306_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_80 N_SLEEP_c_66_n N_X_c_301_n 0.0116078f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_81 SLEEP N_X_c_301_n 0.00382705f $X=0.615 $Y=1.105 $X2=0 $Y2=0
cc_82 N_SLEEP_c_65_n N_X_c_302_n 0.00243049f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_83 SLEEP N_X_c_302_n 0.0307947f $X=0.615 $Y=1.105 $X2=0 $Y2=0
cc_84 N_SLEEP_c_67_n N_X_c_302_n 0.00480108f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_85 N_SLEEP_c_69_n N_X_c_303_n 2.31783e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_86 SLEEP N_X_c_303_n 0.0060396f $X=0.615 $Y=1.105 $X2=0 $Y2=0
cc_87 N_SLEEP_c_67_n N_X_c_303_n 0.00177364f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_88 N_SLEEP_c_66_n N_X_c_315_n 5.32212e-19 $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_89 N_SLEEP_c_65_n N_VGND_c_348_n 0.0047492f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_90 N_SLEEP_c_65_n N_VGND_c_349_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_91 N_SLEEP_c_66_n N_VGND_c_349_n 0.00437852f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_92 N_SLEEP_c_66_n N_VGND_c_350_n 0.00268723f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_93 N_SLEEP_c_65_n N_VGND_c_358_n 0.0107167f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_94 N_SLEEP_c_66_n N_VGND_c_358_n 0.00615622f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_271_21#_c_116_n N_A_c_186_n 0.0109669f $X=2.68 $Y=2.28 $X2=0 $Y2=0
cc_96 N_A_271_21#_c_117_n N_A_c_186_n 0.00498925f $X=2.68 $Y=1.53 $X2=0 $Y2=0
cc_97 N_A_271_21#_c_116_n N_A_c_187_n 0.00616634f $X=2.68 $Y=2.28 $X2=0 $Y2=0
cc_98 N_A_271_21#_c_105_n A 5.27444e-19 $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_271_21#_c_106_n A 7.3318e-19 $X=2.522 $Y=1.075 $X2=0 $Y2=0
cc_100 N_A_271_21#_c_107_n A 0.00241106f $X=2.545 $Y=1.445 $X2=0 $Y2=0
cc_101 N_A_271_21#_c_110_n A 0.0156885f $X=2.522 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_271_21#_c_116_n A 0.0114011f $X=2.68 $Y=2.28 $X2=0 $Y2=0
cc_103 N_A_271_21#_c_117_n A 0.00573082f $X=2.68 $Y=1.53 $X2=0 $Y2=0
cc_104 N_A_271_21#_c_105_n N_A_c_184_n 0.00852167f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_271_21#_c_107_n N_A_c_184_n 0.00540325f $X=2.545 $Y=1.445 $X2=0 $Y2=0
cc_106 N_A_271_21#_c_110_n N_A_c_184_n 6.86672e-19 $X=2.522 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_271_21#_c_106_n N_A_c_185_n 0.00511173f $X=2.522 $Y=1.075 $X2=0 $Y2=0
cc_108 N_A_271_21#_c_108_n N_A_c_185_n 8.48614e-19 $X=2.68 $Y=0.725 $X2=0 $Y2=0
cc_109 N_A_271_21#_c_109_n N_A_c_185_n 5.53506e-19 $X=2.68 $Y=0.81 $X2=0 $Y2=0
cc_110 N_A_271_21#_c_111_n N_A_27_297#_c_220_n 3.6609e-19 $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_111 N_A_271_21#_c_111_n N_A_27_297#_c_229_n 0.0137768f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_112 N_A_271_21#_c_112_n N_A_27_297#_c_229_n 0.0143578f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_113 N_A_271_21#_c_112_n N_A_27_297#_c_221_n 9.92045e-19 $X=1.925 $Y=1.41
+ $X2=0 $Y2=0
cc_114 N_A_271_21#_c_104_n N_A_27_297#_c_221_n 0.0152874f $X=2.415 $Y=1.16 $X2=0
+ $Y2=0
cc_115 N_A_271_21#_c_105_n N_A_27_297#_c_221_n 0.00724241f $X=2.24 $Y=1.16 $X2=0
+ $Y2=0
cc_116 N_A_271_21#_c_116_n N_A_27_297#_c_221_n 0.0142206f $X=2.68 $Y=2.28 $X2=0
+ $Y2=0
cc_117 N_A_271_21#_c_117_n N_A_27_297#_c_221_n 0.0137022f $X=2.68 $Y=1.53 $X2=0
+ $Y2=0
cc_118 N_A_271_21#_c_104_n N_A_27_297#_c_222_n 9.87727e-19 $X=2.415 $Y=1.16
+ $X2=0 $Y2=0
cc_119 N_A_271_21#_c_105_n N_A_27_297#_c_222_n 6.15165e-19 $X=2.24 $Y=1.16 $X2=0
+ $Y2=0
cc_120 N_A_271_21#_c_116_n N_A_27_297#_c_222_n 0.0226472f $X=2.68 $Y=2.28 $X2=0
+ $Y2=0
cc_121 N_A_271_21#_c_116_n N_A_27_297#_c_223_n 0.00984583f $X=2.68 $Y=2.28 $X2=0
+ $Y2=0
cc_122 N_A_271_21#_c_111_n N_VPWR_c_264_n 0.00429453f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_123 N_A_271_21#_c_112_n N_VPWR_c_264_n 0.00429453f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_124 N_A_271_21#_c_116_n N_VPWR_c_264_n 0.0114468f $X=2.68 $Y=2.28 $X2=0 $Y2=0
cc_125 N_A_271_21#_M1006_s N_VPWR_c_261_n 0.00549296f $X=2.555 $Y=2.065 $X2=0
+ $Y2=0
cc_126 N_A_271_21#_c_111_n N_VPWR_c_261_n 0.00609021f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_127 N_A_271_21#_c_112_n N_VPWR_c_261_n 0.00734734f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A_271_21#_c_116_n N_VPWR_c_261_n 0.00645481f $X=2.68 $Y=2.28 $X2=0
+ $Y2=0
cc_129 N_A_271_21#_c_101_n N_X_c_301_n 0.0120386f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_271_21#_c_101_n N_X_c_303_n 0.00285675f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_271_21#_c_111_n N_X_c_303_n 0.00891542f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_271_21#_c_112_n N_X_c_303_n 8.90078e-19 $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_271_21#_c_102_n N_X_c_303_n 0.0014257f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_271_21#_c_103_n N_X_c_303_n 0.0366118f $X=2.025 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_271_21#_c_104_n N_X_c_303_n 0.00929334f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_271_21#_c_106_n N_X_c_303_n 0.00556966f $X=2.522 $Y=1.075 $X2=0 $Y2=0
cc_137 N_A_271_21#_c_107_n N_X_c_303_n 0.00579092f $X=2.545 $Y=1.445 $X2=0 $Y2=0
cc_138 N_A_271_21#_c_101_n N_X_c_304_n 0.00207804f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_271_21#_c_101_n N_X_c_315_n 0.00644736f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_271_21#_c_101_n N_VGND_c_350_n 0.00268723f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_141 N_A_271_21#_c_102_n N_VGND_c_351_n 0.00461069f $X=1.95 $Y=0.995 $X2=0
+ $Y2=0
cc_142 N_A_271_21#_c_104_n N_VGND_c_351_n 0.0129839f $X=2.415 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_271_21#_c_105_n N_VGND_c_351_n 0.00429275f $X=2.24 $Y=1.16 $X2=0
+ $Y2=0
cc_144 N_A_271_21#_c_108_n N_VGND_c_351_n 0.0119909f $X=2.68 $Y=0.725 $X2=0
+ $Y2=0
cc_145 N_A_271_21#_c_109_n N_VGND_c_351_n 0.0132324f $X=2.68 $Y=0.81 $X2=0 $Y2=0
cc_146 N_A_271_21#_c_108_n N_VGND_c_352_n 0.00846051f $X=2.68 $Y=0.725 $X2=0
+ $Y2=0
cc_147 N_A_271_21#_c_101_n N_VGND_c_353_n 0.00423334f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_271_21#_c_102_n N_VGND_c_353_n 0.00585385f $X=1.95 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_271_21#_c_108_n N_VGND_c_355_n 0.00509579f $X=2.68 $Y=0.725 $X2=0
+ $Y2=0
cc_150 N_A_271_21#_c_109_n N_VGND_c_355_n 0.00273515f $X=2.68 $Y=0.81 $X2=0
+ $Y2=0
cc_151 N_A_271_21#_c_101_n N_VGND_c_358_n 0.00598581f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_271_21#_c_102_n N_VGND_c_358_n 0.0121055f $X=1.95 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_271_21#_c_108_n N_VGND_c_358_n 0.0055979f $X=2.68 $Y=0.725 $X2=0
+ $Y2=0
cc_154 N_A_271_21#_c_109_n N_VGND_c_358_n 0.00480544f $X=2.68 $Y=0.81 $X2=0
+ $Y2=0
cc_155 N_A_c_186_n N_A_27_297#_c_221_n 8.51322e-19 $X=2.915 $Y=1.89 $X2=0 $Y2=0
cc_156 N_A_c_187_n N_VPWR_c_263_n 0.00479105f $X=2.915 $Y=1.99 $X2=0 $Y2=0
cc_157 N_A_c_187_n N_VPWR_c_264_n 0.00743866f $X=2.915 $Y=1.99 $X2=0 $Y2=0
cc_158 A N_VPWR_c_266_n 0.00343264f $X=3.34 $Y=1.445 $X2=0 $Y2=0
cc_159 N_A_c_187_n N_VPWR_c_261_n 0.0154317f $X=2.915 $Y=1.99 $X2=0 $Y2=0
cc_160 A N_VPWR_c_261_n 0.0058652f $X=3.34 $Y=1.445 $X2=0 $Y2=0
cc_161 N_A_c_185_n N_VGND_c_351_n 0.00722462f $X=2.982 $Y=0.995 $X2=0 $Y2=0
cc_162 A N_VGND_c_352_n 0.0171282f $X=3.34 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A_c_184_n N_VGND_c_352_n 0.00306423f $X=2.965 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_c_185_n N_VGND_c_352_n 0.0154087f $X=2.982 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_185_n N_VGND_c_355_n 0.00585385f $X=2.982 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_c_185_n N_VGND_c_358_n 0.0132862f $X=2.982 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_27_297#_c_219_n N_VPWR_M1000_d 0.00188315f $X=1.095 $Y=1.55 $X2=-0.19
+ $Y2=1.305
cc_168 N_A_27_297#_c_219_n N_VPWR_c_262_n 0.0145257f $X=1.095 $Y=1.55 $X2=0
+ $Y2=0
cc_169 N_A_27_297#_c_243_p N_VPWR_c_264_n 0.015002f $X=1.22 $Y=2.295 $X2=0 $Y2=0
cc_170 N_A_27_297#_c_229_n N_VPWR_c_264_n 0.0386815f $X=2.035 $Y=2.38 $X2=0
+ $Y2=0
cc_171 N_A_27_297#_c_223_n N_VPWR_c_264_n 0.0191283f $X=2.18 $Y=2.295 $X2=0
+ $Y2=0
cc_172 N_A_27_297#_M1000_s N_VPWR_c_261_n 0.00303344f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_173 N_A_27_297#_M1007_s N_VPWR_c_261_n 0.00297222f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_174 N_A_27_297#_M1003_d N_VPWR_c_261_n 0.00217519f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_175 N_A_27_297#_c_218_n N_VPWR_c_261_n 0.0122467f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_176 N_A_27_297#_c_243_p N_VPWR_c_261_n 0.00962794f $X=1.22 $Y=2.295 $X2=0
+ $Y2=0
cc_177 N_A_27_297#_c_229_n N_VPWR_c_261_n 0.0239144f $X=2.035 $Y=2.38 $X2=0
+ $Y2=0
cc_178 N_A_27_297#_c_223_n N_VPWR_c_261_n 0.0111575f $X=2.18 $Y=2.295 $X2=0
+ $Y2=0
cc_179 N_A_27_297#_c_218_n N_VPWR_c_268_n 0.0211751f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_180 N_A_27_297#_c_229_n N_X_M1002_s 0.00352392f $X=2.035 $Y=2.38 $X2=0 $Y2=0
cc_181 N_A_27_297#_c_219_n N_X_c_301_n 0.00338008f $X=1.095 $Y=1.55 $X2=0 $Y2=0
cc_182 N_A_27_297#_c_220_n N_X_c_301_n 0.00932875f $X=1.22 $Y=1.655 $X2=0 $Y2=0
cc_183 N_A_27_297#_c_220_n N_X_c_303_n 0.00915792f $X=1.22 $Y=1.655 $X2=0 $Y2=0
cc_184 N_A_27_297#_c_229_n N_X_c_303_n 0.0147284f $X=2.035 $Y=2.38 $X2=0 $Y2=0
cc_185 N_A_27_297#_c_221_n N_X_c_303_n 0.00262991f $X=2.16 $Y=1.63 $X2=0 $Y2=0
cc_186 N_A_27_297#_c_217_n N_VGND_c_348_n 0.0114749f $X=0.245 $Y=1.655 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_261_n N_X_M1002_s 0.00232895f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_188 N_X_c_301_n N_VGND_M1009_s 0.00161804f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_189 N_X_c_302_n N_VGND_c_348_n 0.00752789f $X=0.915 $Y=0.81 $X2=0 $Y2=0
cc_190 N_X_c_306_n N_VGND_c_349_n 0.0231581f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_191 N_X_c_301_n N_VGND_c_349_n 0.00253779f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_192 N_X_c_301_n N_VGND_c_350_n 0.0122105f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_193 N_X_c_304_n N_VGND_c_351_n 6.33233e-19 $X=1.665 $Y=0.81 $X2=0 $Y2=0
cc_194 N_X_c_301_n N_VGND_c_353_n 0.00198102f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_195 N_X_c_315_n N_VGND_c_353_n 0.023237f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_196 N_X_M1004_d N_VGND_c_358_n 0.00304143f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_197 N_X_M1005_s N_VGND_c_358_n 0.00364931f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_198 N_X_c_306_n N_VGND_c_358_n 0.0143294f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_199 N_X_c_301_n N_VGND_c_358_n 0.00945827f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_200 N_X_c_315_n N_VGND_c_358_n 0.0143471f $X=1.69 $Y=0.39 $X2=0 $Y2=0
