* NGSPICE file created from sky130_fd_sc_hdll__nand3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nand3b_2 A_N B C VGND VNB VPB VPWR Y
M1000 VGND C a_228_47# VNB nshort w=650000u l=150000u
+  ad=4.295e+11p pd=4.01e+06u as=4.485e+11p ps=3.98e+06u
M1001 Y a_27_47# a_448_47# VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=5.46e+11p ps=5.58e+06u
M1002 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=1.4657e+12p pd=1.303e+07u as=1.134e+11p ps=1.38e+06u
M1003 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=0p ps=0u
M1004 a_448_47# B a_228_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_228_47# B a_448_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_228_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_448_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends

