* File: sky130_fd_sc_hdll__a221oi_4.pxi.spice
* Created: Wed Sep  2 08:18:16 2020
* 
x_PM_SKY130_FD_SC_HDLL__A221OI_4%C1 N_C1_c_128_n N_C1_M1003_g N_C1_c_122_n
+ N_C1_M1007_g N_C1_c_129_n N_C1_M1010_g N_C1_c_123_n N_C1_M1020_g N_C1_c_130_n
+ N_C1_M1016_g N_C1_c_124_n N_C1_M1024_g N_C1_c_131_n N_C1_M1028_g N_C1_c_125_n
+ N_C1_M1033_g C1 N_C1_c_126_n N_C1_c_127_n PM_SKY130_FD_SC_HDLL__A221OI_4%C1
x_PM_SKY130_FD_SC_HDLL__A221OI_4%B2 N_B2_c_198_n N_B2_M1001_g N_B2_c_199_n
+ N_B2_M1015_g N_B2_c_206_n N_B2_M1014_g N_B2_c_200_n N_B2_M1027_g N_B2_c_207_n
+ N_B2_M1018_g N_B2_c_208_n N_B2_M1030_g N_B2_c_201_n N_B2_M1034_g N_B2_c_202_n
+ N_B2_M1036_g N_B2_c_203_n N_B2_c_204_n N_B2_c_205_n N_B2_c_213_n B2 B2
+ PM_SKY130_FD_SC_HDLL__A221OI_4%B2
x_PM_SKY130_FD_SC_HDLL__A221OI_4%B1 N_B1_c_319_n N_B1_M1021_g N_B1_c_325_n
+ N_B1_M1004_g N_B1_c_320_n N_B1_M1022_g N_B1_c_326_n N_B1_M1012_g N_B1_c_321_n
+ N_B1_M1029_g N_B1_c_327_n N_B1_M1026_g N_B1_c_328_n N_B1_M1032_g N_B1_c_322_n
+ N_B1_M1038_g B1 N_B1_c_323_n N_B1_c_324_n B1 PM_SKY130_FD_SC_HDLL__A221OI_4%B1
x_PM_SKY130_FD_SC_HDLL__A221OI_4%A2 N_A2_c_385_n N_A2_M1005_g N_A2_c_386_n
+ N_A2_M1006_g N_A2_c_387_n N_A2_M1009_g N_A2_c_396_n N_A2_M1008_g N_A2_c_388_n
+ N_A2_M1025_g N_A2_c_397_n N_A2_M1013_g N_A2_c_389_n N_A2_M1037_g N_A2_c_398_n
+ N_A2_M1023_g N_A2_c_399_n N_A2_c_390_n N_A2_c_391_n N_A2_c_392_n A2
+ N_A2_c_393_n N_A2_c_394_n A2 PM_SKY130_FD_SC_HDLL__A221OI_4%A2
x_PM_SKY130_FD_SC_HDLL__A221OI_4%A1 N_A1_c_507_n N_A1_M1002_g N_A1_c_513_n
+ N_A1_M1000_g N_A1_c_508_n N_A1_M1011_g N_A1_c_514_n N_A1_M1019_g N_A1_c_509_n
+ N_A1_M1017_g N_A1_c_515_n N_A1_M1031_g N_A1_c_516_n N_A1_M1035_g N_A1_c_510_n
+ N_A1_M1039_g A1 N_A1_c_511_n N_A1_c_512_n A1 PM_SKY130_FD_SC_HDLL__A221OI_4%A1
x_PM_SKY130_FD_SC_HDLL__A221OI_4%A_27_297# N_A_27_297#_M1003_s
+ N_A_27_297#_M1010_s N_A_27_297#_M1028_s N_A_27_297#_M1014_s
+ N_A_27_297#_M1030_s N_A_27_297#_M1012_d N_A_27_297#_M1032_d
+ N_A_27_297#_c_567_n N_A_27_297#_c_568_n N_A_27_297#_c_576_n
+ N_A_27_297#_c_606_p N_A_27_297#_c_578_n N_A_27_297#_c_569_n
+ N_A_27_297#_c_570_n N_A_27_297#_c_571_n N_A_27_297#_c_572_n
+ N_A_27_297#_c_590_n N_A_27_297#_c_591_n N_A_27_297#_c_592_n
+ N_A_27_297#_c_635_p PM_SKY130_FD_SC_HDLL__A221OI_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A221OI_4%Y N_Y_M1007_d N_Y_M1024_d N_Y_M1021_s
+ N_Y_M1029_s N_Y_M1002_s N_Y_M1017_s N_Y_M1003_d N_Y_M1016_d N_Y_c_661_n
+ N_Y_c_734_n N_Y_c_657_n N_Y_c_658_n N_Y_c_648_n N_Y_c_649_n N_Y_c_676_n
+ N_Y_c_738_n N_Y_c_650_n N_Y_c_651_n N_Y_c_652_n N_Y_c_700_n N_Y_c_726_n
+ N_Y_c_653_n N_Y_c_659_n N_Y_c_660_n N_Y_c_702_n N_Y_c_654_n N_Y_c_655_n
+ N_Y_c_656_n Y PM_SKY130_FD_SC_HDLL__A221OI_4%Y
x_PM_SKY130_FD_SC_HDLL__A221OI_4%A_511_297# N_A_511_297#_M1014_d
+ N_A_511_297#_M1018_d N_A_511_297#_M1004_s N_A_511_297#_M1026_s
+ N_A_511_297#_M1034_d N_A_511_297#_M1000_d N_A_511_297#_M1031_d
+ N_A_511_297#_M1008_s N_A_511_297#_M1023_s N_A_511_297#_c_842_n
+ N_A_511_297#_c_844_n N_A_511_297#_c_800_n N_A_511_297#_c_805_n
+ N_A_511_297#_c_866_p N_A_511_297#_c_814_n N_A_511_297#_c_860_p
+ N_A_511_297#_c_819_n N_A_511_297#_c_795_n N_A_511_297#_c_796_n
+ N_A_511_297#_c_873_p N_A_511_297#_c_831_n
+ PM_SKY130_FD_SC_HDLL__A221OI_4%A_511_297#
x_PM_SKY130_FD_SC_HDLL__A221OI_4%VPWR N_VPWR_M1005_d N_VPWR_M1019_s
+ N_VPWR_M1035_s N_VPWR_M1013_d N_VPWR_c_890_n N_VPWR_c_891_n N_VPWR_c_892_n
+ N_VPWR_c_893_n N_VPWR_c_894_n VPWR N_VPWR_c_895_n N_VPWR_c_896_n
+ N_VPWR_c_889_n N_VPWR_c_898_n PM_SKY130_FD_SC_HDLL__A221OI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A221OI_4%VGND N_VGND_M1007_s N_VGND_M1020_s
+ N_VGND_M1033_s N_VGND_M1015_s N_VGND_M1036_s N_VGND_M1009_s N_VGND_M1037_s
+ N_VGND_c_997_n N_VGND_c_998_n N_VGND_c_999_n N_VGND_c_1000_n N_VGND_c_1001_n
+ N_VGND_c_1002_n N_VGND_c_1003_n N_VGND_c_1004_n N_VGND_c_1005_n
+ N_VGND_c_1006_n N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n
+ N_VGND_c_1010_n N_VGND_c_1011_n N_VGND_c_1012_n N_VGND_c_1013_n
+ N_VGND_c_1014_n VGND N_VGND_c_1015_n N_VGND_c_1016_n N_VGND_c_1017_n
+ PM_SKY130_FD_SC_HDLL__A221OI_4%VGND
x_PM_SKY130_FD_SC_HDLL__A221OI_4%A_503_47# N_A_503_47#_M1001_d
+ N_A_503_47#_M1027_d N_A_503_47#_M1022_d N_A_503_47#_M1038_d
+ N_A_503_47#_c_1140_n N_A_503_47#_c_1141_n N_A_503_47#_c_1143_n
+ N_A_503_47#_c_1144_n N_A_503_47#_c_1145_n
+ PM_SKY130_FD_SC_HDLL__A221OI_4%A_503_47#
x_PM_SKY130_FD_SC_HDLL__A221OI_4%A_1375_47# N_A_1375_47#_M1006_d
+ N_A_1375_47#_M1011_d N_A_1375_47#_M1039_d N_A_1375_47#_M1025_d
+ N_A_1375_47#_c_1178_n N_A_1375_47#_c_1179_n N_A_1375_47#_c_1176_n
+ N_A_1375_47#_c_1177_n N_A_1375_47#_c_1190_n
+ PM_SKY130_FD_SC_HDLL__A221OI_4%A_1375_47#
cc_1 VNB N_C1_c_122_n 0.0221022f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB N_C1_c_123_n 0.0167451f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_3 VNB N_C1_c_124_n 0.0167287f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.995
cc_4 VNB N_C1_c_125_n 0.017295f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_5 VNB N_C1_c_126_n 0.0134887f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=1.16
cc_6 VNB N_C1_c_127_n 0.0901852f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_7 VNB N_B2_c_198_n 0.0169232f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_8 VNB N_B2_c_199_n 0.0165913f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_9 VNB N_B2_c_200_n 0.020402f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_10 VNB N_B2_c_201_n 0.0213486f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_11 VNB N_B2_c_202_n 0.0175607f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_12 VNB N_B2_c_203_n 0.00331183f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_13 VNB N_B2_c_204_n 0.0057377f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_14 VNB N_B2_c_205_n 0.0865617f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_15 VNB N_B1_c_319_n 0.0207849f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_16 VNB N_B1_c_320_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_17 VNB N_B1_c_321_n 0.0174167f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_18 VNB N_B1_c_322_n 0.0176283f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_19 VNB N_B1_c_323_n 0.00219191f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=1.202
cc_20 VNB N_B1_c_324_n 0.0733353f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_21 VNB N_A2_c_385_n 0.0219152f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_22 VNB N_A2_c_386_n 0.0171042f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_23 VNB N_A2_c_387_n 0.0164927f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_24 VNB N_A2_c_388_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_25 VNB N_A2_c_389_n 0.0218461f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_26 VNB N_A2_c_390_n 2.86539e-19 $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_27 VNB N_A2_c_391_n 0.00352367f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_28 VNB N_A2_c_392_n 0.00188267f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=1.16
cc_29 VNB N_A2_c_393_n 0.0133375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A2_c_394_n 0.0656014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A1_c_507_n 0.0167267f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_32 VNB N_A1_c_508_n 0.0169715f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_33 VNB N_A1_c_509_n 0.0174157f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_34 VNB N_A1_c_510_n 0.0171706f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_35 VNB N_A1_c_511_n 0.00262678f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=1.16
cc_36 VNB N_A1_c_512_n 0.0730066f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_37 VNB N_Y_c_648_n 0.00264748f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=1.16
cc_38 VNB N_Y_c_649_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=1.16
cc_39 VNB N_Y_c_650_n 0.00159487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_651_n 0.00878555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_652_n 0.00169546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_Y_c_653_n 0.0013877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_654_n 7.82359e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Y_c_655_n 0.00784774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_Y_c_656_n 0.00270091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VPWR_c_889_n 0.440529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_997_n 0.0106747f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_48 VNB N_VGND_c_998_n 0.0316509f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_49 VNB N_VGND_c_999_n 0.0199148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_1000_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_51 VNB N_VGND_c_1001_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=1.16
cc_52 VNB N_VGND_c_1002_n 0.00197226f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.202
cc_53 VNB N_VGND_c_1003_n 0.00469188f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.202
cc_54 VNB N_VGND_c_1004_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1005_n 0.0132827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1006_n 0.00697284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1007_n 0.0201004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1008_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1009_n 0.00140268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1010_n 0.00404437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1011_n 0.0958324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1012_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1013_n 0.0608286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1014_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1015_n 0.0184128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1016_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1017_n 0.489681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1375_47#_c_1176_n 0.00326213f $X=-0.19 $Y=-0.24 $X2=1.925
+ $Y2=1.985
cc_69 VNB N_A_1375_47#_c_1177_n 0.00499593f $X=-0.19 $Y=-0.24 $X2=1.925
+ $Y2=1.985
cc_70 VPB N_C1_c_128_n 0.0200174f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_71 VPB N_C1_c_129_n 0.0158724f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_72 VPB N_C1_c_130_n 0.0158628f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_73 VPB N_C1_c_131_n 0.0196979f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_74 VPB N_C1_c_127_n 0.055155f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_75 VPB N_B2_c_206_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_76 VPB N_B2_c_207_n 0.0162441f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_77 VPB N_B2_c_208_n 0.0159879f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.995
cc_78 VPB N_B2_c_201_n 0.0249939f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_79 VPB N_B2_c_203_n 0.00236005f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_80 VPB N_B2_c_204_n 0.00194983f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.202
cc_81 VPB N_B2_c_205_n 0.0505654f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_82 VPB N_B2_c_213_n 0.0101902f $X=-0.19 $Y=1.305 $X2=1.27 $Y2=1.16
cc_83 VPB N_B1_c_325_n 0.0159748f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_84 VPB N_B1_c_326_n 0.0158725f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_85 VPB N_B1_c_327_n 0.0158728f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.995
cc_86 VPB N_B1_c_328_n 0.015977f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_87 VPB N_B1_c_324_n 0.0449447f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_88 VPB N_A2_c_385_n 0.0250485f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_89 VPB N_A2_c_396_n 0.015606f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_90 VPB N_A2_c_397_n 0.0158836f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.995
cc_91 VPB N_A2_c_398_n 0.0201091f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.995
cc_92 VPB N_A2_c_399_n 0.0121431f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_93 VPB N_A2_c_390_n 0.00137605f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_94 VPB N_A2_c_391_n 0.00272122f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_95 VPB N_A2_c_394_n 0.0369838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A1_c_513_n 0.014886f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_97 VPB N_A1_c_514_n 0.0148232f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_98 VPB N_A1_c_515_n 0.0148054f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.995
cc_99 VPB N_A1_c_516_n 0.0148676f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_100 VPB N_A1_c_512_n 0.0449781f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_101 VPB N_A_27_297#_c_567_n 0.00753428f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.995
cc_102 VPB N_A_27_297#_c_568_n 0.0360658f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_103 VPB N_A_27_297#_c_569_n 0.00196379f $X=-0.19 $Y=1.305 $X2=1.27 $Y2=1.16
cc_104 VPB N_A_27_297#_c_570_n 0.00762043f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.202
cc_105 VPB N_A_27_297#_c_571_n 0.0148655f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.202
cc_106 VPB N_A_27_297#_c_572_n 0.00307685f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_107 VPB N_Y_c_657_n 0.00196322f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.202
cc_108 VPB N_Y_c_658_n 0.00184379f $X=-0.19 $Y=1.305 $X2=1.27 $Y2=1.202
cc_109 VPB N_Y_c_659_n 0.00112154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_Y_c_660_n 6.96187e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_511_297#_c_795_n 0.00656714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_511_297#_c_796_n 0.00115709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_890_n 0.00420672f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_114 VPB N_VPWR_c_891_n 0.00417211f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.56
cc_115 VPB N_VPWR_c_892_n 0.156448f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_116 VPB N_VPWR_c_893_n 0.0171758f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_117 VPB N_VPWR_c_894_n 0.00324402f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_118 VPB N_VPWR_c_895_n 0.022126f $X=-0.19 $Y=1.305 $X2=1.27 $Y2=1.202
cc_119 VPB N_VPWR_c_896_n 0.0209718f $X=-0.19 $Y=1.305 $X2=1.27 $Y2=1.175
cc_120 VPB N_VPWR_c_889_n 0.0566639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_898_n 0.00409747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 N_C1_c_125_n N_B2_c_198_n 0.0181726f $X=1.95 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_123 N_C1_c_127_n N_B2_c_205_n 0.0181726f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_124 N_C1_c_128_n N_A_27_297#_c_568_n 9.99407e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_125 N_C1_c_126_n N_A_27_297#_c_568_n 0.0264267f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_126 N_C1_c_127_n N_A_27_297#_c_568_n 0.00195514f $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_127 N_C1_c_128_n N_A_27_297#_c_576_n 0.0143578f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_128 N_C1_c_129_n N_A_27_297#_c_576_n 0.0143578f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_129 N_C1_c_130_n N_A_27_297#_c_578_n 0.0143578f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_130 N_C1_c_131_n N_A_27_297#_c_578_n 0.0143578f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_131 N_C1_c_131_n N_A_27_297#_c_572_n 0.0016132f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_132 N_C1_c_122_n N_Y_c_661_n 0.00738878f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_133 N_C1_c_129_n N_Y_c_657_n 0.015669f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_134 N_C1_c_130_n N_Y_c_657_n 0.0170044f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_135 N_C1_c_126_n N_Y_c_657_n 0.0395588f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_136 N_C1_c_127_n N_Y_c_657_n 0.00883832f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_137 N_C1_c_128_n N_Y_c_658_n 4.00176e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_138 N_C1_c_126_n N_Y_c_658_n 0.020385f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_139 N_C1_c_127_n N_Y_c_658_n 0.00663436f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_140 N_C1_c_123_n N_Y_c_648_n 0.0109479f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_141 N_C1_c_124_n N_Y_c_648_n 0.00666956f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_142 N_C1_c_126_n N_Y_c_648_n 0.0370948f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_143 N_C1_c_127_n N_Y_c_648_n 0.00345541f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_144 N_C1_c_122_n N_Y_c_649_n 0.00435558f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_145 N_C1_c_126_n N_Y_c_649_n 0.0305116f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_146 N_C1_c_127_n N_Y_c_649_n 0.00358305f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_147 N_C1_c_123_n N_Y_c_676_n 5.82315e-19 $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_148 N_C1_c_124_n N_Y_c_676_n 0.00850899f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_149 N_C1_c_124_n N_Y_c_650_n 0.00211295f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_150 N_C1_c_125_n N_Y_c_650_n 0.00201157f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_151 N_C1_c_126_n N_Y_c_650_n 0.00116136f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_152 N_C1_c_127_n N_Y_c_650_n 0.0106273f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_153 N_C1_c_127_n N_Y_c_651_n 0.0203077f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_154 N_C1_c_124_n N_Y_c_653_n 0.00352025f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_155 N_C1_c_125_n N_Y_c_653_n 2.01404e-19 $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_156 N_C1_c_127_n N_Y_c_653_n 3.16161e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_157 N_C1_c_130_n N_Y_c_659_n 7.90806e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_158 N_C1_c_131_n N_Y_c_659_n 0.00162979f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_159 N_C1_c_127_n N_Y_c_659_n 0.0144805f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_160 N_C1_c_131_n N_Y_c_660_n 0.00351929f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_161 N_C1_c_127_n N_Y_c_660_n 0.00307505f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_162 N_C1_c_126_n Y 0.0123026f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_163 N_C1_c_127_n Y 0.00635817f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_164 N_C1_c_128_n N_VPWR_c_892_n 0.00429453f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_165 N_C1_c_129_n N_VPWR_c_892_n 0.00429453f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_166 N_C1_c_130_n N_VPWR_c_892_n 0.00429453f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_167 N_C1_c_131_n N_VPWR_c_892_n 0.00429453f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_168 N_C1_c_128_n N_VPWR_c_889_n 0.00699455f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_169 N_C1_c_129_n N_VPWR_c_889_n 0.00606499f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_170 N_C1_c_130_n N_VPWR_c_889_n 0.00606499f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_171 N_C1_c_131_n N_VPWR_c_889_n 0.00734734f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_172 N_C1_c_122_n N_VGND_c_998_n 0.0064202f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_173 N_C1_c_126_n N_VGND_c_998_n 0.020187f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_174 N_C1_c_127_n N_VGND_c_998_n 9.96531e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_175 N_C1_c_122_n N_VGND_c_999_n 0.00465454f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_176 N_C1_c_123_n N_VGND_c_999_n 0.00437852f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_177 N_C1_c_123_n N_VGND_c_1000_n 0.00276126f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_178 N_C1_c_124_n N_VGND_c_1000_n 0.00359159f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_179 N_C1_c_125_n N_VGND_c_1001_n 0.00309199f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_180 N_C1_c_125_n N_VGND_c_1002_n 0.00160437f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_181 N_C1_c_124_n N_VGND_c_1007_n 0.00396605f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_182 N_C1_c_125_n N_VGND_c_1007_n 0.00585385f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_183 N_C1_c_122_n N_VGND_c_1017_n 0.00891695f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_184 N_C1_c_123_n N_VGND_c_1017_n 0.00614065f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_185 N_C1_c_124_n N_VGND_c_1017_n 0.00581484f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_186 N_C1_c_125_n N_VGND_c_1017_n 0.0108539f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B2_c_208_n N_B1_c_325_n 0.0374168f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B2_c_204_n N_B1_c_325_n 8.17193e-19 $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B2_c_213_n N_B1_c_325_n 0.0129351f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_190 N_B2_c_213_n N_B1_c_326_n 0.0122688f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_191 N_B2_c_213_n N_B1_c_327_n 0.0122688f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_192 N_B2_c_201_n N_B1_c_328_n 0.037179f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B2_c_203_n N_B1_c_328_n 7.96475e-19 $X=6.23 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B2_c_213_n N_B1_c_328_n 0.0122258f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_195 N_B2_c_202_n N_B1_c_322_n 0.0219111f $X=6.28 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B2_c_201_n N_B1_c_323_n 7.88936e-19 $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B2_c_203_n N_B1_c_323_n 0.0160446f $X=6.23 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B2_c_204_n N_B1_c_323_n 0.0237848f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B2_c_205_n N_B1_c_323_n 2.46885e-19 $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B2_c_213_n N_B1_c_323_n 0.112534f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_201 N_B2_c_201_n N_B1_c_324_n 0.0250948f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B2_c_203_n N_B1_c_324_n 0.0038839f $X=6.23 $Y=1.16 $X2=0 $Y2=0
cc_203 N_B2_c_204_n N_B1_c_324_n 0.00556182f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B2_c_205_n N_B1_c_324_n 0.0219886f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B2_c_213_n N_B1_c_324_n 0.0232076f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_206 N_B2_c_201_n N_A2_c_385_n 0.0443456f $X=6.255 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_207 N_B2_c_203_n N_A2_c_385_n 0.00113245f $X=6.23 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_208 N_B2_c_213_n N_A2_c_385_n 5.68289e-19 $X=6.065 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_209 N_B2_c_202_n N_A2_c_386_n 0.0186142f $X=6.28 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B2_c_201_n N_A2_c_391_n 0.00178688f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B2_c_203_n N_A2_c_391_n 0.0305615f $X=6.23 $Y=1.16 $X2=0 $Y2=0
cc_212 N_B2_c_213_n N_A2_c_391_n 0.0144432f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_213 N_B2_c_204_n N_A_27_297#_M1030_s 0.00140009f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_214 N_B2_c_213_n N_A_27_297#_M1030_s 7.3922e-19 $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_215 N_B2_c_213_n N_A_27_297#_M1012_d 0.00209843f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_216 N_B2_c_213_n N_A_27_297#_M1032_d 0.00209198f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_217 N_B2_c_206_n N_A_27_297#_c_570_n 0.00475474f $X=2.965 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B2_c_206_n N_A_27_297#_c_571_n 0.0140935f $X=2.965 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B2_c_207_n N_A_27_297#_c_571_n 6.83314e-19 $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_220 N_B2_c_204_n N_A_27_297#_c_571_n 0.00318935f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_221 N_B2_c_205_n N_A_27_297#_c_571_n 0.0210586f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B2_c_206_n N_A_27_297#_c_590_n 0.00287251f $X=2.965 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B2_c_206_n N_A_27_297#_c_591_n 0.00813791f $X=2.965 $Y=1.41 $X2=0 $Y2=0
cc_224 N_B2_c_207_n N_A_27_297#_c_592_n 0.0132705f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B2_c_208_n N_A_27_297#_c_592_n 0.0125727f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_226 N_B2_c_201_n N_A_27_297#_c_592_n 0.00317006f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_227 N_B2_c_204_n N_A_27_297#_c_592_n 0.0153529f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_228 N_B2_c_205_n N_A_27_297#_c_592_n 0.00538323f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_229 N_B2_c_213_n N_A_27_297#_c_592_n 0.0884371f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_230 N_B2_c_205_n N_Y_c_650_n 5.32366e-19 $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_231 N_B2_c_204_n N_Y_c_651_n 0.0146462f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_232 N_B2_c_205_n N_Y_c_651_n 0.054193f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_233 N_B2_c_199_n N_Y_c_652_n 4.24414e-19 $X=2.91 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B2_c_200_n N_Y_c_652_n 0.00595921f $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B2_c_204_n N_Y_c_652_n 0.00739304f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_236 N_B2_c_205_n N_Y_c_652_n 0.0107761f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_237 N_B2_c_200_n N_Y_c_700_n 0.00779761f $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B2_c_205_n N_Y_c_659_n 2.65049e-19 $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_239 N_B2_c_201_n N_Y_c_702_n 3.45898e-19 $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_240 N_B2_c_203_n N_Y_c_702_n 0.00259121f $X=6.23 $Y=1.16 $X2=0 $Y2=0
cc_241 N_B2_c_204_n N_Y_c_702_n 0.0304856f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_242 N_B2_c_205_n N_Y_c_702_n 0.00823233f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B2_c_213_n N_Y_c_702_n 0.00821641f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_244 N_B2_c_201_n N_Y_c_654_n 0.00254901f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_245 N_B2_c_202_n N_Y_c_654_n 0.00892152f $X=6.28 $Y=0.995 $X2=0 $Y2=0
cc_246 N_B2_c_203_n N_Y_c_654_n 0.0232935f $X=6.23 $Y=1.16 $X2=0 $Y2=0
cc_247 N_B2_c_201_n N_Y_c_655_n 0.00123166f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B2_c_202_n N_Y_c_655_n 0.00651024f $X=6.28 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B2_c_213_n N_A_511_297#_M1004_s 0.00209843f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_250 N_B2_c_213_n N_A_511_297#_M1026_s 0.00209843f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_251 N_B2_c_213_n N_A_511_297#_M1034_d 0.00118227f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_252 N_B2_c_206_n N_A_511_297#_c_800_n 0.0134692f $X=2.965 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B2_c_207_n N_A_511_297#_c_800_n 0.0112654f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B2_c_208_n N_A_511_297#_c_800_n 0.0112018f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B2_c_201_n N_A_511_297#_c_800_n 0.0134026f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B2_c_213_n N_A_511_297#_c_800_n 0.00435428f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_257 N_B2_c_213_n N_A_511_297#_c_805_n 4.44748e-19 $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_258 N_B2_c_201_n N_VPWR_c_891_n 0.00102327f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B2_c_206_n N_VPWR_c_892_n 0.00429453f $X=2.965 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B2_c_207_n N_VPWR_c_892_n 0.00429453f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B2_c_208_n N_VPWR_c_892_n 0.00429453f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B2_c_201_n N_VPWR_c_892_n 0.00429453f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B2_c_206_n N_VPWR_c_889_n 0.00734734f $X=2.965 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B2_c_207_n N_VPWR_c_889_n 0.00606499f $X=3.435 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B2_c_208_n N_VPWR_c_889_n 0.00609118f $X=3.905 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B2_c_201_n N_VPWR_c_889_n 0.00623066f $X=6.255 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B2_c_198_n N_VGND_c_1001_n 0.00825648f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_268 N_B2_c_202_n N_VGND_c_1003_n 0.00526373f $X=6.28 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B2_c_200_n N_VGND_c_1009_n 0.00206565f $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B2_c_205_n N_VGND_c_1009_n 0.00333976f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_271 N_B2_c_198_n N_VGND_c_1010_n 0.0155874f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_272 N_B2_c_199_n N_VGND_c_1010_n 0.0123914f $X=2.91 $Y=0.995 $X2=0 $Y2=0
cc_273 N_B2_c_205_n N_VGND_c_1010_n 0.00358041f $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_274 N_B2_c_198_n N_VGND_c_1011_n 0.00389931f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_275 N_B2_c_199_n N_VGND_c_1011_n 0.00357877f $X=2.91 $Y=0.995 $X2=0 $Y2=0
cc_276 N_B2_c_200_n N_VGND_c_1011_n 0.00357877f $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_277 N_B2_c_202_n N_VGND_c_1011_n 0.00432885f $X=6.28 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B2_c_198_n N_VGND_c_1017_n 0.00584654f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_279 N_B2_c_199_n N_VGND_c_1017_n 0.00548399f $X=2.91 $Y=0.995 $X2=0 $Y2=0
cc_280 N_B2_c_200_n N_VGND_c_1017_n 0.00668309f $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_281 N_B2_c_202_n N_VGND_c_1017_n 0.00632328f $X=6.28 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B2_c_198_n N_A_503_47#_c_1140_n 0.00491153f $X=2.44 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_B2_c_200_n N_A_503_47#_c_1141_n 0.00625674f $X=3.38 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_B2_c_205_n N_A_503_47#_c_1141_n 4.01412e-19 $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B2_c_205_n N_A_503_47#_c_1143_n 2.232e-19 $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_286 N_B2_c_199_n N_A_503_47#_c_1144_n 0.00173979f $X=2.91 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_B2_c_199_n N_A_503_47#_c_1145_n 0.00721438f $X=2.91 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_B2_c_200_n N_A_503_47#_c_1145_n 0.00378632f $X=3.38 $Y=0.995 $X2=0
+ $Y2=0
cc_289 N_B2_c_205_n N_A_503_47#_c_1145_n 3.07254e-19 $X=3.85 $Y=1.16 $X2=0 $Y2=0
cc_290 N_B1_c_325_n N_A_27_297#_c_592_n 0.0113499f $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_291 N_B1_c_326_n N_A_27_297#_c_592_n 0.0113499f $X=4.845 $Y=1.41 $X2=0 $Y2=0
cc_292 N_B1_c_327_n N_A_27_297#_c_592_n 0.0113499f $X=5.315 $Y=1.41 $X2=0 $Y2=0
cc_293 N_B1_c_328_n N_A_27_297#_c_592_n 0.0113499f $X=5.785 $Y=1.41 $X2=0 $Y2=0
cc_294 N_B1_c_319_n N_Y_c_652_n 0.0036334f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_295 N_B1_c_319_n N_Y_c_702_n 0.0115069f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_296 N_B1_c_320_n N_Y_c_702_n 0.00882716f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B1_c_321_n N_Y_c_702_n 0.00882716f $X=5.29 $Y=0.995 $X2=0 $Y2=0
cc_298 N_B1_c_322_n N_Y_c_702_n 0.00877034f $X=5.81 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B1_c_323_n N_Y_c_702_n 0.0970818f $X=5.67 $Y=1.16 $X2=0 $Y2=0
cc_300 N_B1_c_324_n N_Y_c_702_n 0.010511f $X=5.785 $Y=1.202 $X2=0 $Y2=0
cc_301 N_B1_c_322_n N_Y_c_654_n 0.00220022f $X=5.81 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B1_c_325_n N_A_511_297#_c_800_n 0.0112018f $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_303 N_B1_c_326_n N_A_511_297#_c_800_n 0.0112654f $X=4.845 $Y=1.41 $X2=0 $Y2=0
cc_304 N_B1_c_327_n N_A_511_297#_c_800_n 0.0112654f $X=5.315 $Y=1.41 $X2=0 $Y2=0
cc_305 N_B1_c_328_n N_A_511_297#_c_800_n 0.0112018f $X=5.785 $Y=1.41 $X2=0 $Y2=0
cc_306 N_B1_c_325_n N_VPWR_c_892_n 0.00429453f $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_307 N_B1_c_326_n N_VPWR_c_892_n 0.00429453f $X=4.845 $Y=1.41 $X2=0 $Y2=0
cc_308 N_B1_c_327_n N_VPWR_c_892_n 0.00429453f $X=5.315 $Y=1.41 $X2=0 $Y2=0
cc_309 N_B1_c_328_n N_VPWR_c_892_n 0.00429453f $X=5.785 $Y=1.41 $X2=0 $Y2=0
cc_310 N_B1_c_325_n N_VPWR_c_889_n 0.00609118f $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_311 N_B1_c_326_n N_VPWR_c_889_n 0.00606499f $X=4.845 $Y=1.41 $X2=0 $Y2=0
cc_312 N_B1_c_327_n N_VPWR_c_889_n 0.00606499f $X=5.315 $Y=1.41 $X2=0 $Y2=0
cc_313 N_B1_c_328_n N_VPWR_c_889_n 0.00609118f $X=5.785 $Y=1.41 $X2=0 $Y2=0
cc_314 N_B1_c_319_n N_VGND_c_1011_n 0.00357877f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_315 N_B1_c_320_n N_VGND_c_1011_n 0.00357877f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_316 N_B1_c_321_n N_VGND_c_1011_n 0.00357877f $X=5.29 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B1_c_322_n N_VGND_c_1011_n 0.00357877f $X=5.81 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B1_c_319_n N_VGND_c_1017_n 0.00668309f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_319 N_B1_c_320_n N_VGND_c_1017_n 0.00548399f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_320 N_B1_c_321_n N_VGND_c_1017_n 0.00560377f $X=5.29 $Y=0.995 $X2=0 $Y2=0
cc_321 N_B1_c_322_n N_VGND_c_1017_n 0.00562222f $X=5.81 $Y=0.995 $X2=0 $Y2=0
cc_322 N_B1_c_319_n N_A_503_47#_c_1143_n 0.00931157f $X=4.35 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_B1_c_320_n N_A_503_47#_c_1143_n 0.00931157f $X=4.82 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_B1_c_321_n N_A_503_47#_c_1143_n 0.00964761f $X=5.29 $Y=0.995 $X2=0
+ $Y2=0
cc_325 N_B1_c_322_n N_A_503_47#_c_1143_n 0.00964761f $X=5.81 $Y=0.995 $X2=0
+ $Y2=0
cc_326 N_A2_c_386_n N_A1_c_507_n 0.0260114f $X=6.8 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_327 N_A2_c_385_n N_A1_c_513_n 0.0368713f $X=6.775 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A2_c_399_n N_A1_c_513_n 0.0112841f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_329 N_A2_c_391_n N_A1_c_513_n 0.00101445f $X=6.75 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A2_c_399_n N_A1_c_514_n 0.011867f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_331 N_A2_c_399_n N_A1_c_515_n 0.01191f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_332 N_A2_c_396_n N_A1_c_516_n 0.0362875f $X=9.125 $Y=1.41 $X2=0 $Y2=0
cc_333 N_A2_c_399_n N_A1_c_516_n 0.011867f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_334 N_A2_c_390_n N_A1_c_516_n 6.69584e-19 $X=9.05 $Y=1.445 $X2=0 $Y2=0
cc_335 N_A2_c_387_n N_A1_c_510_n 0.0167003f $X=9.1 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A2_c_385_n N_A1_c_511_n 2.32333e-19 $X=6.775 $Y=1.41 $X2=0 $Y2=0
cc_337 N_A2_c_399_n N_A1_c_511_n 0.113835f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_338 N_A2_c_391_n N_A1_c_511_n 0.0160817f $X=6.75 $Y=1.16 $X2=0 $Y2=0
cc_339 N_A2_c_392_n N_A1_c_511_n 0.0150453f $X=9.135 $Y=1.175 $X2=0 $Y2=0
cc_340 N_A2_c_394_n N_A1_c_511_n 2.24197e-19 $X=10.04 $Y=1.202 $X2=0 $Y2=0
cc_341 N_A2_c_385_n N_A1_c_512_n 0.0263635f $X=6.775 $Y=1.41 $X2=0 $Y2=0
cc_342 N_A2_c_399_n N_A1_c_512_n 0.0231495f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_343 N_A2_c_390_n N_A1_c_512_n 0.00271099f $X=9.05 $Y=1.445 $X2=0 $Y2=0
cc_344 N_A2_c_391_n N_A1_c_512_n 0.00395386f $X=6.75 $Y=1.16 $X2=0 $Y2=0
cc_345 N_A2_c_392_n N_A1_c_512_n 8.29323e-19 $X=9.135 $Y=1.175 $X2=0 $Y2=0
cc_346 N_A2_c_394_n N_A1_c_512_n 0.0167003f $X=10.04 $Y=1.202 $X2=0 $Y2=0
cc_347 N_A2_c_386_n N_Y_c_654_n 3.06774e-19 $X=6.8 $Y=0.995 $X2=0 $Y2=0
cc_348 N_A2_c_385_n N_Y_c_655_n 0.00437142f $X=6.775 $Y=1.41 $X2=0 $Y2=0
cc_349 N_A2_c_386_n N_Y_c_655_n 0.011749f $X=6.8 $Y=0.995 $X2=0 $Y2=0
cc_350 N_A2_c_391_n N_Y_c_655_n 0.0293248f $X=6.75 $Y=1.16 $X2=0 $Y2=0
cc_351 N_A2_c_386_n N_Y_c_656_n 0.00138626f $X=6.8 $Y=0.995 $X2=0 $Y2=0
cc_352 N_A2_c_399_n N_Y_c_656_n 0.00576346f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_353 N_A2_c_391_n N_A_511_297#_M1034_d 0.00161602f $X=6.75 $Y=1.16 $X2=0 $Y2=0
cc_354 N_A2_c_399_n N_A_511_297#_M1000_d 0.00187547f $X=8.965 $Y=1.53 $X2=0
+ $Y2=0
cc_355 N_A2_c_399_n N_A_511_297#_M1031_d 0.00187547f $X=8.965 $Y=1.53 $X2=0
+ $Y2=0
cc_356 N_A2_c_391_n N_A_511_297#_c_805_n 0.00372315f $X=6.75 $Y=1.16 $X2=0 $Y2=0
cc_357 N_A2_c_385_n N_A_511_297#_c_814_n 0.0140027f $X=6.775 $Y=1.41 $X2=0 $Y2=0
cc_358 N_A2_c_396_n N_A_511_297#_c_814_n 0.0146399f $X=9.125 $Y=1.41 $X2=0 $Y2=0
cc_359 N_A2_c_399_n N_A_511_297#_c_814_n 0.120813f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_360 N_A2_c_391_n N_A_511_297#_c_814_n 0.0172816f $X=6.75 $Y=1.16 $X2=0 $Y2=0
cc_361 N_A2_c_393_n N_A_511_297#_c_814_n 0.00313515f $X=9.97 $Y=1.16 $X2=0 $Y2=0
cc_362 N_A2_c_396_n N_A_511_297#_c_819_n 0.00358083f $X=9.125 $Y=1.41 $X2=0
+ $Y2=0
cc_363 N_A2_c_397_n N_A_511_297#_c_819_n 0.00447126f $X=9.595 $Y=1.41 $X2=0
+ $Y2=0
cc_364 N_A2_c_398_n N_A_511_297#_c_819_n 4.63712e-19 $X=10.065 $Y=1.41 $X2=0
+ $Y2=0
cc_365 N_A2_c_397_n N_A_511_297#_c_795_n 0.0137916f $X=9.595 $Y=1.41 $X2=0 $Y2=0
cc_366 N_A2_c_398_n N_A_511_297#_c_795_n 0.0185973f $X=10.065 $Y=1.41 $X2=0
+ $Y2=0
cc_367 N_A2_c_393_n N_A_511_297#_c_795_n 0.0647834f $X=9.97 $Y=1.16 $X2=0 $Y2=0
cc_368 N_A2_c_394_n N_A_511_297#_c_795_n 0.00895735f $X=10.04 $Y=1.202 $X2=0
+ $Y2=0
cc_369 N_A2_c_396_n N_A_511_297#_c_796_n 0.00134335f $X=9.125 $Y=1.41 $X2=0
+ $Y2=0
cc_370 N_A2_c_397_n N_A_511_297#_c_796_n 0.00190955f $X=9.595 $Y=1.41 $X2=0
+ $Y2=0
cc_371 N_A2_c_399_n N_A_511_297#_c_796_n 0.0122348f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_372 N_A2_c_393_n N_A_511_297#_c_796_n 0.0137036f $X=9.97 $Y=1.16 $X2=0 $Y2=0
cc_373 N_A2_c_394_n N_A_511_297#_c_796_n 0.00415172f $X=10.04 $Y=1.202 $X2=0
+ $Y2=0
cc_374 N_A2_c_397_n N_A_511_297#_c_831_n 0.00358587f $X=9.595 $Y=1.41 $X2=0
+ $Y2=0
cc_375 N_A2_c_393_n N_A_511_297#_c_831_n 0.00272072f $X=9.97 $Y=1.16 $X2=0 $Y2=0
cc_376 N_A2_c_394_n N_A_511_297#_c_831_n 0.00157245f $X=10.04 $Y=1.202 $X2=0
+ $Y2=0
cc_377 N_A2_c_399_n N_VPWR_M1005_d 0.00172342f $X=8.965 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_378 N_A2_c_391_n N_VPWR_M1005_d 7.76441e-19 $X=6.75 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_379 N_A2_c_399_n N_VPWR_M1019_s 0.00187547f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_380 N_A2_c_399_n N_VPWR_M1035_s 0.00186949f $X=8.965 $Y=1.53 $X2=0 $Y2=0
cc_381 N_A2_c_397_n N_VPWR_c_890_n 0.00438957f $X=9.595 $Y=1.41 $X2=0 $Y2=0
cc_382 N_A2_c_398_n N_VPWR_c_890_n 0.00571916f $X=10.065 $Y=1.41 $X2=0 $Y2=0
cc_383 N_A2_c_385_n N_VPWR_c_891_n 0.00931192f $X=6.775 $Y=1.41 $X2=0 $Y2=0
cc_384 N_A2_c_385_n N_VPWR_c_892_n 0.00401422f $X=6.775 $Y=1.41 $X2=0 $Y2=0
cc_385 N_A2_c_396_n N_VPWR_c_893_n 0.00372695f $X=9.125 $Y=1.41 $X2=0 $Y2=0
cc_386 N_A2_c_397_n N_VPWR_c_893_n 0.00681844f $X=9.595 $Y=1.41 $X2=0 $Y2=0
cc_387 N_A2_c_398_n N_VPWR_c_896_n 0.00702461f $X=10.065 $Y=1.41 $X2=0 $Y2=0
cc_388 N_A2_c_385_n N_VPWR_c_889_n 0.00478117f $X=6.775 $Y=1.41 $X2=0 $Y2=0
cc_389 N_A2_c_396_n N_VPWR_c_889_n 0.00434988f $X=9.125 $Y=1.41 $X2=0 $Y2=0
cc_390 N_A2_c_397_n N_VPWR_c_889_n 0.0118965f $X=9.595 $Y=1.41 $X2=0 $Y2=0
cc_391 N_A2_c_398_n N_VPWR_c_889_n 0.0135527f $X=10.065 $Y=1.41 $X2=0 $Y2=0
cc_392 N_A2_c_396_n N_VPWR_c_898_n 0.00912658f $X=9.125 $Y=1.41 $X2=0 $Y2=0
cc_393 N_A2_c_397_n N_VPWR_c_898_n 5.82546e-19 $X=9.595 $Y=1.41 $X2=0 $Y2=0
cc_394 N_A2_c_386_n N_VGND_c_1003_n 0.00497791f $X=6.8 $Y=0.995 $X2=0 $Y2=0
cc_395 N_A2_c_387_n N_VGND_c_1004_n 0.00378935f $X=9.1 $Y=0.995 $X2=0 $Y2=0
cc_396 N_A2_c_388_n N_VGND_c_1004_n 0.00276126f $X=9.57 $Y=0.995 $X2=0 $Y2=0
cc_397 N_A2_c_389_n N_VGND_c_1006_n 0.00482457f $X=10.04 $Y=0.995 $X2=0 $Y2=0
cc_398 N_A2_c_393_n N_VGND_c_1006_n 0.014178f $X=9.97 $Y=1.16 $X2=0 $Y2=0
cc_399 N_A2_c_394_n N_VGND_c_1006_n 0.00112974f $X=10.04 $Y=1.202 $X2=0 $Y2=0
cc_400 N_A2_c_386_n N_VGND_c_1013_n 0.00395831f $X=6.8 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A2_c_387_n N_VGND_c_1013_n 0.00421816f $X=9.1 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A2_c_388_n N_VGND_c_1015_n 0.00423334f $X=9.57 $Y=0.995 $X2=0 $Y2=0
cc_403 N_A2_c_389_n N_VGND_c_1015_n 0.00541359f $X=10.04 $Y=0.995 $X2=0 $Y2=0
cc_404 N_A2_c_386_n N_VGND_c_1017_n 0.0058621f $X=6.8 $Y=0.995 $X2=0 $Y2=0
cc_405 N_A2_c_387_n N_VGND_c_1017_n 0.00600232f $X=9.1 $Y=0.995 $X2=0 $Y2=0
cc_406 N_A2_c_388_n N_VGND_c_1017_n 0.00597024f $X=9.57 $Y=0.995 $X2=0 $Y2=0
cc_407 N_A2_c_389_n N_VGND_c_1017_n 0.0106434f $X=10.04 $Y=0.995 $X2=0 $Y2=0
cc_408 N_A2_c_386_n N_A_1375_47#_c_1178_n 0.00509899f $X=6.8 $Y=0.995 $X2=0
+ $Y2=0
cc_409 N_A2_c_387_n N_A_1375_47#_c_1179_n 0.00282739f $X=9.1 $Y=0.995 $X2=0
+ $Y2=0
cc_410 N_A2_c_387_n N_A_1375_47#_c_1176_n 0.00513774f $X=9.1 $Y=0.995 $X2=0
+ $Y2=0
cc_411 N_A2_c_388_n N_A_1375_47#_c_1176_n 4.74935e-19 $X=9.57 $Y=0.995 $X2=0
+ $Y2=0
cc_412 N_A2_c_399_n N_A_1375_47#_c_1176_n 0.00600976f $X=8.965 $Y=1.53 $X2=0
+ $Y2=0
cc_413 N_A2_c_392_n N_A_1375_47#_c_1176_n 0.00799416f $X=9.135 $Y=1.175 $X2=0
+ $Y2=0
cc_414 N_A2_c_387_n N_A_1375_47#_c_1177_n 0.00901419f $X=9.1 $Y=0.995 $X2=0
+ $Y2=0
cc_415 N_A2_c_388_n N_A_1375_47#_c_1177_n 0.0101253f $X=9.57 $Y=0.995 $X2=0
+ $Y2=0
cc_416 N_A2_c_389_n N_A_1375_47#_c_1177_n 0.00266157f $X=10.04 $Y=0.995 $X2=0
+ $Y2=0
cc_417 N_A2_c_392_n N_A_1375_47#_c_1177_n 0.00596758f $X=9.135 $Y=1.175 $X2=0
+ $Y2=0
cc_418 N_A2_c_393_n N_A_1375_47#_c_1177_n 0.0648321f $X=9.97 $Y=1.16 $X2=0 $Y2=0
cc_419 N_A2_c_394_n N_A_1375_47#_c_1177_n 0.00703846f $X=10.04 $Y=1.202 $X2=0
+ $Y2=0
cc_420 N_A2_c_387_n N_A_1375_47#_c_1190_n 5.24597e-19 $X=9.1 $Y=0.995 $X2=0
+ $Y2=0
cc_421 N_A2_c_388_n N_A_1375_47#_c_1190_n 0.00651696f $X=9.57 $Y=0.995 $X2=0
+ $Y2=0
cc_422 N_A2_c_389_n N_A_1375_47#_c_1190_n 0.00539651f $X=10.04 $Y=0.995 $X2=0
+ $Y2=0
cc_423 N_A1_c_507_n N_Y_c_726_n 0.00864619f $X=7.22 $Y=0.995 $X2=0 $Y2=0
cc_424 N_A1_c_508_n N_Y_c_726_n 0.00929111f $X=7.69 $Y=0.995 $X2=0 $Y2=0
cc_425 N_A1_c_509_n N_Y_c_726_n 0.00929111f $X=8.16 $Y=0.995 $X2=0 $Y2=0
cc_426 N_A1_c_511_n N_Y_c_726_n 0.065269f $X=8.09 $Y=1.16 $X2=0 $Y2=0
cc_427 N_A1_c_512_n N_Y_c_726_n 0.0109421f $X=8.655 $Y=1.202 $X2=0 $Y2=0
cc_428 N_A1_c_507_n N_Y_c_656_n 8.89068e-19 $X=7.22 $Y=0.995 $X2=0 $Y2=0
cc_429 N_A1_c_513_n N_A_511_297#_c_814_n 0.0124275f $X=7.245 $Y=1.41 $X2=0 $Y2=0
cc_430 N_A1_c_514_n N_A_511_297#_c_814_n 0.0124936f $X=7.715 $Y=1.41 $X2=0 $Y2=0
cc_431 N_A1_c_515_n N_A_511_297#_c_814_n 0.0124936f $X=8.185 $Y=1.41 $X2=0 $Y2=0
cc_432 N_A1_c_516_n N_A_511_297#_c_814_n 0.0124275f $X=8.655 $Y=1.41 $X2=0 $Y2=0
cc_433 N_A1_c_513_n N_VPWR_c_895_n 0.0190585f $X=7.245 $Y=1.41 $X2=0 $Y2=0
cc_434 N_A1_c_514_n N_VPWR_c_895_n 0.0190916f $X=7.715 $Y=1.41 $X2=0 $Y2=0
cc_435 N_A1_c_515_n N_VPWR_c_895_n 0.0190916f $X=8.185 $Y=1.41 $X2=0 $Y2=0
cc_436 N_A1_c_516_n N_VPWR_c_895_n 0.0190585f $X=8.655 $Y=1.41 $X2=0 $Y2=0
cc_437 N_A1_c_507_n N_VGND_c_1013_n 0.00357877f $X=7.22 $Y=0.995 $X2=0 $Y2=0
cc_438 N_A1_c_508_n N_VGND_c_1013_n 0.00357877f $X=7.69 $Y=0.995 $X2=0 $Y2=0
cc_439 N_A1_c_509_n N_VGND_c_1013_n 0.00357877f $X=8.16 $Y=0.995 $X2=0 $Y2=0
cc_440 N_A1_c_510_n N_VGND_c_1013_n 0.00357877f $X=8.68 $Y=0.995 $X2=0 $Y2=0
cc_441 N_A1_c_507_n N_VGND_c_1017_n 0.00538422f $X=7.22 $Y=0.995 $X2=0 $Y2=0
cc_442 N_A1_c_508_n N_VGND_c_1017_n 0.00548399f $X=7.69 $Y=0.995 $X2=0 $Y2=0
cc_443 N_A1_c_509_n N_VGND_c_1017_n 0.00560377f $X=8.16 $Y=0.995 $X2=0 $Y2=0
cc_444 N_A1_c_510_n N_VGND_c_1017_n 0.005504f $X=8.68 $Y=0.995 $X2=0 $Y2=0
cc_445 N_A1_c_507_n N_A_1375_47#_c_1178_n 0.00931157f $X=7.22 $Y=0.995 $X2=0
+ $Y2=0
cc_446 N_A1_c_508_n N_A_1375_47#_c_1178_n 0.00931157f $X=7.69 $Y=0.995 $X2=0
+ $Y2=0
cc_447 N_A1_c_509_n N_A_1375_47#_c_1178_n 0.00964761f $X=8.16 $Y=0.995 $X2=0
+ $Y2=0
cc_448 N_A1_c_510_n N_A_1375_47#_c_1178_n 0.0117007f $X=8.68 $Y=0.995 $X2=0
+ $Y2=0
cc_449 N_A1_c_511_n N_A_1375_47#_c_1178_n 0.00393303f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_450 N_A1_c_510_n N_A_1375_47#_c_1176_n 6.06509e-19 $X=8.68 $Y=0.995 $X2=0
+ $Y2=0
cc_451 N_A_27_297#_c_576_n N_Y_M1003_d 0.00352392f $X=1.095 $Y=2.38 $X2=0 $Y2=0
cc_452 N_A_27_297#_c_578_n N_Y_M1016_d 0.00352392f $X=2.075 $Y=2.38 $X2=0 $Y2=0
cc_453 N_A_27_297#_c_576_n N_Y_c_734_n 0.0134104f $X=1.095 $Y=2.38 $X2=0 $Y2=0
cc_454 N_A_27_297#_M1010_s N_Y_c_657_n 0.00187091f $X=1.075 $Y=1.485 $X2=0 $Y2=0
cc_455 N_A_27_297#_c_606_p N_Y_c_657_n 0.0143191f $X=1.22 $Y=1.96 $X2=0 $Y2=0
cc_456 N_A_27_297#_c_568_n N_Y_c_658_n 0.00286441f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_457 N_A_27_297#_c_578_n N_Y_c_738_n 0.0134104f $X=2.075 $Y=2.38 $X2=0 $Y2=0
cc_458 N_A_27_297#_c_571_n N_Y_c_651_n 0.0740177f $X=3.035 $Y=1.53 $X2=0 $Y2=0
cc_459 N_A_27_297#_c_572_n N_Y_c_651_n 0.0211976f $X=2.325 $Y=1.53 $X2=0 $Y2=0
cc_460 N_A_27_297#_c_592_n N_Y_c_651_n 0.00651545f $X=6.02 $Y=1.96 $X2=0 $Y2=0
cc_461 N_A_27_297#_c_572_n N_Y_c_660_n 0.0122341f $X=2.325 $Y=1.53 $X2=0 $Y2=0
cc_462 N_A_27_297#_c_571_n N_A_511_297#_M1014_d 0.00411964f $X=3.035 $Y=1.53
+ $X2=-0.19 $Y2=1.305
cc_463 N_A_27_297#_c_592_n N_A_511_297#_M1018_d 0.00463783f $X=6.02 $Y=1.96
+ $X2=0 $Y2=0
cc_464 N_A_27_297#_c_592_n N_A_511_297#_M1004_s 0.0036976f $X=6.02 $Y=1.96 $X2=0
+ $Y2=0
cc_465 N_A_27_297#_c_592_n N_A_511_297#_M1026_s 0.0036976f $X=6.02 $Y=1.96 $X2=0
+ $Y2=0
cc_466 N_A_27_297#_c_569_n N_A_511_297#_c_842_n 0.0121718f $X=2.2 $Y=2.295 $X2=0
+ $Y2=0
cc_467 N_A_27_297#_c_570_n N_A_511_297#_c_842_n 0.00526703f $X=2.16 $Y=1.63
+ $X2=0 $Y2=0
cc_468 N_A_27_297#_c_570_n N_A_511_297#_c_844_n 0.0256826f $X=2.16 $Y=1.63 $X2=0
+ $Y2=0
cc_469 N_A_27_297#_c_571_n N_A_511_297#_c_844_n 0.019309f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_470 N_A_27_297#_c_590_n N_A_511_297#_c_844_n 0.0138894f $X=3.182 $Y=1.835
+ $X2=0 $Y2=0
cc_471 N_A_27_297#_c_591_n N_A_511_297#_c_844_n 0.00244225f $X=3.2 $Y=1.62 $X2=0
+ $Y2=0
cc_472 N_A_27_297#_M1014_s N_A_511_297#_c_800_n 0.00356605f $X=3.055 $Y=1.485
+ $X2=0 $Y2=0
cc_473 N_A_27_297#_M1030_s N_A_511_297#_c_800_n 0.00357068f $X=3.995 $Y=1.485
+ $X2=0 $Y2=0
cc_474 N_A_27_297#_M1012_d N_A_511_297#_c_800_n 0.00357068f $X=4.935 $Y=1.485
+ $X2=0 $Y2=0
cc_475 N_A_27_297#_M1032_d N_A_511_297#_c_800_n 0.00357068f $X=5.875 $Y=1.485
+ $X2=0 $Y2=0
cc_476 N_A_27_297#_c_571_n N_A_511_297#_c_800_n 0.00395611f $X=3.035 $Y=1.53
+ $X2=0 $Y2=0
cc_477 N_A_27_297#_c_590_n N_A_511_297#_c_800_n 0.0153108f $X=3.182 $Y=1.835
+ $X2=0 $Y2=0
cc_478 N_A_27_297#_c_592_n N_A_511_297#_c_800_n 0.150886f $X=6.02 $Y=1.96 $X2=0
+ $Y2=0
cc_479 N_A_27_297#_c_592_n N_A_511_297#_c_805_n 0.0148798f $X=6.02 $Y=1.96 $X2=0
+ $Y2=0
cc_480 N_A_27_297#_c_567_n N_VPWR_c_892_n 0.0209238f $X=0.247 $Y=2.295 $X2=0
+ $Y2=0
cc_481 N_A_27_297#_c_576_n N_VPWR_c_892_n 0.0386815f $X=1.095 $Y=2.38 $X2=0
+ $Y2=0
cc_482 N_A_27_297#_c_578_n N_VPWR_c_892_n 0.0400924f $X=2.075 $Y=2.38 $X2=0
+ $Y2=0
cc_483 N_A_27_297#_c_569_n N_VPWR_c_892_n 0.0176351f $X=2.2 $Y=2.295 $X2=0 $Y2=0
cc_484 N_A_27_297#_c_635_p N_VPWR_c_892_n 0.015002f $X=1.22 $Y=2.38 $X2=0 $Y2=0
cc_485 N_A_27_297#_M1003_s N_VPWR_c_889_n 0.00233915f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_486 N_A_27_297#_M1010_s N_VPWR_c_889_n 0.00231264f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_487 N_A_27_297#_M1028_s N_VPWR_c_889_n 0.00217523f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_488 N_A_27_297#_M1014_s N_VPWR_c_889_n 0.00232895f $X=3.055 $Y=1.485 $X2=0
+ $Y2=0
cc_489 N_A_27_297#_M1030_s N_VPWR_c_889_n 0.00232895f $X=3.995 $Y=1.485 $X2=0
+ $Y2=0
cc_490 N_A_27_297#_M1012_d N_VPWR_c_889_n 0.00232895f $X=4.935 $Y=1.485 $X2=0
+ $Y2=0
cc_491 N_A_27_297#_M1032_d N_VPWR_c_889_n 0.00232895f $X=5.875 $Y=1.485 $X2=0
+ $Y2=0
cc_492 N_A_27_297#_c_567_n N_VPWR_c_889_n 0.012126f $X=0.247 $Y=2.295 $X2=0
+ $Y2=0
cc_493 N_A_27_297#_c_576_n N_VPWR_c_889_n 0.0239144f $X=1.095 $Y=2.38 $X2=0
+ $Y2=0
cc_494 N_A_27_297#_c_578_n N_VPWR_c_889_n 0.0253962f $X=2.075 $Y=2.38 $X2=0
+ $Y2=0
cc_495 N_A_27_297#_c_569_n N_VPWR_c_889_n 0.00962794f $X=2.2 $Y=2.295 $X2=0
+ $Y2=0
cc_496 N_A_27_297#_c_635_p N_VPWR_c_889_n 0.00962794f $X=1.22 $Y=2.38 $X2=0
+ $Y2=0
cc_497 N_Y_M1003_d N_VPWR_c_889_n 0.00232895f $X=0.605 $Y=1.485 $X2=0 $Y2=0
cc_498 N_Y_M1016_d N_VPWR_c_889_n 0.00232895f $X=1.545 $Y=1.485 $X2=0 $Y2=0
cc_499 N_Y_c_648_n N_VGND_M1020_s 0.00251047f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_500 N_Y_c_655_n N_VGND_M1036_s 0.00353543f $X=6.96 $Y=0.775 $X2=0 $Y2=0
cc_501 N_Y_c_661_n N_VGND_c_998_n 0.0360647f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_502 N_Y_c_649_n N_VGND_c_998_n 0.0137446f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_503 N_Y_c_661_n N_VGND_c_999_n 0.023074f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_504 N_Y_c_648_n N_VGND_c_999_n 0.00254521f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_505 N_Y_c_648_n N_VGND_c_1000_n 0.0127273f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_506 N_Y_c_676_n N_VGND_c_1000_n 0.0223967f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_507 N_Y_c_650_n N_VGND_c_1002_n 0.00139066f $X=1.755 $Y=1.095 $X2=0 $Y2=0
cc_508 N_Y_c_651_n N_VGND_c_1002_n 0.0144144f $X=3.375 $Y=1.185 $X2=0 $Y2=0
cc_509 N_Y_c_653_n N_VGND_c_1002_n 0.00148154f $X=1.665 $Y=0.815 $X2=0 $Y2=0
cc_510 N_Y_c_655_n N_VGND_c_1003_n 0.0125492f $X=6.96 $Y=0.775 $X2=0 $Y2=0
cc_511 N_Y_c_648_n N_VGND_c_1007_n 0.00199443f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_512 N_Y_c_676_n N_VGND_c_1007_n 0.0231119f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_513 N_Y_c_652_n N_VGND_c_1009_n 0.00838459f $X=3.485 $Y=1.095 $X2=0 $Y2=0
cc_514 N_Y_c_700_n N_VGND_c_1009_n 0.0152956f $X=3.595 $Y=0.732 $X2=0 $Y2=0
cc_515 N_Y_c_651_n N_VGND_c_1010_n 0.0711431f $X=3.375 $Y=1.185 $X2=0 $Y2=0
cc_516 N_Y_c_654_n N_VGND_c_1011_n 0.00142251f $X=6.28 $Y=0.775 $X2=0 $Y2=0
cc_517 N_Y_c_655_n N_VGND_c_1011_n 0.00201105f $X=6.96 $Y=0.775 $X2=0 $Y2=0
cc_518 N_Y_c_655_n N_VGND_c_1013_n 0.00195107f $X=6.96 $Y=0.775 $X2=0 $Y2=0
cc_519 N_Y_M1007_d N_VGND_c_1017_n 0.00263993f $X=0.615 $Y=0.235 $X2=0 $Y2=0
cc_520 N_Y_M1024_d N_VGND_c_1017_n 0.00324782f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_521 N_Y_M1021_s N_VGND_c_1017_n 0.00256987f $X=4.425 $Y=0.235 $X2=0 $Y2=0
cc_522 N_Y_M1029_s N_VGND_c_1017_n 0.00297142f $X=5.365 $Y=0.235 $X2=0 $Y2=0
cc_523 N_Y_M1002_s N_VGND_c_1017_n 0.00256987f $X=7.295 $Y=0.235 $X2=0 $Y2=0
cc_524 N_Y_M1017_s N_VGND_c_1017_n 0.00297142f $X=8.235 $Y=0.235 $X2=0 $Y2=0
cc_525 N_Y_c_661_n N_VGND_c_1017_n 0.0141066f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_526 N_Y_c_648_n N_VGND_c_1017_n 0.00977515f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_527 N_Y_c_676_n N_VGND_c_1017_n 0.0141157f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_528 N_Y_c_702_n N_VGND_c_1017_n 0.00705923f $X=6.11 $Y=0.775 $X2=0 $Y2=0
cc_529 N_Y_c_655_n N_VGND_c_1017_n 0.00932591f $X=6.96 $Y=0.775 $X2=0 $Y2=0
cc_530 N_Y_c_652_n N_A_503_47#_M1027_d 0.00117859f $X=3.485 $Y=1.095 $X2=0 $Y2=0
cc_531 N_Y_c_700_n N_A_503_47#_M1027_d 8.85226e-19 $X=3.595 $Y=0.732 $X2=0 $Y2=0
cc_532 N_Y_c_702_n N_A_503_47#_M1027_d 0.0174347f $X=6.11 $Y=0.775 $X2=0 $Y2=0
cc_533 N_Y_c_702_n N_A_503_47#_M1022_d 0.00401748f $X=6.11 $Y=0.775 $X2=0 $Y2=0
cc_534 N_Y_c_702_n N_A_503_47#_M1038_d 0.00472948f $X=6.11 $Y=0.775 $X2=0 $Y2=0
cc_535 N_Y_c_654_n N_A_503_47#_M1038_d 0.00132244f $X=6.28 $Y=0.775 $X2=0 $Y2=0
cc_536 N_Y_c_651_n N_A_503_47#_c_1141_n 9.37998e-19 $X=3.375 $Y=1.185 $X2=0
+ $Y2=0
cc_537 N_Y_c_700_n N_A_503_47#_c_1141_n 0.012237f $X=3.595 $Y=0.732 $X2=0 $Y2=0
cc_538 N_Y_M1021_s N_A_503_47#_c_1143_n 0.00400389f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_539 N_Y_M1029_s N_A_503_47#_c_1143_n 0.00507817f $X=5.365 $Y=0.235 $X2=0
+ $Y2=0
cc_540 N_Y_c_702_n N_A_503_47#_c_1143_n 0.145037f $X=6.11 $Y=0.775 $X2=0 $Y2=0
cc_541 N_Y_c_651_n N_A_503_47#_c_1145_n 0.00228037f $X=3.375 $Y=1.185 $X2=0
+ $Y2=0
cc_542 N_Y_c_655_n N_A_1375_47#_M1006_d 3.3779e-19 $X=6.96 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_543 N_Y_c_656_n N_A_1375_47#_M1006_d 0.00255149f $X=7.13 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_544 N_Y_c_726_n N_A_1375_47#_M1011_d 0.00434237f $X=8.42 $Y=0.73 $X2=0 $Y2=0
cc_545 N_Y_M1002_s N_A_1375_47#_c_1178_n 0.00400389f $X=7.295 $Y=0.235 $X2=0
+ $Y2=0
cc_546 N_Y_M1017_s N_A_1375_47#_c_1178_n 0.00507817f $X=8.235 $Y=0.235 $X2=0
+ $Y2=0
cc_547 N_Y_c_655_n N_A_1375_47#_c_1178_n 0.00493364f $X=6.96 $Y=0.775 $X2=0
+ $Y2=0
cc_548 N_Y_c_656_n N_A_1375_47#_c_1178_n 0.0859508f $X=7.13 $Y=0.775 $X2=0 $Y2=0
cc_549 N_A_511_297#_c_814_n N_VPWR_M1005_d 0.00370129f $X=9.275 $Y=1.915
+ $X2=-0.19 $Y2=1.305
cc_550 N_A_511_297#_c_814_n N_VPWR_M1019_s 0.00350737f $X=9.275 $Y=1.915 $X2=0
+ $Y2=0
cc_551 N_A_511_297#_c_814_n N_VPWR_M1035_s 0.0037405f $X=9.275 $Y=1.915 $X2=0
+ $Y2=0
cc_552 N_A_511_297#_c_795_n N_VPWR_M1013_d 0.00182924f $X=10.175 $Y=1.53 $X2=0
+ $Y2=0
cc_553 N_A_511_297#_c_860_p N_VPWR_c_890_n 0.0200543f $X=9.36 $Y=2.3 $X2=0 $Y2=0
cc_554 N_A_511_297#_c_795_n N_VPWR_c_890_n 0.0130962f $X=10.175 $Y=1.53 $X2=0
+ $Y2=0
cc_555 N_A_511_297#_c_831_n N_VPWR_c_890_n 0.0160874f $X=9.36 $Y=1.96 $X2=0
+ $Y2=0
cc_556 N_A_511_297#_c_814_n N_VPWR_c_891_n 0.12896f $X=9.275 $Y=1.915 $X2=0
+ $Y2=0
cc_557 N_A_511_297#_c_842_n N_VPWR_c_892_n 0.0175612f $X=2.69 $Y=2.215 $X2=0
+ $Y2=0
cc_558 N_A_511_297#_c_800_n N_VPWR_c_892_n 0.203204f $X=6.405 $Y=2.34 $X2=0
+ $Y2=0
cc_559 N_A_511_297#_c_866_p N_VPWR_c_892_n 0.0166395f $X=6.53 $Y=2.215 $X2=0
+ $Y2=0
cc_560 N_A_511_297#_c_814_n N_VPWR_c_892_n 0.00239818f $X=9.275 $Y=1.915 $X2=0
+ $Y2=0
cc_561 N_A_511_297#_c_814_n N_VPWR_c_893_n 0.00250917f $X=9.275 $Y=1.915 $X2=0
+ $Y2=0
cc_562 N_A_511_297#_c_860_p N_VPWR_c_893_n 0.0118139f $X=9.36 $Y=2.3 $X2=0 $Y2=0
cc_563 N_A_511_297#_c_831_n N_VPWR_c_893_n 8.748e-19 $X=9.36 $Y=1.96 $X2=0 $Y2=0
cc_564 N_A_511_297#_M1000_d N_VPWR_c_895_n 0.00194857f $X=7.335 $Y=1.485 $X2=0
+ $Y2=0
cc_565 N_A_511_297#_M1031_d N_VPWR_c_895_n 0.00194857f $X=8.275 $Y=1.485 $X2=0
+ $Y2=0
cc_566 N_A_511_297#_c_873_p N_VPWR_c_896_n 0.0161853f $X=10.3 $Y=1.82 $X2=0
+ $Y2=0
cc_567 N_A_511_297#_M1014_d N_VPWR_c_889_n 0.00293228f $X=2.555 $Y=1.485 $X2=0
+ $Y2=0
cc_568 N_A_511_297#_M1018_d N_VPWR_c_889_n 0.00231289f $X=3.525 $Y=1.485 $X2=0
+ $Y2=0
cc_569 N_A_511_297#_M1004_s N_VPWR_c_889_n 0.00231289f $X=4.465 $Y=1.485 $X2=0
+ $Y2=0
cc_570 N_A_511_297#_M1026_s N_VPWR_c_889_n 0.00231289f $X=5.405 $Y=1.485 $X2=0
+ $Y2=0
cc_571 N_A_511_297#_M1034_d N_VPWR_c_889_n 0.00283685f $X=6.345 $Y=1.485 $X2=0
+ $Y2=0
cc_572 N_A_511_297#_M1008_s N_VPWR_c_889_n 0.00279492f $X=9.215 $Y=1.485 $X2=0
+ $Y2=0
cc_573 N_A_511_297#_M1023_s N_VPWR_c_889_n 0.00380522f $X=10.155 $Y=1.485 $X2=0
+ $Y2=0
cc_574 N_A_511_297#_c_842_n N_VPWR_c_889_n 0.00962421f $X=2.69 $Y=2.215 $X2=0
+ $Y2=0
cc_575 N_A_511_297#_c_800_n N_VPWR_c_889_n 0.127685f $X=6.405 $Y=2.34 $X2=0
+ $Y2=0
cc_576 N_A_511_297#_c_866_p N_VPWR_c_889_n 0.00962794f $X=6.53 $Y=2.215 $X2=0
+ $Y2=0
cc_577 N_A_511_297#_c_814_n N_VPWR_c_889_n 0.0179807f $X=9.275 $Y=1.915 $X2=0
+ $Y2=0
cc_578 N_A_511_297#_c_860_p N_VPWR_c_889_n 0.00646998f $X=9.36 $Y=2.3 $X2=0
+ $Y2=0
cc_579 N_A_511_297#_c_873_p N_VPWR_c_889_n 0.00955092f $X=10.3 $Y=1.82 $X2=0
+ $Y2=0
cc_580 N_A_511_297#_c_831_n N_VPWR_c_889_n 0.00216775f $X=9.36 $Y=1.96 $X2=0
+ $Y2=0
cc_581 N_A_511_297#_c_860_p N_VPWR_c_898_n 0.0179477f $X=9.36 $Y=2.3 $X2=0 $Y2=0
cc_582 N_VGND_c_1010_n N_A_503_47#_M1001_d 0.00214831f $X=3.035 $Y=0.76
+ $X2=-0.19 $Y2=-0.24
cc_583 N_VGND_c_1017_n N_A_503_47#_M1001_d 0.00255381f $X=10.35 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_584 N_VGND_c_1017_n N_A_503_47#_M1027_d 0.00664657f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_585 N_VGND_c_1017_n N_A_503_47#_M1022_d 0.00255381f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_586 N_VGND_c_1017_n N_A_503_47#_M1038_d 0.00262586f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_1001_n N_A_503_47#_c_1140_n 0.0155832f $X=2.16 $Y=0.39 $X2=0
+ $Y2=0
cc_588 N_VGND_c_1010_n N_A_503_47#_c_1140_n 0.0220992f $X=3.035 $Y=0.76 $X2=0
+ $Y2=0
cc_589 N_VGND_c_1011_n N_A_503_47#_c_1140_n 0.216556f $X=6.455 $Y=0 $X2=0 $Y2=0
cc_590 N_VGND_c_1017_n N_A_503_47#_c_1140_n 0.13538f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_591 N_VGND_M1015_s N_A_503_47#_c_1145_n 0.00441779f $X=2.985 $Y=0.235 $X2=0
+ $Y2=0
cc_592 N_VGND_c_1009_n N_A_503_47#_c_1145_n 0.0116976f $X=3.12 $Y=0.76 $X2=0
+ $Y2=0
cc_593 N_VGND_c_1010_n N_A_503_47#_c_1145_n 0.0064979f $X=3.035 $Y=0.76 $X2=0
+ $Y2=0
cc_594 N_VGND_c_1017_n N_A_1375_47#_M1006_d 0.00215227f $X=10.35 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_595 N_VGND_c_1017_n N_A_1375_47#_M1011_d 0.00255381f $X=10.35 $Y=0 $X2=0
+ $Y2=0
cc_596 N_VGND_c_1017_n N_A_1375_47#_M1039_d 0.00215206f $X=10.35 $Y=0 $X2=0
+ $Y2=0
cc_597 N_VGND_c_1017_n N_A_1375_47#_M1025_d 0.0025535f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_c_1003_n N_A_1375_47#_c_1178_n 0.0171345f $X=6.54 $Y=0.39 $X2=0
+ $Y2=0
cc_599 N_VGND_c_1013_n N_A_1375_47#_c_1178_n 0.113411f $X=9.275 $Y=0 $X2=0 $Y2=0
cc_600 N_VGND_c_1017_n N_A_1375_47#_c_1178_n 0.0718274f $X=10.35 $Y=0 $X2=0
+ $Y2=0
cc_601 N_VGND_c_1004_n N_A_1375_47#_c_1179_n 0.0141571f $X=9.36 $Y=0.39 $X2=0
+ $Y2=0
cc_602 N_VGND_c_1013_n N_A_1375_47#_c_1179_n 0.0152108f $X=9.275 $Y=0 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1017_n N_A_1375_47#_c_1179_n 0.00940698f $X=10.35 $Y=0 $X2=0
+ $Y2=0
cc_604 N_VGND_c_1004_n N_A_1375_47#_c_1176_n 0.00471242f $X=9.36 $Y=0.39 $X2=0
+ $Y2=0
cc_605 N_VGND_M1009_s N_A_1375_47#_c_1177_n 0.00251047f $X=9.175 $Y=0.235 $X2=0
+ $Y2=0
cc_606 N_VGND_c_1004_n N_A_1375_47#_c_1177_n 0.0127273f $X=9.36 $Y=0.39 $X2=0
+ $Y2=0
cc_607 N_VGND_c_1006_n N_A_1375_47#_c_1177_n 0.00830019f $X=10.25 $Y=0.39 $X2=0
+ $Y2=0
cc_608 N_VGND_c_1013_n N_A_1375_47#_c_1177_n 0.00266636f $X=9.275 $Y=0 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1015_n N_A_1375_47#_c_1177_n 0.00198695f $X=10.165 $Y=0 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1017_n N_A_1375_47#_c_1177_n 0.00972452f $X=10.35 $Y=0 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1015_n N_A_1375_47#_c_1190_n 0.0223596f $X=10.165 $Y=0 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1017_n N_A_1375_47#_c_1190_n 0.0141302f $X=10.35 $Y=0 $X2=0
+ $Y2=0
