* File: sky130_fd_sc_hdll__mux2i_2.pxi.spice
* Created: Thu Aug 27 19:11:08 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%S N_S_c_85_n N_S_M1005_g N_S_c_80_n N_S_M1011_g
+ N_S_c_86_n N_S_M1001_g N_S_c_81_n N_S_M1002_g N_S_c_87_n N_S_M1014_g
+ N_S_c_82_n N_S_M1016_g S S N_S_c_84_n PM_SKY130_FD_SC_HDLL__MUX2I_2%S
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%A_27_47# N_A_27_47#_M1011_s N_A_27_47#_M1005_s
+ N_A_27_47#_c_153_n N_A_27_47#_M1006_g N_A_27_47#_M1008_g N_A_27_47#_c_154_n
+ N_A_27_47#_M1009_g N_A_27_47#_M1012_g N_A_27_47#_c_149_n N_A_27_47#_c_168_n
+ N_A_27_47#_c_156_n N_A_27_47#_c_176_n N_A_27_47#_c_150_n N_A_27_47#_c_157_n
+ N_A_27_47#_c_158_n N_A_27_47#_c_159_n N_A_27_47#_c_179_n N_A_27_47#_c_151_n
+ N_A_27_47#_c_152_n PM_SKY130_FD_SC_HDLL__MUX2I_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%A0 N_A0_c_248_n N_A0_M1004_g N_A0_c_243_n
+ N_A0_M1000_g N_A0_c_249_n N_A0_M1015_g N_A0_c_244_n N_A0_M1003_g A0 A0 A0
+ N_A0_c_246_n N_A0_c_247_n A0 A0 A0 PM_SKY130_FD_SC_HDLL__MUX2I_2%A0
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%A1 N_A1_c_297_n N_A1_M1007_g N_A1_c_301_n
+ N_A1_M1010_g N_A1_c_298_n N_A1_M1017_g N_A1_c_302_n N_A1_M1013_g A1 A1
+ N_A1_c_299_n N_A1_c_300_n PM_SKY130_FD_SC_HDLL__MUX2I_2%A1
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%VPWR N_VPWR_M1005_d N_VPWR_M1014_s
+ N_VPWR_M1009_d N_VPWR_c_341_n N_VPWR_c_342_n VPWR N_VPWR_c_343_n
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_340_n N_VPWR_c_347_n N_VPWR_c_348_n
+ N_VPWR_c_349_n PM_SKY130_FD_SC_HDLL__MUX2I_2%VPWR
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%A_211_297# N_A_211_297#_M1001_d
+ N_A_211_297#_M1004_d N_A_211_297#_c_412_n N_A_211_297#_c_415_n
+ N_A_211_297#_c_416_n N_A_211_297#_c_429_n N_A_211_297#_c_411_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_2%A_211_297#
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%A_399_297# N_A_399_297#_M1006_s
+ N_A_399_297#_M1010_s N_A_399_297#_c_463_n N_A_399_297#_c_460_n
+ N_A_399_297#_c_458_n N_A_399_297#_c_459_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_2%A_399_297#
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%Y N_Y_M1000_d N_Y_M1003_d N_Y_M1017_s
+ N_Y_M1004_s N_Y_M1015_s N_Y_M1013_d N_Y_c_494_n Y Y N_Y_c_498_n Y Y
+ PM_SKY130_FD_SC_HDLL__MUX2I_2%Y
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%VGND N_VGND_M1011_d N_VGND_M1016_s
+ N_VGND_M1012_d N_VGND_c_549_n N_VGND_c_550_n N_VGND_c_551_n N_VGND_c_552_n
+ N_VGND_c_553_n VGND N_VGND_c_554_n N_VGND_c_555_n N_VGND_c_556_n
+ N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_2%VGND
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%A_213_47# N_A_213_47#_M1002_d
+ N_A_213_47#_M1007_d N_A_213_47#_c_623_n N_A_213_47#_c_624_n
+ N_A_213_47#_c_625_n N_A_213_47#_c_626_n N_A_213_47#_c_627_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_2%A_213_47#
x_PM_SKY130_FD_SC_HDLL__MUX2I_2%A_401_47# N_A_401_47#_M1008_s
+ N_A_401_47#_M1000_s N_A_401_47#_c_690_n N_A_401_47#_c_687_n
+ N_A_401_47#_c_688_n N_A_401_47#_c_689_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_2%A_401_47#
cc_1 VNB N_S_c_80_n 0.019229f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_S_c_81_n 0.0169082f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_S_c_82_n 0.0166785f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_4 VNB S 0.00205484f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_5 VNB N_S_c_84_n 0.0611882f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_6 VNB N_A_27_47#_M1008_g 0.018531f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_7 VNB N_A_27_47#_M1012_g 0.0233108f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.765
cc_8 VNB N_A_27_47#_c_149_n 0.027306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_150_n 0.01296f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.85
cc_10 VNB N_A_27_47#_c_151_n 0.00229698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_152_n 0.0353714f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A0_c_243_n 0.0216975f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_13 VNB N_A0_c_244_n 0.0167702f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_14 VNB A0 0.00581408f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_15 VNB N_A0_c_246_n 0.0473559f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.765
cc_16 VNB N_A0_c_247_n 0.0341629f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_17 VNB N_A1_c_297_n 0.016323f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_18 VNB N_A1_c_298_n 0.0201933f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_19 VNB N_A1_c_299_n 0.0560162f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_20 VNB N_A1_c_300_n 0.00328207f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_21 VNB N_VPWR_c_340_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.19
cc_22 VNB N_Y_c_494_n 0.00990813f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.765
cc_23 VNB Y 0.0351475f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_24 VNB N_VGND_c_549_n 0.00275138f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_25 VNB N_VGND_c_550_n 0.0210182f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_26 VNB N_VGND_c_551_n 0.00621771f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_27 VNB N_VGND_c_552_n 0.0193309f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_28 VNB N_VGND_c_553_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_29 VNB N_VGND_c_554_n 0.0154495f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_30 VNB N_VGND_c_555_n 0.0696979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_556_n 0.278986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_557_n 0.00554944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_558_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_559_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_213_47#_c_623_n 0.0186754f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_36 VNB N_A_213_47#_c_624_n 0.00352753f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_37 VNB N_A_213_47#_c_625_n 0.00822332f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_38 VNB N_A_213_47#_c_626_n 0.00310931f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_39 VNB N_A_213_47#_c_627_n 0.00322305f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_40 VNB N_A_401_47#_c_687_n 0.00106438f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_41 VNB N_A_401_47#_c_688_n 0.00120415f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_42 VNB N_A_401_47#_c_689_n 0.0104335f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_43 VPB N_S_c_85_n 0.0187457f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_44 VPB N_S_c_86_n 0.0160781f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_45 VPB N_S_c_87_n 0.0151596f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_46 VPB S 0.00219871f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_47 VPB N_S_c_84_n 0.0333731f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.202
cc_48 VPB N_A_27_47#_c_153_n 0.0162168f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_49 VPB N_A_27_47#_c_154_n 0.0210879f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_50 VPB N_A_27_47#_c_149_n 0.00909759f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_156_n 0.0033713f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_52 VPB N_A_27_47#_c_157_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_158_n 0.0128993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_159_n 0.0169831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_151_n 0.00316123f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_152_n 0.0231139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A0_c_248_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_58 VPB N_A0_c_249_n 0.0167504f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_59 VPB N_A0_c_247_n 0.0243624f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_60 VPB N_A1_c_301_n 0.016779f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_61 VPB N_A1_c_302_n 0.019327f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_62 VPB N_A1_c_299_n 0.0322253f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_63 VPB N_A1_c_300_n 0.00330882f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_64 VPB N_VPWR_c_341_n 0.0176419f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_65 VPB N_VPWR_c_342_n 0.00916705f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_66 VPB N_VPWR_c_343_n 0.0150788f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_67 VPB N_VPWR_c_344_n 0.0139346f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_68 VPB N_VPWR_c_345_n 0.0674102f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_69 VPB N_VPWR_c_340_n 0.0472638f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.19
cc_70 VPB N_VPWR_c_347_n 0.00547281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_348_n 0.00547281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_349_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_211_297#_c_411_n 0.00583938f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_74 VPB N_A_399_297#_c_458_n 0.00609927f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_75 VPB N_A_399_297#_c_459_n 0.00219389f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_76 VPB Y 0.0367211f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_77 VPB Y 0.00219582f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_78 VPB N_Y_c_498_n 0.00762094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 N_S_c_87_n N_A_27_47#_c_153_n 0.0368923f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_80 N_S_c_82_n N_A_27_47#_M1008_g 0.0118845f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_81 N_S_c_85_n N_A_27_47#_c_149_n 0.00302677f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_82 N_S_c_80_n N_A_27_47#_c_149_n 0.00680542f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_83 S N_A_27_47#_c_149_n 0.0335266f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_84 N_S_c_84_n N_A_27_47#_c_149_n 0.0123555f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_85 N_S_c_85_n N_A_27_47#_c_168_n 0.0182811f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_86 N_S_c_86_n N_A_27_47#_c_168_n 0.0203972f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_87 N_S_c_87_n N_A_27_47#_c_168_n 0.00819184f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_88 S N_A_27_47#_c_168_n 0.0275105f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_89 N_S_c_84_n N_A_27_47#_c_168_n 0.00838399f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_90 N_S_c_86_n N_A_27_47#_c_156_n 0.00147276f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_91 N_S_c_87_n N_A_27_47#_c_156_n 0.00202709f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_92 N_S_c_84_n N_A_27_47#_c_156_n 0.00410836f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_93 S N_A_27_47#_c_176_n 0.00575572f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_94 N_S_c_84_n N_A_27_47#_c_176_n 0.0137142f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_95 N_S_c_85_n N_A_27_47#_c_159_n 0.0163567f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_96 N_S_c_84_n N_A_27_47#_c_179_n 5.74744e-19 $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_97 N_S_c_84_n N_A_27_47#_c_152_n 0.0209873f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_98 N_S_c_85_n N_VPWR_c_343_n 0.00429282f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_99 N_S_c_86_n N_VPWR_c_344_n 0.00554924f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_100 N_S_c_87_n N_VPWR_c_344_n 0.0032009f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_101 N_S_c_85_n N_VPWR_c_340_n 0.00824125f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_102 N_S_c_86_n N_VPWR_c_340_n 0.00826794f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_103 N_S_c_87_n N_VPWR_c_340_n 0.00390148f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_104 N_S_c_85_n N_VPWR_c_347_n 0.0119938f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_105 N_S_c_86_n N_VPWR_c_347_n 0.00846253f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_106 N_S_c_87_n N_VPWR_c_347_n 0.00106505f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_107 N_S_c_86_n N_VPWR_c_348_n 0.00118604f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_108 N_S_c_87_n N_VPWR_c_348_n 0.0112739f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_109 N_S_c_85_n N_A_211_297#_c_412_n 8.47478e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_110 N_S_c_86_n N_A_211_297#_c_412_n 0.00668236f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_111 N_S_c_87_n N_A_211_297#_c_412_n 0.0111799f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_112 N_S_c_87_n N_A_211_297#_c_415_n 0.00343832f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_113 N_S_c_87_n N_A_211_297#_c_416_n 6.53439e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_114 S N_VGND_M1011_d 0.00434139f $X=0.66 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_115 N_S_c_80_n N_VGND_c_549_n 0.0162081f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_116 N_S_c_81_n N_VGND_c_549_n 0.00310434f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_117 S N_VGND_c_549_n 0.0179379f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_118 N_S_c_84_n N_VGND_c_549_n 6.07153e-19 $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_119 N_S_c_81_n N_VGND_c_550_n 0.00585385f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_120 N_S_c_82_n N_VGND_c_550_n 0.00585385f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_121 N_S_c_82_n N_VGND_c_551_n 0.00304374f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_122 N_S_c_80_n N_VGND_c_554_n 0.00271402f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_123 N_S_c_80_n N_VGND_c_556_n 0.00600638f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_124 N_S_c_81_n N_VGND_c_556_n 0.0108216f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_125 N_S_c_82_n N_VGND_c_556_n 0.00653348f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_126 S N_VGND_c_556_n 8.77277e-19 $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_127 N_S_c_82_n N_A_213_47#_c_623_n 0.00392239f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_128 N_S_c_81_n N_A_213_47#_c_624_n 0.00412164f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_129 N_S_c_82_n N_A_213_47#_c_624_n 0.00184102f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_130 S N_A_213_47#_c_624_n 0.00732065f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_131 N_S_c_84_n N_A_213_47#_c_624_n 0.00393542f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_132 N_S_c_81_n N_A_213_47#_c_627_n 7.31634e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_133 N_S_c_82_n N_A_213_47#_c_627_n 0.00138038f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_134 S N_A_213_47#_c_627_n 0.00649219f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_135 N_S_c_84_n N_A_213_47#_c_627_n 0.00419187f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_179_n A0 0.00639636f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_152_n A0 9.64383e-19 $X=2.375 $Y=1.217 $X2=0 $Y2=0
cc_138 N_A_27_47#_M1012_g N_A0_c_246_n 0.0179705f $X=2.4 $Y=0.56 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_179_n N_A0_c_246_n 2.57595e-19 $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_168_n N_VPWR_M1005_d 0.0049392f $X=1.325 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A_27_47#_c_153_n N_VPWR_c_341_n 0.00574732f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_c_154_n N_VPWR_c_341_n 0.00523784f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_c_154_n N_VPWR_c_342_n 0.00604513f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_c_158_n N_VPWR_c_343_n 0.0179125f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_145 N_A_27_47#_M1005_s N_VPWR_c_340_n 0.00425811f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_c_153_n N_VPWR_c_340_n 0.00878938f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_c_154_n N_VPWR_c_340_n 0.0081693f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_158_n N_VPWR_c_340_n 0.00987844f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_168_n N_VPWR_c_347_n 0.00786103f $X=1.325 $Y=1.58 $X2=0
+ $Y2=0
cc_150 N_A_27_47#_c_158_n N_VPWR_c_347_n 0.0161786f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_153_n N_VPWR_c_348_n 0.00787181f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_154_n N_VPWR_c_348_n 0.00107191f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_168_n N_A_211_297#_M1001_d 0.00412421f $X=1.325 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_154 N_A_27_47#_c_153_n N_A_211_297#_c_412_n 0.00622416f $X=1.905 $Y=1.41
+ $X2=0 $Y2=0
cc_155 N_A_27_47#_c_168_n N_A_211_297#_c_412_n 0.0308469f $X=1.325 $Y=1.58 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_151_n N_A_211_297#_c_412_n 0.00509811f $X=1.805 $Y=1.2 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_153_n N_A_211_297#_c_415_n 0.00463061f $X=1.905 $Y=1.41
+ $X2=0 $Y2=0
cc_158 N_A_27_47#_c_154_n N_A_211_297#_c_415_n 8.67348e-19 $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_159 N_A_27_47#_c_153_n N_A_211_297#_c_416_n 0.00319588f $X=1.905 $Y=1.41
+ $X2=0 $Y2=0
cc_160 N_A_27_47#_c_151_n N_A_211_297#_c_416_n 0.0106271f $X=1.805 $Y=1.2 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_153_n N_A_211_297#_c_411_n 0.0100999f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_154_n N_A_211_297#_c_411_n 0.0161745f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_179_n N_A_211_297#_c_411_n 0.0188545f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_152_n N_A_211_297#_c_411_n 0.00648147f $X=2.375 $Y=1.217
+ $X2=0 $Y2=0
cc_165 N_A_27_47#_c_153_n N_A_399_297#_c_460_n 0.00423074f $X=1.905 $Y=1.41
+ $X2=0 $Y2=0
cc_166 N_A_27_47#_c_154_n N_A_399_297#_c_458_n 0.0152363f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_154_n N_A_399_297#_c_459_n 0.00233762f $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_168 N_A_27_47#_c_150_n N_VGND_c_549_n 0.015377f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_169 N_A_27_47#_M1008_g N_VGND_c_551_n 0.00322323f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_179_n N_VGND_c_551_n 0.00121936f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_151_n N_VGND_c_551_n 0.00871156f $X=1.805 $Y=1.2 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_152_n N_VGND_c_551_n 0.00107349f $X=2.375 $Y=1.217 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_M1008_g N_VGND_c_552_n 0.00585385f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A_27_47#_M1012_g N_VGND_c_552_n 0.00439206f $X=2.4 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1012_g N_VGND_c_553_n 0.00438629f $X=2.4 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_150_n N_VGND_c_554_n 0.0113284f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_177 N_A_27_47#_M1011_s N_VGND_c_556_n 0.00611128f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_M1008_g N_VGND_c_556_n 0.00647025f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_179 N_A_27_47#_M1012_g N_VGND_c_556_n 0.00702789f $X=2.4 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_150_n N_VGND_c_556_n 0.00939877f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_181 N_A_27_47#_M1008_g N_A_213_47#_c_623_n 0.00511627f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_M1012_g N_A_213_47#_c_623_n 0.00251402f $X=2.4 $Y=0.56 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_176_n N_A_213_47#_c_623_n 0.00588571f $X=1.545 $Y=1.24 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_179_n N_A_213_47#_c_623_n 0.013236f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_151_n N_A_213_47#_c_623_n 0.00714923f $X=1.805 $Y=1.2 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_152_n N_A_213_47#_c_623_n 0.00523968f $X=2.375 $Y=1.217
+ $X2=0 $Y2=0
cc_187 N_A_27_47#_M1008_g N_A_213_47#_c_624_n 2.01873e-19 $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_168_n N_A_213_47#_c_624_n 0.00479736f $X=1.325 $Y=1.58 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_176_n N_A_213_47#_c_624_n 0.00296915f $X=1.545 $Y=1.24 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_168_n N_A_213_47#_c_627_n 0.00350752f $X=1.325 $Y=1.58 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_176_n N_A_213_47#_c_627_n 0.00152247f $X=1.545 $Y=1.24 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1012_g N_A_401_47#_c_690_n 0.0049342f $X=2.4 $Y=0.56 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_M1008_g N_A_401_47#_c_687_n 0.00131581f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_179_n N_A_401_47#_c_687_n 0.00859309f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_152_n N_A_401_47#_c_687_n 0.0031979f $X=2.375 $Y=1.217 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_M1012_g N_A_401_47#_c_689_n 0.0149303f $X=2.4 $Y=0.56 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_152_n N_A_401_47#_c_689_n 2.60861e-19 $X=2.375 $Y=1.217
+ $X2=0 $Y2=0
cc_198 N_A0_c_244_n N_A1_c_297_n 0.0231532f $X=3.86 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_199 N_A0_c_249_n N_A1_c_301_n 0.0359664f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_200 A0 N_A1_c_299_n 0.00538576f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_201 N_A0_c_247_n N_A1_c_299_n 0.022136f $X=3.835 $Y=1.202 $X2=0 $Y2=0
cc_202 N_A0_c_248_n N_VPWR_c_342_n 0.00283134f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A0_c_248_n N_VPWR_c_345_n 0.00439333f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A0_c_249_n N_VPWR_c_345_n 0.00439333f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A0_c_248_n N_VPWR_c_340_n 0.00736527f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A0_c_249_n N_VPWR_c_340_n 0.00620037f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A0_c_248_n N_A_211_297#_c_429_n 0.00558766f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A0_c_249_n N_A_211_297#_c_429_n 0.00507402f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A0_c_247_n N_A_211_297#_c_429_n 0.00649224f $X=3.835 $Y=1.202 $X2=0
+ $Y2=0
cc_210 N_A0_c_248_n N_A_211_297#_c_411_n 0.0093264f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_211 A0 N_A_211_297#_c_411_n 0.0531344f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_212 N_A0_c_246_n N_A_211_297#_c_411_n 0.0117285f $X=3.265 $Y=1.145 $X2=0
+ $Y2=0
cc_213 N_A0_c_248_n N_A_399_297#_c_463_n 0.0140002f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A0_c_249_n N_A_399_297#_c_463_n 0.0144075f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_215 A0 N_A_399_297#_c_463_n 0.00558315f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_216 N_A0_c_248_n N_A_399_297#_c_459_n 0.00341345f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A0_c_243_n N_Y_c_494_n 0.00846157f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A0_c_244_n N_Y_c_494_n 0.00996531f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_219 A0 N_Y_c_494_n 0.00219523f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_220 N_A0_c_248_n Y 0.0092122f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A0_c_249_n Y 0.0092122f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A0_c_243_n N_VGND_c_553_n 0.00223443f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A0_c_243_n N_VGND_c_555_n 0.00366111f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A0_c_244_n N_VGND_c_555_n 0.00366111f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A0_c_243_n N_VGND_c_556_n 0.00664141f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A0_c_244_n N_VGND_c_556_n 0.00543797f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A0_c_243_n N_A_213_47#_c_623_n 0.00168096f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A0_c_244_n N_A_213_47#_c_623_n 0.00449987f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_229 A0 N_A_213_47#_c_623_n 0.0333114f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_230 N_A0_c_246_n N_A_213_47#_c_623_n 0.0151175f $X=3.265 $Y=1.145 $X2=0 $Y2=0
cc_231 N_A0_c_247_n N_A_213_47#_c_623_n 0.00446818f $X=3.835 $Y=1.202 $X2=0
+ $Y2=0
cc_232 N_A0_c_244_n N_A_213_47#_c_625_n 0.0014135f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A0_c_244_n N_A_213_47#_c_626_n 0.00145722f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A0_c_243_n N_A_401_47#_c_688_n 0.00705448f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A0_c_244_n N_A_401_47#_c_688_n 5.84999e-19 $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A0_c_247_n N_A_401_47#_c_688_n 0.00340407f $X=3.835 $Y=1.202 $X2=0
+ $Y2=0
cc_237 N_A0_c_243_n N_A_401_47#_c_689_n 0.00685935f $X=3.39 $Y=0.995 $X2=0 $Y2=0
cc_238 A0 N_A_401_47#_c_689_n 0.0657531f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_239 N_A0_c_246_n N_A_401_47#_c_689_n 0.0143083f $X=3.265 $Y=1.145 $X2=0 $Y2=0
cc_240 N_A1_c_301_n N_VPWR_c_345_n 0.00439333f $X=4.345 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A1_c_302_n N_VPWR_c_345_n 0.00439333f $X=4.82 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A1_c_301_n N_VPWR_c_340_n 0.00621361f $X=4.345 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A1_c_302_n N_VPWR_c_340_n 0.00715012f $X=4.82 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A1_c_301_n N_A_211_297#_c_429_n 9.91692e-19 $X=4.345 $Y=1.41 $X2=0
+ $Y2=0
cc_245 N_A1_c_301_n N_A_399_297#_c_463_n 0.0154152f $X=4.345 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A1_c_302_n N_A_399_297#_c_463_n 0.00365011f $X=4.82 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A1_c_299_n N_A_399_297#_c_463_n 0.00581419f $X=4.82 $Y=1.202 $X2=0
+ $Y2=0
cc_248 N_A1_c_300_n N_A_399_297#_c_463_n 9.36343e-19 $X=4.95 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A1_c_300_n N_Y_M1013_d 0.00394172f $X=4.95 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A1_c_297_n N_Y_c_494_n 0.008274f $X=4.32 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A1_c_298_n N_Y_c_494_n 0.0136127f $X=4.795 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A1_c_299_n N_Y_c_494_n 0.00291747f $X=4.82 $Y=1.202 $X2=0 $Y2=0
cc_253 N_A1_c_300_n N_Y_c_494_n 0.00966005f $X=4.95 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A1_c_298_n Y 0.012736f $X=4.795 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A1_c_302_n Y 0.0170776f $X=4.82 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A1_c_299_n Y 0.00990156f $X=4.82 $Y=1.202 $X2=0 $Y2=0
cc_257 N_A1_c_300_n Y 0.0478942f $X=4.95 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A1_c_301_n Y 0.00924199f $X=4.345 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A1_c_302_n Y 0.0115484f $X=4.82 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A1_c_300_n Y 0.00747058f $X=4.95 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A1_c_297_n N_VGND_c_555_n 0.00366111f $X=4.32 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A1_c_298_n N_VGND_c_555_n 0.00366111f $X=4.795 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A1_c_297_n N_VGND_c_556_n 0.00540196f $X=4.32 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A1_c_298_n N_VGND_c_556_n 0.00659174f $X=4.795 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A1_c_297_n N_A_213_47#_c_625_n 0.00650596f $X=4.32 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A1_c_298_n N_A_213_47#_c_625_n 4.62395e-19 $X=4.795 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A1_c_297_n N_A_213_47#_c_626_n 0.0114758f $X=4.32 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A1_c_298_n N_A_213_47#_c_626_n 0.00617504f $X=4.795 $Y=0.995 $X2=0
+ $Y2=0
cc_269 N_A1_c_299_n N_A_213_47#_c_626_n 0.00560309f $X=4.82 $Y=1.202 $X2=0 $Y2=0
cc_270 N_A1_c_300_n N_A_213_47#_c_626_n 0.00224159f $X=4.95 $Y=1.16 $X2=0 $Y2=0
cc_271 N_VPWR_c_340_n N_A_211_297#_M1001_d 0.0037272f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_272 N_VPWR_c_340_n N_A_211_297#_M1004_d 0.00235479f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_273 N_VPWR_M1014_s N_A_211_297#_c_412_n 0.00456705f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_341_n N_A_211_297#_c_412_n 7.38269e-19 $X=2.525 $Y=2.72 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_344_n N_A_211_297#_c_412_n 0.00595845f $X=1.455 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_340_n N_A_211_297#_c_412_n 0.0145702f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_348_n N_A_211_297#_c_412_n 0.0143686f $X=1.67 $Y=2.34 $X2=0
+ $Y2=0
cc_278 N_VPWR_M1014_s N_A_211_297#_c_415_n 0.00197555f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_279 N_VPWR_M1014_s N_A_211_297#_c_416_n 0.00193612f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_280 N_VPWR_M1009_d N_A_211_297#_c_411_n 0.00693642f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_340_n N_A_399_297#_M1006_s 0.00432871f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_282 N_VPWR_c_340_n N_A_399_297#_M1010_s 0.00239539f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_341_n N_A_399_297#_c_460_n 0.0137694f $X=2.525 $Y=2.72 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_340_n N_A_399_297#_c_460_n 0.00861434f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_348_n N_A_399_297#_c_460_n 0.0131787f $X=1.67 $Y=2.34 $X2=0
+ $Y2=0
cc_286 N_VPWR_M1009_d N_A_399_297#_c_458_n 0.00525552f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_341_n N_A_399_297#_c_458_n 0.00299202f $X=2.525 $Y=2.72 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_342_n N_A_399_297#_c_458_n 0.0194775f $X=2.61 $Y=2.34 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_345_n N_A_399_297#_c_458_n 0.0029367f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_340_n N_A_399_297#_c_458_n 0.0116347f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_340_n N_Y_M1004_s 0.0021994f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_340_n N_Y_M1015_s 0.00266335f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_293 N_VPWR_c_340_n N_Y_M1013_d 0.00381498f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_c_342_n Y 0.0134692f $X=2.61 $Y=2.34 $X2=0 $Y2=0
cc_295 N_VPWR_c_345_n Y 0.101709f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_296 N_VPWR_c_340_n Y 0.0775947f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_297 N_VPWR_c_345_n N_Y_c_498_n 0.0126008f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_298 N_VPWR_c_340_n N_Y_c_498_n 0.00848438f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_299 N_A_211_297#_c_411_n N_A_399_297#_M1006_s 0.00382328f $X=3.385 $Y=1.605
+ $X2=-0.19 $Y2=1.305
cc_300 N_A_211_297#_M1004_d N_A_399_297#_c_463_n 0.00363051f $X=3.455 $Y=1.485
+ $X2=0 $Y2=0
cc_301 N_A_211_297#_c_429_n N_A_399_297#_c_463_n 0.0169588f $X=3.6 $Y=1.63 $X2=0
+ $Y2=0
cc_302 N_A_211_297#_c_411_n N_A_399_297#_c_463_n 0.00996357f $X=3.385 $Y=1.605
+ $X2=0 $Y2=0
cc_303 N_A_211_297#_c_412_n N_A_399_297#_c_460_n 0.0119525f $X=1.715 $Y=1.92
+ $X2=0 $Y2=0
cc_304 N_A_211_297#_c_411_n N_A_399_297#_c_460_n 0.0115274f $X=3.385 $Y=1.605
+ $X2=0 $Y2=0
cc_305 N_A_211_297#_c_411_n N_A_399_297#_c_458_n 0.0577788f $X=3.385 $Y=1.605
+ $X2=0 $Y2=0
cc_306 N_A_211_297#_c_411_n N_Y_M1004_s 0.0052299f $X=3.385 $Y=1.605 $X2=0 $Y2=0
cc_307 N_A_211_297#_M1004_d Y 0.00367601f $X=3.455 $Y=1.485 $X2=0 $Y2=0
cc_308 N_A_211_297#_c_411_n N_A_213_47#_c_623_n 0.0121415f $X=3.385 $Y=1.605
+ $X2=0 $Y2=0
cc_309 N_A_211_297#_c_411_n N_A_401_47#_c_687_n 6.95363e-19 $X=3.385 $Y=1.605
+ $X2=0 $Y2=0
cc_310 N_A_211_297#_c_411_n N_A_401_47#_c_689_n 0.00676562f $X=3.385 $Y=1.605
+ $X2=0 $Y2=0
cc_311 N_A_399_297#_c_463_n N_Y_M1004_s 0.00178471f $X=4.585 $Y=2 $X2=0 $Y2=0
cc_312 N_A_399_297#_c_459_n N_Y_M1004_s 0.00490776f $X=3.135 $Y=1.96 $X2=0 $Y2=0
cc_313 N_A_399_297#_c_463_n N_Y_M1015_s 0.0097009f $X=4.585 $Y=2 $X2=0 $Y2=0
cc_314 N_A_399_297#_c_463_n Y 0.00631114f $X=4.585 $Y=2 $X2=0 $Y2=0
cc_315 N_A_399_297#_M1010_s Y 0.00378044f $X=4.435 $Y=1.485 $X2=0 $Y2=0
cc_316 N_A_399_297#_c_459_n Y 0.0931964f $X=3.135 $Y=1.96 $X2=0 $Y2=0
cc_317 N_Y_c_494_n N_VGND_c_553_n 0.0100248f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_318 N_Y_c_494_n N_VGND_c_555_n 0.114284f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_319 N_Y_M1000_d N_VGND_c_556_n 0.0020813f $X=3.005 $Y=0.235 $X2=0 $Y2=0
cc_320 N_Y_M1003_d N_VGND_c_556_n 0.00202839f $X=3.935 $Y=0.235 $X2=0 $Y2=0
cc_321 N_Y_M1017_s N_VGND_c_556_n 0.00415481f $X=4.87 $Y=0.235 $X2=0 $Y2=0
cc_322 N_Y_c_494_n N_VGND_c_556_n 0.0576677f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_323 N_Y_c_494_n N_A_213_47#_M1007_d 0.00431812f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_324 N_Y_M1003_d N_A_213_47#_c_623_n 0.0016435f $X=3.935 $Y=0.235 $X2=0 $Y2=0
cc_325 N_Y_c_494_n N_A_213_47#_c_623_n 0.00905399f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_326 N_Y_M1003_d N_A_213_47#_c_625_n 9.37216e-19 $X=3.935 $Y=0.235 $X2=0 $Y2=0
cc_327 N_Y_c_494_n N_A_213_47#_c_625_n 0.00261211f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_328 N_Y_c_494_n N_A_213_47#_c_626_n 0.0229179f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_329 Y N_A_213_47#_c_626_n 0.00555158f $X=5.2 $Y=1.785 $X2=0 $Y2=0
cc_330 N_Y_c_494_n N_A_401_47#_M1000_s 0.00412092f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_331 N_Y_c_494_n N_A_401_47#_c_688_n 0.0165395f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_332 N_Y_M1000_d N_A_401_47#_c_689_n 0.00429312f $X=3.005 $Y=0.235 $X2=0 $Y2=0
cc_333 N_Y_c_494_n N_A_401_47#_c_689_n 0.0141755f $X=5.255 $Y=0.38 $X2=0 $Y2=0
cc_334 N_VGND_c_556_n N_A_213_47#_M1002_d 0.00433793f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_335 N_VGND_c_556_n N_A_213_47#_M1007_d 0.00249538f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_336 N_VGND_M1016_s N_A_213_47#_c_623_n 9.36802e-19 $X=1.535 $Y=0.235 $X2=0
+ $Y2=0
cc_337 N_VGND_c_551_n N_A_213_47#_c_623_n 0.0136805f $X=1.67 $Y=0.38 $X2=0 $Y2=0
cc_338 N_VGND_c_553_n N_A_213_47#_c_623_n 8.4091e-19 $X=2.61 $Y=0.38 $X2=0 $Y2=0
cc_339 N_VGND_c_556_n N_A_213_47#_c_623_n 0.126297f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_340 N_VGND_c_551_n N_A_213_47#_c_624_n 0.00114639f $X=1.67 $Y=0.38 $X2=0
+ $Y2=0
cc_341 N_VGND_c_556_n N_A_213_47#_c_624_n 0.0148735f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_342 N_VGND_c_556_n N_A_213_47#_c_625_n 0.0171571f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_343 N_VGND_c_550_n N_A_213_47#_c_627_n 0.00472818f $X=1.585 $Y=0 $X2=0 $Y2=0
cc_344 N_VGND_c_551_n N_A_213_47#_c_627_n 0.00338192f $X=1.67 $Y=0.38 $X2=0
+ $Y2=0
cc_345 N_VGND_c_556_n N_A_213_47#_c_627_n 0.00317372f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_556_n N_A_401_47#_M1008_s 0.00280589f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_347 N_VGND_c_556_n N_A_401_47#_M1000_s 0.00213276f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_348 N_VGND_c_552_n N_A_401_47#_c_690_n 0.00915794f $X=2.525 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_c_556_n N_A_401_47#_c_690_n 0.00300001f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_350 N_VGND_c_551_n N_A_401_47#_c_687_n 0.00296978f $X=1.67 $Y=0.38 $X2=0
+ $Y2=0
cc_351 N_VGND_M1012_d N_A_401_47#_c_689_n 0.00319634f $X=2.475 $Y=0.235 $X2=0
+ $Y2=0
cc_352 N_VGND_c_552_n N_A_401_47#_c_689_n 0.00337093f $X=2.525 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_553_n N_A_401_47#_c_689_n 0.0102463f $X=2.61 $Y=0.38 $X2=0 $Y2=0
cc_354 N_VGND_c_555_n N_A_401_47#_c_689_n 0.00399916f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_355 N_VGND_c_556_n N_A_401_47#_c_689_n 0.00749316f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_356 N_A_213_47#_c_623_n N_A_401_47#_M1008_s 6.95505e-19 $X=4.14 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_357 N_A_213_47#_c_623_n N_A_401_47#_c_687_n 0.0096269f $X=4.14 $Y=0.85 $X2=0
+ $Y2=0
cc_358 N_A_213_47#_c_623_n N_A_401_47#_c_688_n 0.0148111f $X=4.14 $Y=0.85 $X2=0
+ $Y2=0
cc_359 N_A_213_47#_c_625_n N_A_401_47#_c_688_n 0.00125486f $X=4.285 $Y=0.85
+ $X2=0 $Y2=0
cc_360 N_A_213_47#_c_626_n N_A_401_47#_c_688_n 0.00228781f $X=4.285 $Y=0.85
+ $X2=0 $Y2=0
cc_361 N_A_213_47#_c_623_n N_A_401_47#_c_689_n 0.0410939f $X=4.14 $Y=0.85 $X2=0
+ $Y2=0
