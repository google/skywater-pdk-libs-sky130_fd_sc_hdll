* File: sky130_fd_sc_hdll__nand2_4.pxi.spice
* Created: Thu Aug 27 19:12:55 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2_4%B N_B_c_65_n N_B_M1001_g N_B_c_59_n N_B_M1002_g
+ N_B_c_66_n N_B_M1006_g N_B_c_60_n N_B_M1010_g N_B_c_67_n N_B_M1009_g
+ N_B_c_61_n N_B_M1011_g N_B_c_68_n N_B_M1014_g N_B_c_62_n N_B_M1015_g B B B B
+ N_B_c_63_n B B B B PM_SKY130_FD_SC_HDLL__NAND2_4%B
x_PM_SKY130_FD_SC_HDLL__NAND2_4%A N_A_c_143_n N_A_M1005_g N_A_c_149_n
+ N_A_M1000_g N_A_c_144_n N_A_M1008_g N_A_c_150_n N_A_M1003_g N_A_c_145_n
+ N_A_M1012_g N_A_c_151_n N_A_M1004_g N_A_c_152_n N_A_M1007_g N_A_c_146_n
+ N_A_M1013_g A A N_A_c_147_n N_A_c_148_n A A PM_SKY130_FD_SC_HDLL__NAND2_4%A
x_PM_SKY130_FD_SC_HDLL__NAND2_4%VPWR N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_M1014_d N_VPWR_M1003_d N_VPWR_M1007_d N_VPWR_c_218_n N_VPWR_c_219_n
+ N_VPWR_c_220_n N_VPWR_c_221_n N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n
+ N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n
+ VPWR N_VPWR_c_230_n N_VPWR_c_217_n N_VPWR_c_232_n N_VPWR_c_233_n
+ PM_SKY130_FD_SC_HDLL__NAND2_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2_4%Y N_Y_M1005_s N_Y_M1012_s N_Y_M1001_s
+ N_Y_M1009_s N_Y_M1000_s N_Y_M1004_s N_Y_c_291_n N_Y_c_295_n N_Y_c_298_n
+ N_Y_c_302_n N_Y_c_305_n N_Y_c_307_n N_Y_c_320_n N_Y_c_324_n N_Y_c_328_n
+ N_Y_c_332_n N_Y_c_308_n N_Y_c_335_n Y Y PM_SKY130_FD_SC_HDLL__NAND2_4%Y
x_PM_SKY130_FD_SC_HDLL__NAND2_4%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1010_d
+ N_A_27_47#_M1015_d N_A_27_47#_M1008_d N_A_27_47#_M1013_d N_A_27_47#_c_382_n
+ N_A_27_47#_c_383_n N_A_27_47#_c_384_n N_A_27_47#_c_396_n N_A_27_47#_c_385_n
+ N_A_27_47#_c_402_n N_A_27_47#_c_386_n N_A_27_47#_c_408_n N_A_27_47#_c_387_n
+ N_A_27_47#_c_388_n N_A_27_47#_c_389_n PM_SKY130_FD_SC_HDLL__NAND2_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND2_4%VGND N_VGND_M1002_s N_VGND_M1011_s
+ N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n VGND N_VGND_c_455_n
+ N_VGND_c_456_n N_VGND_c_457_n N_VGND_c_458_n
+ PM_SKY130_FD_SC_HDLL__NAND2_4%VGND
cc_1 VNB N_B_c_59_n 0.0219752f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_B_c_60_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_B_c_61_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_4 VNB N_B_c_62_n 0.0164854f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_B_c_63_n 0.0970829f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_6 VNB B 0.00932659f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.19
cc_7 VNB N_A_c_143_n 0.0162503f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_A_c_144_n 0.0169272f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_9 VNB N_A_c_145_n 0.0174114f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_10 VNB N_A_c_146_n 0.0229091f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_11 VNB N_A_c_147_n 0.0122746f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_12 VNB N_A_c_148_n 0.0821252f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_13 VNB N_VPWR_c_217_n 0.193827f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.19
cc_14 VNB Y 0.00106016f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.2
cc_15 VNB N_A_27_47#_c_382_n 0.0182049f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_16 VNB N_A_27_47#_c_383_n 0.00258613f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_17 VNB N_A_27_47#_c_384_n 0.0102713f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_18 VNB N_A_27_47#_c_385_n 0.00264996f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_19 VNB N_A_27_47#_c_386_n 0.00370326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_387_n 0.00914706f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_21 VNB N_A_27_47#_c_388_n 0.0201677f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_22 VNB N_A_27_47#_c_389_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_23 VNB N_VGND_c_452_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_24 VNB N_VGND_c_453_n 0.0192454f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_25 VNB N_VGND_c_454_n 0.00467885f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_26 VNB N_VGND_c_455_n 0.070111f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_27 VNB N_VGND_c_456_n 0.251358f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_28 VNB N_VGND_c_457_n 0.0219327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_458_n 0.003239f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.202
cc_30 VPB N_B_c_65_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_31 VPB N_B_c_66_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_32 VPB N_B_c_67_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_33 VPB N_B_c_68_n 0.0164383f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_34 VPB N_B_c_63_n 0.0574824f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_35 VPB B 7.73822e-19 $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.19
cc_36 VPB N_A_c_149_n 0.0161146f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_37 VPB N_A_c_150_n 0.0162386f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_38 VPB N_A_c_151_n 0.016261f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_39 VPB N_A_c_152_n 0.0210879f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_40 VPB N_A_c_147_n 0.00528555f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_41 VPB N_A_c_148_n 0.0489731f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_42 VPB N_VPWR_c_218_n 0.00994749f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_43 VPB N_VPWR_c_219_n 0.0428682f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_44 VPB N_VPWR_c_220_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_45 VPB N_VPWR_c_221_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_46 VPB N_VPWR_c_222_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.105
cc_47 VPB N_VPWR_c_223_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_224_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_49 VPB N_VPWR_c_225_n 0.0310182f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.202
cc_50 VPB N_VPWR_c_226_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.67 $Y2=1.16
cc_51 VPB N_VPWR_c_227_n 0.00324069f $X=-0.19 $Y=1.305 $X2=1.67 $Y2=1.16
cc_52 VPB N_VPWR_c_228_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.202
cc_53 VPB N_VPWR_c_229_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_54 VPB N_VPWR_c_230_n 0.0153494f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.2
cc_55 VPB N_VPWR_c_217_n 0.0562661f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.19
cc_56 VPB N_VPWR_c_232_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_233_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB Y 0.00155805f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.2
cc_59 N_B_c_62_n N_A_c_143_n 0.0171111f $X=1.93 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_60 N_B_c_68_n N_A_c_149_n 0.0230725f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_61 N_B_c_63_n N_A_c_148_n 0.0171111f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_62 B N_A_c_148_n 9.46922e-19 $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_63 N_B_c_65_n N_VPWR_c_219_n 0.00777002f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_64 N_B_c_63_n N_VPWR_c_219_n 0.00545118f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_65 B N_VPWR_c_219_n 0.0190002f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_66 N_B_c_65_n N_VPWR_c_220_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_67 N_B_c_66_n N_VPWR_c_220_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_68 N_B_c_66_n N_VPWR_c_221_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_69 N_B_c_67_n N_VPWR_c_221_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_70 N_B_c_67_n N_VPWR_c_222_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_71 N_B_c_68_n N_VPWR_c_222_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_72 N_B_c_68_n N_VPWR_c_223_n 0.0052072f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_73 N_B_c_65_n N_VPWR_c_217_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_B_c_66_n N_VPWR_c_217_n 0.0118438f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_75 N_B_c_67_n N_VPWR_c_217_n 0.00999457f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_76 N_B_c_68_n N_VPWR_c_217_n 0.011869f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_77 N_B_c_65_n N_Y_c_291_n 0.00347232f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_78 N_B_c_66_n N_Y_c_291_n 5.79575e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_79 N_B_c_63_n N_Y_c_291_n 0.00651614f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_80 B N_Y_c_291_n 0.0253353f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_81 N_B_c_65_n N_Y_c_295_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B_c_66_n N_Y_c_295_n 0.0106251f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B_c_67_n N_Y_c_295_n 6.24674e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B_c_66_n N_Y_c_298_n 0.0137916f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B_c_67_n N_Y_c_298_n 0.0101048f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B_c_63_n N_Y_c_298_n 0.00635951f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_87 B N_Y_c_298_n 0.0356113f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_88 N_B_c_66_n N_Y_c_302_n 6.48386e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B_c_67_n N_Y_c_302_n 0.0130707f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B_c_68_n N_Y_c_302_n 0.0106251f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B_c_68_n N_Y_c_305_n 0.015284f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_92 B N_Y_c_305_n 0.00310934f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_93 N_B_c_68_n N_Y_c_307_n 6.48386e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_c_67_n N_Y_c_308_n 0.00210477f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B_c_68_n N_Y_c_308_n 5.79575e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B_c_63_n N_Y_c_308_n 0.00651614f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_97 B N_Y_c_308_n 0.0253353f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_98 N_B_c_68_n Y 4.25242e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B_c_62_n Y 0.0023522f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_100 B Y 0.00792228f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_101 N_B_c_59_n N_A_27_47#_c_383_n 0.0113247f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B_c_60_n N_A_27_47#_c_383_n 0.00640878f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_103 N_B_c_63_n N_A_27_47#_c_383_n 0.0040376f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_104 B N_A_27_47#_c_383_n 0.0406647f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_105 N_B_c_63_n N_A_27_47#_c_384_n 0.00815985f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_106 B N_A_27_47#_c_384_n 0.0259684f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_107 N_B_c_59_n N_A_27_47#_c_396_n 5.79378e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B_c_60_n N_A_27_47#_c_396_n 0.00837042f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B_c_61_n N_A_27_47#_c_385_n 0.0111264f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B_c_62_n N_A_27_47#_c_385_n 0.00700013f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B_c_63_n N_A_27_47#_c_385_n 0.00346f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_112 B N_A_27_47#_c_385_n 0.0375301f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_113 N_B_c_62_n N_A_27_47#_c_402_n 0.00359564f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B_c_61_n N_A_27_47#_c_386_n 5.18407e-19 $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B_c_62_n N_A_27_47#_c_386_n 0.00861768f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B_c_60_n N_A_27_47#_c_389_n 0.00281161f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B_c_63_n N_A_27_47#_c_389_n 0.00358305f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_118 B N_A_27_47#_c_389_n 0.030974f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_119 N_B_c_59_n N_VGND_c_452_n 0.00276126f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B_c_60_n N_VGND_c_452_n 0.0035663f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B_c_60_n N_VGND_c_453_n 0.00395968f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B_c_61_n N_VGND_c_453_n 0.00436487f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_61_n N_VGND_c_454_n 0.00276126f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B_c_62_n N_VGND_c_454_n 0.00356343f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B_c_62_n N_VGND_c_455_n 0.0039445f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B_c_59_n N_VGND_c_456_n 0.00698799f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_c_60_n N_VGND_c_456_n 0.0058034f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B_c_61_n N_VGND_c_456_n 0.0061161f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B_c_62_n N_VGND_c_456_n 0.00571271f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B_c_59_n N_VGND_c_457_n 0.00436487f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_149_n N_VPWR_c_223_n 0.004751f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_c_150_n N_VPWR_c_224_n 0.0052072f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_151_n N_VPWR_c_224_n 0.004751f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_152_n N_VPWR_c_225_n 0.00722921f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_147_n N_VPWR_c_225_n 0.00689375f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_149_n N_VPWR_c_226_n 0.00597712f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_c_150_n N_VPWR_c_226_n 0.00673617f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_151_n N_VPWR_c_228_n 0.00597712f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_152_n N_VPWR_c_228_n 0.00673617f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_149_n N_VPWR_c_217_n 0.0100198f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_150_n N_VPWR_c_217_n 0.0118438f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_151_n N_VPWR_c_217_n 0.00999457f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_152_n N_VPWR_c_217_n 0.0131262f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_149_n N_Y_c_302_n 6.24674e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_149_n N_Y_c_305_n 0.0133907f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_149_n N_Y_c_307_n 0.0130707f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_150_n N_Y_c_307_n 0.0106251f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_151_n N_Y_c_307_n 6.24674e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_144_n N_Y_c_320_n 0.0123878f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_c_145_n N_Y_c_320_n 0.00922871f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_c_147_n N_Y_c_320_n 0.0372461f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_c_148_n N_Y_c_320_n 0.00759225f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_153 N_A_c_150_n N_Y_c_324_n 0.0165098f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_151_n N_Y_c_324_n 0.0101048f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_147_n N_Y_c_324_n 0.0293587f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_c_148_n N_Y_c_324_n 0.00635951f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_157 N_A_c_151_n N_Y_c_328_n 0.00210477f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_152_n N_Y_c_328_n 0.00827826f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_147_n N_Y_c_328_n 0.0253353f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_c_148_n N_Y_c_328_n 0.00631893f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_161 N_A_c_150_n N_Y_c_332_n 6.48386e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_c_151_n N_Y_c_332_n 0.0130707f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_c_152_n N_Y_c_332_n 0.0153658f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_c_143_n N_Y_c_335_n 0.00219421f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_143_n Y 0.003837f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_c_149_n Y 0.00253311f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_144_n Y 0.00297612f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_c_150_n Y 0.00220286f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_147_n Y 0.019661f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_c_148_n Y 0.0351365f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_171 N_A_c_149_n Y 0.00110455f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_c_150_n Y 0.00129054f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_c_148_n Y 0.00128221f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_174 N_A_c_143_n N_A_27_47#_c_408_n 0.0127822f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_c_144_n N_A_27_47#_c_408_n 0.00903374f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_c_145_n N_A_27_47#_c_408_n 0.00935436f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_146_n N_A_27_47#_c_408_n 0.0114382f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_147_n N_A_27_47#_c_408_n 0.00475263f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_c_148_n N_A_27_47#_c_408_n 4.68623e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_180 N_A_c_147_n N_A_27_47#_c_388_n 0.013698f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_c_143_n N_VGND_c_455_n 0.00357877f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_c_144_n N_VGND_c_455_n 0.00357877f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_c_145_n N_VGND_c_455_n 0.00357877f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_c_146_n N_VGND_c_455_n 0.00357877f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_c_143_n N_VGND_c_456_n 0.00538422f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_c_144_n N_VGND_c_456_n 0.00548399f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_145_n N_VGND_c_456_n 0.00560377f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_146_n N_VGND_c_456_n 0.00662792f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_189 N_VPWR_c_217_n N_Y_M1001_s 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_190 N_VPWR_c_217_n N_Y_M1009_s 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_191 N_VPWR_c_217_n N_Y_M1000_s 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_217_n N_Y_M1004_s 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_219_n N_Y_c_291_n 0.0137498f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_194 N_VPWR_c_219_n N_Y_c_295_n 0.0615045f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_195 N_VPWR_c_220_n N_Y_c_295_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_196 N_VPWR_c_221_n N_Y_c_295_n 0.0385613f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_197 N_VPWR_c_217_n N_Y_c_295_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_M1006_d N_Y_c_298_n 0.00325884f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_199 N_VPWR_c_221_n N_Y_c_298_n 0.0136682f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_200 N_VPWR_c_221_n N_Y_c_302_n 0.0470327f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_201 N_VPWR_c_222_n N_Y_c_302_n 0.0223557f $X=2.055 $Y=2.72 $X2=0 $Y2=0
cc_202 N_VPWR_c_223_n N_Y_c_302_n 0.0385613f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_203 N_VPWR_c_217_n N_Y_c_302_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_204 N_VPWR_M1014_d N_Y_c_305_n 0.0051962f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_205 N_VPWR_c_223_n N_Y_c_305_n 0.0136682f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_206 N_VPWR_c_223_n N_Y_c_307_n 0.0470327f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_207 N_VPWR_c_224_n N_Y_c_307_n 0.0385613f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_208 N_VPWR_c_226_n N_Y_c_307_n 0.0223557f $X=2.995 $Y=2.72 $X2=0 $Y2=0
cc_209 N_VPWR_c_217_n N_Y_c_307_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_210 N_VPWR_M1003_d N_Y_c_324_n 0.00325884f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_211 N_VPWR_c_224_n N_Y_c_324_n 0.0136682f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_212 N_VPWR_c_224_n N_Y_c_332_n 0.0470327f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_213 N_VPWR_c_225_n N_Y_c_332_n 0.0396855f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_214 N_VPWR_c_228_n N_Y_c_332_n 0.0223557f $X=3.935 $Y=2.72 $X2=0 $Y2=0
cc_215 N_VPWR_c_217_n N_Y_c_332_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_216 N_VPWR_c_219_n N_A_27_47#_c_384_n 7.42972e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_217 N_Y_c_320_n N_A_27_47#_M1008_d 0.00439968f $X=3.55 $Y=0.72 $X2=0 $Y2=0
cc_218 N_Y_c_305_n N_A_27_47#_c_385_n 0.00108863f $X=2.395 $Y=1.58 $X2=0 $Y2=0
cc_219 N_Y_c_305_n N_A_27_47#_c_386_n 0.00881009f $X=2.395 $Y=1.58 $X2=0 $Y2=0
cc_220 Y N_A_27_47#_c_386_n 0.00456405f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_221 N_Y_M1005_s N_A_27_47#_c_408_n 0.00399738f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_222 N_Y_M1012_s N_A_27_47#_c_408_n 0.00507102f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_223 N_Y_c_320_n N_A_27_47#_c_408_n 0.0518873f $X=3.55 $Y=0.72 $X2=0 $Y2=0
cc_224 N_Y_c_335_n N_A_27_47#_c_408_n 0.0182216f $X=2.545 $Y=0.805 $X2=0 $Y2=0
cc_225 N_Y_M1005_s N_VGND_c_456_n 0.00256987f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_226 N_Y_M1012_s N_VGND_c_456_n 0.00297142f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_383_n N_VGND_M1002_s 0.0025045f $X=0.985 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_228 N_A_27_47#_c_385_n N_VGND_M1011_s 0.0025045f $X=1.925 $Y=0.81 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_383_n N_VGND_c_452_n 0.0127393f $X=0.985 $Y=0.81 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_396_n N_VGND_c_452_n 0.0216501f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_383_n N_VGND_c_453_n 0.0020445f $X=0.985 $Y=0.81 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_396_n N_VGND_c_453_n 0.023074f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_385_n N_VGND_c_453_n 0.00260993f $X=1.925 $Y=0.81 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_385_n N_VGND_c_454_n 0.0127393f $X=1.925 $Y=0.81 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_402_n N_VGND_c_454_n 0.0165057f $X=2.075 $Y=0.465 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_386_n N_VGND_c_454_n 0.00582645f $X=2.075 $Y=0.715 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_385_n N_VGND_c_455_n 0.0020445f $X=1.925 $Y=0.81 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_402_n N_VGND_c_455_n 0.0186086f $X=2.075 $Y=0.465 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_408_n N_VGND_c_455_n 0.0958611f $X=3.935 $Y=0.36 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_387_n N_VGND_c_455_n 0.0172955f $X=4.06 $Y=0.465 $X2=0 $Y2=0
cc_241 N_A_27_47#_M1002_d N_VGND_c_456_n 0.00258669f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_M1010_d N_VGND_c_456_n 0.0026371f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_M1015_d N_VGND_c_456_n 0.00215206f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_M1008_d N_VGND_c_456_n 0.00255381f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_M1013_d N_VGND_c_456_n 0.00209324f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_382_n N_VGND_c_456_n 0.0128092f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_383_n N_VGND_c_456_n 0.00988931f $X=0.985 $Y=0.81 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_396_n N_VGND_c_456_n 0.0141066f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_385_n N_VGND_c_456_n 0.00988931f $X=1.925 $Y=0.81 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_402_n N_VGND_c_456_n 0.0111017f $X=2.075 $Y=0.465 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_408_n N_VGND_c_456_n 0.0609578f $X=3.935 $Y=0.36 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_387_n N_VGND_c_456_n 0.00960883f $X=4.06 $Y=0.465 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_382_n N_VGND_c_457_n 0.0221535f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_383_n N_VGND_c_457_n 0.00260993f $X=0.985 $Y=0.81 $X2=0
+ $Y2=0
