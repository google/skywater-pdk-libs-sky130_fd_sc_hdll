* File: sky130_fd_sc_hdll__a211o_1.spice
* Created: Wed Sep  2 08:15:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a211o_1.pex.spice"
.subckt sky130_fd_sc_hdll__a211o_1  VNB VPB A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2925 AS=0.17225 PD=1.55 PS=1.83 NRD=23.988 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1007 A_320_47# N_A2_M1007_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65 AD=0.16575
+ AS=0.2925 PD=1.16 PS=1.55 NRD=36.912 NRS=23.988 M=1 R=4.33333 SA=75001.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1006 N_A_80_21#_M1006_d N_A1_M1006_g A_320_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.16575 PD=0.93 PS=1.16 NRD=0.912 NRS=36.912 M=1 R=4.33333
+ SA=75001.9 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_B1_M1001_g N_A_80_21#_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.091 PD=1.03 PS=0.93 NRD=15.684 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1009 N_A_80_21#_M1009_d N_C1_M1009_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.20475 AS=0.1235 PD=1.93 PS=1.03 NRD=9.228 NRS=2.76 M=1 R=4.33333
+ SA=75002.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_80_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.275 PD=2.55 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_227_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.24 AS=0.275 PD=1.48 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1008 N_A_227_297#_M1008_d N_A1_M1008_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.24 PD=1.3 PS=1.48 NRD=1.9503 NRS=37.4103 M=1 R=5.55556 SA=90000.8
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1004 A_546_297# N_B1_M1004_g N_A_227_297#_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=23.6203 NRS=1.9503 M=1 R=5.55556
+ SA=90001.3 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1000 N_A_80_21#_M1000_d N_C1_M1000_g A_546_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.175 PD=2.55 PS=1.35 NRD=1.9503 NRS=23.6203 M=1 R=5.55556
+ SA=90001.9 SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_14 B1 B1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a211o_1.pxi.spice"
*
.ends
*
*
