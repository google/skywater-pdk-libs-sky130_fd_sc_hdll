* File: sky130_fd_sc_hdll__a31oi_4.pxi.spice
* Created: Wed Sep  2 08:20:27 2020
* 
x_PM_SKY130_FD_SC_HDLL__A31OI_4%A3 N_A3_c_88_n N_A3_M1001_g N_A3_c_83_n
+ N_A3_M1002_g N_A3_c_89_n N_A3_M1012_g N_A3_c_84_n N_A3_M1022_g N_A3_c_90_n
+ N_A3_M1021_g N_A3_c_85_n N_A3_M1023_g N_A3_c_91_n N_A3_M1030_g N_A3_c_86_n
+ N_A3_M1031_g A3 A3 A3 A3 N_A3_c_87_n A3 A3 PM_SKY130_FD_SC_HDLL__A31OI_4%A3
x_PM_SKY130_FD_SC_HDLL__A31OI_4%A2 N_A2_c_157_n N_A2_M1010_g N_A2_c_163_n
+ N_A2_M1000_g N_A2_c_158_n N_A2_M1018_g N_A2_c_164_n N_A2_M1003_g N_A2_c_159_n
+ N_A2_M1026_g N_A2_c_165_n N_A2_M1008_g N_A2_c_166_n N_A2_M1017_g N_A2_c_160_n
+ N_A2_M1028_g A2 A2 A2 A2 N_A2_c_161_n A2 A2 A2 A2
+ PM_SKY130_FD_SC_HDLL__A31OI_4%A2
x_PM_SKY130_FD_SC_HDLL__A31OI_4%A1 N_A1_c_238_n N_A1_M1004_g N_A1_c_239_n
+ N_A1_M1011_g N_A1_c_231_n N_A1_M1007_g N_A1_c_240_n N_A1_M1024_g N_A1_c_232_n
+ N_A1_M1013_g N_A1_c_241_n N_A1_M1025_g N_A1_c_233_n N_A1_M1027_g N_A1_c_234_n
+ N_A1_c_235_n N_A1_c_236_n N_A1_M1029_g A1 A1 A1 A1 A1 A1 A1 A1
+ PM_SKY130_FD_SC_HDLL__A31OI_4%A1
x_PM_SKY130_FD_SC_HDLL__A31OI_4%B1 N_B1_c_313_n N_B1_M1005_g N_B1_c_307_n
+ N_B1_M1006_g N_B1_c_314_n N_B1_M1009_g N_B1_c_308_n N_B1_M1014_g N_B1_c_315_n
+ N_B1_M1015_g N_B1_c_309_n N_B1_M1016_g N_B1_c_316_n N_B1_M1020_g N_B1_c_310_n
+ N_B1_M1019_g B1 B1 B1 N_B1_c_312_n B1 B1 B1 PM_SKY130_FD_SC_HDLL__A31OI_4%B1
x_PM_SKY130_FD_SC_HDLL__A31OI_4%A_27_297# N_A_27_297#_M1001_d
+ N_A_27_297#_M1012_d N_A_27_297#_M1030_d N_A_27_297#_M1003_d
+ N_A_27_297#_M1017_d N_A_27_297#_M1011_d N_A_27_297#_M1025_d
+ N_A_27_297#_M1009_d N_A_27_297#_M1020_d N_A_27_297#_c_384_n
+ N_A_27_297#_c_385_n N_A_27_297#_c_389_n N_A_27_297#_c_391_n
+ N_A_27_297#_c_393_n N_A_27_297#_c_397_n N_A_27_297#_c_401_n
+ N_A_27_297#_c_405_n N_A_27_297#_c_407_n N_A_27_297#_c_411_n
+ N_A_27_297#_c_417_n N_A_27_297#_c_421_n N_A_27_297#_c_423_n
+ N_A_27_297#_c_427_n N_A_27_297#_c_435_n N_A_27_297#_c_440_n
+ N_A_27_297#_c_470_p N_A_27_297#_c_497_p N_A_27_297#_c_398_n
+ N_A_27_297#_c_412_n N_A_27_297#_c_413_n N_A_27_297#_c_415_n
+ N_A_27_297#_c_428_n PM_SKY130_FD_SC_HDLL__A31OI_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A31OI_4%VPWR N_VPWR_M1001_s N_VPWR_M1021_s
+ N_VPWR_M1000_s N_VPWR_M1008_s N_VPWR_M1004_s N_VPWR_M1024_s N_VPWR_c_500_n
+ N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n
+ N_VPWR_c_506_n VPWR N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_499_n N_VPWR_c_513_n N_VPWR_c_514_n
+ N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n
+ PM_SKY130_FD_SC_HDLL__A31OI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A31OI_4%Y N_Y_M1007_d N_Y_M1013_d N_Y_M1029_d
+ N_Y_M1014_d N_Y_M1019_d N_Y_M1005_s N_Y_M1015_s N_Y_c_626_n N_Y_c_641_n
+ N_Y_c_646_n N_Y_c_647_n N_Y_c_650_n N_Y_c_684_p N_Y_c_651_n Y Y Y Y
+ N_Y_c_654_n Y Y PM_SKY130_FD_SC_HDLL__A31OI_4%Y
x_PM_SKY130_FD_SC_HDLL__A31OI_4%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1022_d
+ N_A_27_47#_M1031_d N_A_27_47#_M1018_d N_A_27_47#_M1028_d N_A_27_47#_c_703_n
+ N_A_27_47#_c_704_n N_A_27_47#_c_708_n N_A_27_47#_c_710_n N_A_27_47#_c_711_n
+ N_A_27_47#_c_729_p N_A_27_47#_c_702_n N_A_27_47#_c_715_n N_A_27_47#_c_723_n
+ PM_SKY130_FD_SC_HDLL__A31OI_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__A31OI_4%VGND N_VGND_M1002_s N_VGND_M1023_s
+ N_VGND_M1006_s N_VGND_M1016_s N_VGND_c_756_n N_VGND_c_757_n N_VGND_c_758_n
+ N_VGND_c_759_n VGND N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n
+ N_VGND_c_763_n N_VGND_c_764_n N_VGND_c_765_n
+ PM_SKY130_FD_SC_HDLL__A31OI_4%VGND
x_PM_SKY130_FD_SC_HDLL__A31OI_4%A_485_47# N_A_485_47#_M1010_s
+ N_A_485_47#_M1026_s N_A_485_47#_M1007_s N_A_485_47#_M1027_s
+ N_A_485_47#_c_867_n PM_SKY130_FD_SC_HDLL__A31OI_4%A_485_47#
cc_1 VNB N_A3_c_83_n 0.0219558f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_A3_c_84_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_A3_c_85_n 0.0164634f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_4 VNB N_A3_c_86_n 0.0167331f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_A3_c_87_n 0.105734f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_6 VNB N_A2_c_157_n 0.0167331f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_7 VNB N_A2_c_158_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_8 VNB N_A2_c_159_n 0.0174167f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_9 VNB N_A2_c_160_n 0.0229091f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_10 VNB N_A2_c_161_n 0.0726796f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_11 VNB A2 0.00637804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A1_c_231_n 0.022465f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_13 VNB N_A1_c_232_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_14 VNB N_A1_c_233_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_15 VNB N_A1_c_234_n 0.0213478f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_16 VNB N_A1_c_235_n 0.086138f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_17 VNB N_A1_c_236_n 0.0178636f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_18 VNB A1 0.00159364f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B1_c_307_n 0.0166804f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_20 VNB N_B1_c_308_n 0.0169689f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_21 VNB N_B1_c_309_n 0.0164213f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_22 VNB N_B1_c_310_n 0.0219898f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_23 VNB B1 0.00205078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_B1_c_312_n 0.0887686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_499_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_626_n 0.00223563f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_27 VNB Y 0.0010588f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_702_n 0.0031452f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_29 VNB N_VGND_c_756_n 0.00792095f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_30 VNB N_VGND_c_757_n 0.115994f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_31 VNB N_VGND_c_758_n 0.00849831f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_32 VNB N_VGND_c_759_n 0.0134288f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_33 VNB N_VGND_c_760_n 0.0151574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_761_n 0.0134288f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_35 VNB N_VGND_c_762_n 0.0217207f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_36 VNB N_VGND_c_763_n 0.418884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_764_n 0.00792095f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=1.16
cc_38 VNB N_VGND_c_765_n 0.00849831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_485_47#_c_867_n 0.00782917f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_40 VPB N_A3_c_88_n 0.0206372f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_41 VPB N_A3_c_89_n 0.0160921f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_42 VPB N_A3_c_90_n 0.0158129f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_43 VPB N_A3_c_91_n 0.0162737f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_44 VPB N_A3_c_87_n 0.0581273f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_45 VPB N_A2_c_163_n 0.0159944f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_46 VPB N_A2_c_164_n 0.0160921f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_47 VPB N_A2_c_165_n 0.0158129f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_48 VPB N_A2_c_166_n 0.016429f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_49 VPB N_A2_c_161_n 0.0453899f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_50 VPB A2 0.0021736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A1_c_238_n 0.0161497f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_52 VPB N_A1_c_239_n 0.0160921f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_53 VPB N_A1_c_240_n 0.0158129f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_54 VPB N_A1_c_241_n 0.0194863f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_55 VPB N_A1_c_234_n 0.0207701f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_56 VPB N_A1_c_235_n 0.0479333f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_57 VPB N_B1_c_313_n 0.0192858f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_58 VPB N_B1_c_314_n 0.0155986f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_59 VPB N_B1_c_315_n 0.0159124f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_60 VPB N_B1_c_316_n 0.0207585f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_61 VPB B1 0.00240873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_B1_c_312_n 0.0535688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_500_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_64 VPB N_VPWR_c_501_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_65 VPB N_VPWR_c_502_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_503_n 3.22956e-19 $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.202
cc_67 VPB N_VPWR_c_504_n 0.014719f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_68 VPB N_VPWR_c_505_n 3.22956e-19 $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_69 VPB N_VPWR_c_506_n 0.0141085f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.202
cc_70 VPB N_VPWR_c_507_n 0.0159043f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_71 VPB N_VPWR_c_508_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.16
cc_72 VPB N_VPWR_c_509_n 0.0140826f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=1.16
cc_73 VPB N_VPWR_c_510_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_511_n 0.0771679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_499_n 0.0511754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_513_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_514_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_515_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_516_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_517_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_518_n 0.0054644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB Y 0.00105149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 N_A3_c_86_n N_A2_c_157_n 0.0229653f $X=1.93 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_84 N_A3_c_91_n N_A2_c_163_n 0.0213451f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A3_c_87_n N_A2_c_161_n 0.0229653f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_86 A3 N_A2_c_161_n 2.79436e-19 $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_87 N_A3_c_87_n A2 0.00317941f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_88 A3 A2 0.021867f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_89 N_A3_c_88_n N_A_27_297#_c_384_n 0.00836571f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A3_c_88_n N_A_27_297#_c_385_n 0.0166293f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A3_c_89_n N_A_27_297#_c_385_n 0.0168429f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A3_c_87_n N_A_27_297#_c_385_n 0.00635951f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_93 A3 N_A_27_297#_c_385_n 0.0474842f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_94 N_A3_c_87_n N_A_27_297#_c_389_n 0.00396026f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_95 A3 N_A_27_297#_c_389_n 0.0140387f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_96 N_A3_c_89_n N_A_27_297#_c_391_n 0.00722591f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A3_c_90_n N_A_27_297#_c_391_n 0.00682765f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A3_c_90_n N_A_27_297#_c_393_n 0.0155135f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A3_c_91_n N_A_27_297#_c_393_n 0.0202024f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A3_c_87_n N_A_27_297#_c_393_n 0.00635951f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_101 A3 N_A_27_297#_c_393_n 0.0373774f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_102 N_A3_c_91_n N_A_27_297#_c_397_n 0.00722591f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A3_c_87_n N_A_27_297#_c_398_n 0.00411803f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_104 A3 N_A_27_297#_c_398_n 0.0140387f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_105 N_A3_c_88_n N_VPWR_c_500_n 0.0161957f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A3_c_89_n N_VPWR_c_500_n 0.0108266f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A3_c_90_n N_VPWR_c_500_n 5.96427e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A3_c_89_n N_VPWR_c_501_n 6.33692e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A3_c_90_n N_VPWR_c_501_n 0.0144185f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A3_c_91_n N_VPWR_c_501_n 0.0108266f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A3_c_91_n N_VPWR_c_502_n 6.33692e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A3_c_88_n N_VPWR_c_507_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A3_c_89_n N_VPWR_c_508_n 0.00622633f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A3_c_90_n N_VPWR_c_508_n 0.00427505f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A3_c_91_n N_VPWR_c_509_n 0.00622633f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A3_c_88_n N_VPWR_c_499_n 0.0082412f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A3_c_89_n N_VPWR_c_499_n 0.0104011f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A3_c_90_n N_VPWR_c_499_n 0.00732977f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A3_c_91_n N_VPWR_c_499_n 0.0104264f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A3_c_83_n N_A_27_47#_c_703_n 0.00405771f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A3_c_83_n N_A_27_47#_c_704_n 0.0127563f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A3_c_84_n N_A_27_47#_c_704_n 0.0124611f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A3_c_87_n N_A_27_47#_c_704_n 0.00534082f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_124 A3 N_A_27_47#_c_704_n 0.0440221f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_125 N_A3_c_87_n N_A_27_47#_c_708_n 0.00388817f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_126 A3 N_A_27_47#_c_708_n 0.0126663f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_127 N_A3_c_85_n N_A_27_47#_c_710_n 0.00377939f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A3_c_85_n N_A_27_47#_c_711_n 0.0116963f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A3_c_86_n N_A_27_47#_c_711_n 0.0156709f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A3_c_87_n N_A_27_47#_c_711_n 0.00331732f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_131 A3 N_A_27_47#_c_711_n 0.034467f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_132 N_A3_c_87_n N_A_27_47#_c_715_n 0.00297321f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_133 A3 N_A_27_47#_c_715_n 0.0123849f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_134 N_A3_c_86_n N_VGND_c_757_n 0.00425094f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A3_c_83_n N_VGND_c_760_n 0.00198377f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A3_c_84_n N_VGND_c_761_n 0.00425094f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A3_c_85_n N_VGND_c_761_n 0.00198377f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A3_c_83_n N_VGND_c_763_n 0.00358947f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A3_c_84_n N_VGND_c_763_n 0.00584696f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A3_c_85_n N_VGND_c_763_n 0.00271758f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A3_c_86_n N_VGND_c_763_n 0.0057472f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A3_c_83_n N_VGND_c_764_n 0.0112154f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A3_c_84_n N_VGND_c_764_n 0.00162962f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A3_c_84_n N_VGND_c_765_n 5.64511e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A3_c_85_n N_VGND_c_765_n 0.00960147f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A3_c_86_n N_VGND_c_765_n 0.00317372f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A2_c_166_n N_A1_c_238_n 0.0197305f $X=3.785 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_148 N_A2_c_161_n N_A1_c_235_n 0.0191054f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_149 A2 N_A1_c_235_n 0.00284587f $X=3.875 $Y=1.19 $X2=0 $Y2=0
cc_150 N_A2_c_161_n A1 3.47199e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_151 A2 A1 0.0203714f $X=3.875 $Y=1.19 $X2=0 $Y2=0
cc_152 N_A2_c_163_n N_A_27_297#_c_397_n 0.00682765f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A2_c_163_n N_A_27_297#_c_401_n 0.0154704f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_c_164_n N_A_27_297#_c_401_n 0.016886f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A2_c_161_n N_A_27_297#_c_401_n 0.00635951f $X=3.785 $Y=1.202 $X2=0
+ $Y2=0
cc_156 A2 N_A_27_297#_c_401_n 0.0476898f $X=3.875 $Y=1.19 $X2=0 $Y2=0
cc_157 N_A2_c_164_n N_A_27_297#_c_405_n 0.00722591f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A2_c_165_n N_A_27_297#_c_405_n 0.00682765f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A2_c_165_n N_A_27_297#_c_407_n 0.0155135f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A2_c_166_n N_A_27_297#_c_407_n 0.0169558f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A2_c_161_n N_A_27_297#_c_407_n 0.00616252f $X=3.785 $Y=1.202 $X2=0
+ $Y2=0
cc_162 A2 N_A_27_297#_c_407_n 0.0476898f $X=3.875 $Y=1.19 $X2=0 $Y2=0
cc_163 N_A2_c_166_n N_A_27_297#_c_411_n 0.00725278f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_164 A2 N_A_27_297#_c_412_n 0.00780217f $X=3.875 $Y=1.19 $X2=0 $Y2=0
cc_165 N_A2_c_161_n N_A_27_297#_c_413_n 0.00411803f $X=3.785 $Y=1.202 $X2=0
+ $Y2=0
cc_166 A2 N_A_27_297#_c_413_n 0.0140387f $X=3.875 $Y=1.19 $X2=0 $Y2=0
cc_167 A2 N_A_27_297#_c_415_n 0.00130036f $X=3.875 $Y=1.19 $X2=0 $Y2=0
cc_168 N_A2_c_163_n N_VPWR_c_501_n 5.96427e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A2_c_163_n N_VPWR_c_502_n 0.0144185f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A2_c_164_n N_VPWR_c_502_n 0.0108266f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A2_c_165_n N_VPWR_c_502_n 5.96427e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A2_c_164_n N_VPWR_c_503_n 6.33692e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A2_c_165_n N_VPWR_c_503_n 0.0144185f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A2_c_166_n N_VPWR_c_503_n 0.0108937f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A2_c_166_n N_VPWR_c_504_n 0.00622633f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A2_c_166_n N_VPWR_c_505_n 6.38483e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A2_c_163_n N_VPWR_c_509_n 0.00427505f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A2_c_164_n N_VPWR_c_510_n 0.00622633f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A2_c_165_n N_VPWR_c_510_n 0.00427505f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A2_c_163_n N_VPWR_c_499_n 0.00735499f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A2_c_164_n N_VPWR_c_499_n 0.0104011f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A2_c_165_n N_VPWR_c_499_n 0.00732977f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A2_c_166_n N_VPWR_c_499_n 0.0104733f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A2_c_157_n N_A_27_47#_c_702_n 0.0118402f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A2_c_158_n N_A_27_47#_c_702_n 0.0087742f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A2_c_159_n N_A_27_47#_c_702_n 0.00903316f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A2_c_160_n N_A_27_47#_c_702_n 0.00903316f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A2_c_161_n N_A_27_47#_c_702_n 0.0104016f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_189 A2 N_A_27_47#_c_702_n 0.1008f $X=3.875 $Y=1.19 $X2=0 $Y2=0
cc_190 A2 N_A_27_47#_c_723_n 0.00680018f $X=3.875 $Y=1.19 $X2=0 $Y2=0
cc_191 N_A2_c_157_n N_VGND_c_757_n 0.00413298f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_158_n N_VGND_c_757_n 0.00366111f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A2_c_159_n N_VGND_c_757_n 0.00366111f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_160_n N_VGND_c_757_n 0.00366111f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A2_c_157_n N_VGND_c_763_n 0.0058296f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_c_158_n N_VGND_c_763_n 0.00549891f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A2_c_159_n N_VGND_c_763_n 0.00561425f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_c_160_n N_VGND_c_763_n 0.00685947f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A2_c_157_n N_A_485_47#_c_867_n 0.00245853f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A2_c_158_n N_A_485_47#_c_867_n 0.00818766f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A2_c_159_n N_A_485_47#_c_867_n 0.00818766f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A2_c_160_n N_A_485_47#_c_867_n 0.00999448f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A1_c_236_n N_B1_c_307_n 0.0215122f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_204 N_A1_c_241_n B1 0.00312031f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A1_c_234_n B1 0.01172f $X=6.185 $Y=1.167 $X2=0 $Y2=0
cc_206 N_A1_c_235_n B1 0.00268011f $X=5.865 $Y=1.167 $X2=0 $Y2=0
cc_207 N_A1_c_236_n B1 0.00130751f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_208 A1 B1 0.0203743f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_209 N_A1_c_236_n N_B1_c_312_n 0.0215549f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_210 N_A1_c_238_n N_A_27_297#_c_411_n 0.0068226f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A1_c_238_n N_A_27_297#_c_417_n 0.0167067f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A1_c_239_n N_A_27_297#_c_417_n 0.016886f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A1_c_235_n N_A_27_297#_c_417_n 0.00605803f $X=5.865 $Y=1.167 $X2=0
+ $Y2=0
cc_214 A1 N_A_27_297#_c_417_n 0.0423763f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_215 N_A1_c_239_n N_A_27_297#_c_421_n 0.00722591f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A1_c_240_n N_A_27_297#_c_421_n 0.0125395f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A1_c_240_n N_A_27_297#_c_423_n 0.0161777f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A1_c_241_n N_A_27_297#_c_423_n 0.0170288f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A1_c_235_n N_A_27_297#_c_423_n 0.0110937f $X=5.865 $Y=1.167 $X2=0 $Y2=0
cc_220 A1 N_A_27_297#_c_423_n 0.0614851f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_221 N_A1_c_241_n N_A_27_297#_c_427_n 0.0136792f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A1_c_235_n N_A_27_297#_c_428_n 0.00455443f $X=5.865 $Y=1.167 $X2=0
+ $Y2=0
cc_223 A1 N_A_27_297#_c_428_n 0.0140387f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_224 N_A1_c_238_n N_VPWR_c_503_n 5.8529e-19 $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A1_c_238_n N_VPWR_c_504_n 0.00427505f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A1_c_238_n N_VPWR_c_505_n 0.0147392f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A1_c_239_n N_VPWR_c_505_n 0.0108266f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A1_c_240_n N_VPWR_c_505_n 5.96427e-19 $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A1_c_239_n N_VPWR_c_506_n 0.00622633f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A1_c_240_n N_VPWR_c_506_n 0.00429282f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A1_c_241_n N_VPWR_c_511_n 0.0062441f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A1_c_238_n N_VPWR_c_499_n 0.00740194f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A1_c_239_n N_VPWR_c_499_n 0.0104011f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A1_c_240_n N_VPWR_c_499_n 0.00732982f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A1_c_241_n N_VPWR_c_499_n 0.0116835f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A1_c_239_n N_VPWR_c_518_n 5.36535e-19 $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A1_c_240_n N_VPWR_c_518_n 0.0103971f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_238 N_A1_c_241_n N_VPWR_c_518_n 0.00861566f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A1_c_231_n N_Y_c_626_n 0.0087742f $X=4.85 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A1_c_232_n N_Y_c_626_n 0.0087742f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A1_c_233_n N_Y_c_626_n 0.0087742f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A1_c_234_n N_Y_c_626_n 0.00312844f $X=6.185 $Y=1.167 $X2=0 $Y2=0
cc_243 N_A1_c_235_n N_Y_c_626_n 0.0146477f $X=5.865 $Y=1.167 $X2=0 $Y2=0
cc_244 N_A1_c_236_n N_Y_c_626_n 0.0124981f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_245 A1 N_Y_c_626_n 0.0961563f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_246 N_A1_c_235_n N_A_27_47#_c_702_n 3.7827e-19 $X=5.865 $Y=1.167 $X2=0 $Y2=0
cc_247 N_A1_c_236_n N_VGND_c_756_n 0.00197423f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_248 N_A1_c_231_n N_VGND_c_757_n 0.00366111f $X=4.85 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A1_c_232_n N_VGND_c_757_n 0.00366111f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A1_c_233_n N_VGND_c_757_n 0.00366111f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A1_c_236_n N_VGND_c_757_n 0.00425094f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_252 N_A1_c_231_n N_VGND_c_763_n 0.00674413f $X=4.85 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A1_c_232_n N_VGND_c_763_n 0.00549891f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A1_c_233_n N_VGND_c_763_n 0.00549891f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A1_c_236_n N_VGND_c_763_n 0.00611197f $X=6.26 $Y=1.01 $X2=0 $Y2=0
cc_256 N_A1_c_231_n N_A_485_47#_c_867_n 0.00999448f $X=4.85 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A1_c_232_n N_A_485_47#_c_867_n 0.00818766f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A1_c_233_n N_A_485_47#_c_867_n 0.00818766f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A1_c_235_n N_A_485_47#_c_867_n 0.0052885f $X=5.865 $Y=1.167 $X2=0 $Y2=0
cc_260 A1 N_A_485_47#_c_867_n 0.00638061f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_261 B1 N_A_27_297#_M1025_d 0.00898198f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_262 B1 N_A_27_297#_M1009_d 0.00247586f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_263 N_B1_c_313_n N_A_27_297#_c_423_n 0.00149132f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_264 B1 N_A_27_297#_c_423_n 0.00868458f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_265 N_B1_c_313_n N_A_27_297#_c_427_n 0.0130457f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B1_c_313_n N_A_27_297#_c_435_n 0.01488f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B1_c_314_n N_A_27_297#_c_435_n 0.0092122f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_268 N_B1_c_315_n N_A_27_297#_c_435_n 0.0092122f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_269 N_B1_c_316_n N_A_27_297#_c_435_n 0.0128305f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_270 B1 N_A_27_297#_c_435_n 0.0115539f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_271 N_B1_c_313_n N_A_27_297#_c_440_n 8.88013e-19 $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B1_c_313_n N_VPWR_c_511_n 0.00439333f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B1_c_314_n N_VPWR_c_511_n 0.00439333f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B1_c_315_n N_VPWR_c_511_n 0.00439333f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B1_c_316_n N_VPWR_c_511_n 0.00439333f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B1_c_313_n N_VPWR_c_499_n 0.00745558f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B1_c_314_n N_VPWR_c_499_n 0.00608292f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_278 N_B1_c_315_n N_VPWR_c_499_n 0.00608292f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B1_c_316_n N_VPWR_c_499_n 0.00709469f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_280 B1 N_Y_M1005_s 0.00247586f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_281 N_B1_c_307_n N_Y_c_626_n 0.00940277f $X=6.73 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B1_c_308_n N_Y_c_626_n 0.0124611f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_283 B1 N_Y_c_626_n 0.0660108f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_284 N_B1_c_312_n N_Y_c_626_n 0.00556447f $X=8.115 $Y=1.202 $X2=0 $Y2=0
cc_285 N_B1_c_313_n N_Y_c_641_n 0.0107672f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_286 N_B1_c_314_n N_Y_c_641_n 0.0105592f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_287 N_B1_c_315_n N_Y_c_641_n 0.0139313f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_288 B1 N_Y_c_641_n 0.0342985f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_289 N_B1_c_312_n N_Y_c_641_n 0.00375084f $X=8.115 $Y=1.202 $X2=0 $Y2=0
cc_290 N_B1_c_309_n N_Y_c_646_n 0.00377939f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B1_c_309_n N_Y_c_647_n 0.0157858f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_292 B1 N_Y_c_647_n 0.00588732f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_293 N_B1_c_312_n N_Y_c_647_n 5.6965e-19 $X=8.115 $Y=1.202 $X2=0 $Y2=0
cc_294 N_B1_c_310_n N_Y_c_650_n 0.0138332f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_295 B1 N_Y_c_651_n 0.0130015f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_296 N_B1_c_312_n N_Y_c_651_n 0.00297321f $X=8.115 $Y=1.202 $X2=0 $Y2=0
cc_297 N_B1_c_310_n Y 0.00304421f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_298 N_B1_c_316_n N_Y_c_654_n 0.00323163f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_299 N_B1_c_315_n Y 0.00810477f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_300 N_B1_c_309_n Y 0.00464444f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B1_c_316_n Y 0.0130059f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_302 N_B1_c_310_n Y 0.0096592f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_303 B1 Y 0.0384183f $X=7.435 $Y=1.105 $X2=0 $Y2=0
cc_304 N_B1_c_312_n Y 0.0383457f $X=8.115 $Y=1.202 $X2=0 $Y2=0
cc_305 N_B1_c_307_n N_VGND_c_756_n 0.0124455f $X=6.73 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B1_c_308_n N_VGND_c_756_n 0.00162962f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B1_c_307_n N_VGND_c_757_n 0.00198377f $X=6.73 $Y=0.995 $X2=0 $Y2=0
cc_308 N_B1_c_308_n N_VGND_c_758_n 5.64511e-19 $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_309 N_B1_c_309_n N_VGND_c_758_n 0.00960147f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_310 N_B1_c_310_n N_VGND_c_758_n 0.00317372f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_311 N_B1_c_312_n N_VGND_c_758_n 4.99612e-19 $X=8.115 $Y=1.202 $X2=0 $Y2=0
cc_312 N_B1_c_308_n N_VGND_c_759_n 0.00425094f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_313 N_B1_c_309_n N_VGND_c_759_n 0.00198377f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_314 N_B1_c_310_n N_VGND_c_762_n 0.00425075f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_315 N_B1_c_307_n N_VGND_c_763_n 0.00278437f $X=6.73 $Y=0.995 $X2=0 $Y2=0
cc_316 N_B1_c_308_n N_VGND_c_763_n 0.00584696f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B1_c_309_n N_VGND_c_763_n 0.00271758f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B1_c_310_n N_VGND_c_763_n 0.00677732f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_27_297#_c_385_n N_VPWR_M1001_s 0.00369624f $X=1.115 $Y=1.58 $X2=0.495
+ $Y2=1.41
cc_320 N_A_27_297#_c_393_n N_VPWR_M1021_s 0.00369624f $X=2.055 $Y=1.58 $X2=0.495
+ $Y2=1.985
cc_321 N_A_27_297#_c_401_n N_VPWR_M1000_s 0.00369624f $X=2.995 $Y=1.58 $X2=0.495
+ $Y2=1.985
cc_322 N_A_27_297#_c_407_n N_VPWR_M1008_s 0.00369624f $X=3.935 $Y=1.58 $X2=0.52
+ $Y2=0.995
cc_323 N_A_27_297#_c_417_n N_VPWR_M1004_s 0.00368674f $X=4.895 $Y=1.58 $X2=0.52
+ $Y2=0.56
cc_324 N_A_27_297#_c_423_n N_VPWR_M1024_s 0.00493294f $X=5.835 $Y=1.58 $X2=0.52
+ $Y2=0.56
cc_325 N_A_27_297#_c_384_n N_VPWR_c_500_n 0.0410603f $X=0.26 $Y=1.96 $X2=1.905
+ $Y2=1.985
cc_326 N_A_27_297#_c_385_n N_VPWR_c_500_n 0.0156171f $X=1.115 $Y=1.58 $X2=1.905
+ $Y2=1.985
cc_327 N_A_27_297#_c_391_n N_VPWR_c_500_n 0.0336646f $X=1.2 $Y=1.96 $X2=1.905
+ $Y2=1.985
cc_328 N_A_27_297#_c_391_n N_VPWR_c_501_n 0.0410603f $X=1.2 $Y=1.96 $X2=0.15
+ $Y2=1.105
cc_329 N_A_27_297#_c_393_n N_VPWR_c_501_n 0.0156171f $X=2.055 $Y=1.58 $X2=0.15
+ $Y2=1.105
cc_330 N_A_27_297#_c_397_n N_VPWR_c_501_n 0.0336646f $X=2.14 $Y=1.96 $X2=0.15
+ $Y2=1.105
cc_331 N_A_27_297#_c_397_n N_VPWR_c_502_n 0.0410603f $X=2.14 $Y=1.96 $X2=0 $Y2=0
cc_332 N_A_27_297#_c_401_n N_VPWR_c_502_n 0.0156171f $X=2.995 $Y=1.58 $X2=0
+ $Y2=0
cc_333 N_A_27_297#_c_405_n N_VPWR_c_502_n 0.0336646f $X=3.08 $Y=1.96 $X2=0 $Y2=0
cc_334 N_A_27_297#_c_405_n N_VPWR_c_503_n 0.0410603f $X=3.08 $Y=1.96 $X2=0.285
+ $Y2=1.202
cc_335 N_A_27_297#_c_407_n N_VPWR_c_503_n 0.0156171f $X=3.935 $Y=1.58 $X2=0.285
+ $Y2=1.202
cc_336 N_A_27_297#_c_411_n N_VPWR_c_503_n 0.0336646f $X=4.02 $Y=1.96 $X2=0.285
+ $Y2=1.202
cc_337 N_A_27_297#_c_411_n N_VPWR_c_504_n 0.0118139f $X=4.02 $Y=1.96 $X2=0.285
+ $Y2=1.16
cc_338 N_A_27_297#_c_411_n N_VPWR_c_505_n 0.0376795f $X=4.02 $Y=1.96 $X2=0.99
+ $Y2=1.202
cc_339 N_A_27_297#_c_417_n N_VPWR_c_505_n 0.0156171f $X=4.895 $Y=1.58 $X2=0.99
+ $Y2=1.202
cc_340 N_A_27_297#_c_421_n N_VPWR_c_505_n 0.0336646f $X=4.98 $Y=1.96 $X2=0.99
+ $Y2=1.202
cc_341 N_A_27_297#_c_421_n N_VPWR_c_506_n 0.0118139f $X=4.98 $Y=1.96 $X2=1.46
+ $Y2=1.202
cc_342 N_A_27_297#_c_384_n N_VPWR_c_507_n 0.0118139f $X=0.26 $Y=1.96 $X2=1.905
+ $Y2=1.202
cc_343 N_A_27_297#_c_391_n N_VPWR_c_508_n 0.0118139f $X=1.2 $Y=1.96 $X2=0.695
+ $Y2=1.16
cc_344 N_A_27_297#_c_397_n N_VPWR_c_509_n 0.0118139f $X=2.14 $Y=1.96 $X2=1.495
+ $Y2=1.16
cc_345 N_A_27_297#_c_405_n N_VPWR_c_510_n 0.0118139f $X=3.08 $Y=1.96 $X2=0 $Y2=0
cc_346 N_A_27_297#_c_435_n N_VPWR_c_511_n 0.102887f $X=8.265 $Y=2.34 $X2=0 $Y2=0
cc_347 N_A_27_297#_c_440_n N_VPWR_c_511_n 0.0119545f $X=6.005 $Y=2.34 $X2=0
+ $Y2=0
cc_348 N_A_27_297#_c_470_p N_VPWR_c_511_n 0.0139745f $X=8.39 $Y=2.255 $X2=0
+ $Y2=0
cc_349 N_A_27_297#_M1001_d N_VPWR_c_499_n 0.00568146f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_350 N_A_27_297#_M1012_d N_VPWR_c_499_n 0.00647849f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_351 N_A_27_297#_M1030_d N_VPWR_c_499_n 0.00647849f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_352 N_A_27_297#_M1003_d N_VPWR_c_499_n 0.00647849f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_353 N_A_27_297#_M1017_d N_VPWR_c_499_n 0.0073334f $X=3.875 $Y=1.485 $X2=0
+ $Y2=0
cc_354 N_A_27_297#_M1011_d N_VPWR_c_499_n 0.00647849f $X=4.835 $Y=1.485 $X2=0
+ $Y2=0
cc_355 N_A_27_297#_M1025_d N_VPWR_c_499_n 0.00892095f $X=5.775 $Y=1.485 $X2=0
+ $Y2=0
cc_356 N_A_27_297#_M1009_d N_VPWR_c_499_n 0.00233855f $X=7.265 $Y=1.485 $X2=0
+ $Y2=0
cc_357 N_A_27_297#_M1020_d N_VPWR_c_499_n 0.00338835f $X=8.205 $Y=1.485 $X2=0
+ $Y2=0
cc_358 N_A_27_297#_c_384_n N_VPWR_c_499_n 0.00646998f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_359 N_A_27_297#_c_391_n N_VPWR_c_499_n 0.00646998f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_360 N_A_27_297#_c_397_n N_VPWR_c_499_n 0.00646998f $X=2.14 $Y=1.96 $X2=0
+ $Y2=0
cc_361 N_A_27_297#_c_405_n N_VPWR_c_499_n 0.00646998f $X=3.08 $Y=1.96 $X2=0
+ $Y2=0
cc_362 N_A_27_297#_c_411_n N_VPWR_c_499_n 0.00646998f $X=4.02 $Y=1.96 $X2=0
+ $Y2=0
cc_363 N_A_27_297#_c_421_n N_VPWR_c_499_n 0.00646998f $X=4.98 $Y=1.96 $X2=0
+ $Y2=0
cc_364 N_A_27_297#_c_435_n N_VPWR_c_499_n 0.0785579f $X=8.265 $Y=2.34 $X2=0
+ $Y2=0
cc_365 N_A_27_297#_c_440_n N_VPWR_c_499_n 0.006547f $X=6.005 $Y=2.34 $X2=0 $Y2=0
cc_366 N_A_27_297#_c_470_p N_VPWR_c_499_n 0.00943767f $X=8.39 $Y=2.255 $X2=0
+ $Y2=0
cc_367 N_A_27_297#_c_421_n N_VPWR_c_518_n 0.0156776f $X=4.98 $Y=1.96 $X2=0 $Y2=0
cc_368 N_A_27_297#_c_423_n N_VPWR_c_518_n 0.00786103f $X=5.835 $Y=1.58 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_440_n N_VPWR_c_518_n 0.0140804f $X=6.005 $Y=2.34 $X2=0
+ $Y2=0
cc_370 N_A_27_297#_c_435_n N_Y_M1005_s 0.00367601f $X=8.265 $Y=2.34 $X2=0.52
+ $Y2=0.56
cc_371 N_A_27_297#_c_435_n N_Y_M1015_s 0.00366219f $X=8.265 $Y=2.34 $X2=0.965
+ $Y2=1.41
cc_372 N_A_27_297#_M1009_d N_Y_c_641_n 0.00393624f $X=7.265 $Y=1.485 $X2=0 $Y2=0
cc_373 N_A_27_297#_c_435_n N_Y_c_641_n 0.0553837f $X=8.265 $Y=2.34 $X2=0 $Y2=0
cc_374 N_A_27_297#_c_435_n N_Y_c_654_n 0.0136488f $X=8.265 $Y=2.34 $X2=1.615
+ $Y2=1.19
cc_375 N_A_27_297#_c_497_p N_Y_c_654_n 0.0131326f $X=8.35 $Y=1.66 $X2=1.615
+ $Y2=1.19
cc_376 N_A_27_297#_c_497_p Y 0.0297883f $X=8.35 $Y=1.66 $X2=0 $Y2=0
cc_377 N_VPWR_c_499_n N_Y_M1005_s 0.00235479f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_378 N_VPWR_c_499_n N_Y_M1015_s 0.00235479f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_379 N_Y_c_626_n N_A_27_47#_c_702_n 0.0123435f $X=7.325 $Y=0.72 $X2=0 $Y2=0
cc_380 N_Y_c_626_n N_VGND_M1006_s 0.00407492f $X=7.325 $Y=0.72 $X2=0 $Y2=0
cc_381 N_Y_c_647_n N_VGND_M1016_s 0.00179449f $X=7.845 $Y=0.72 $X2=0 $Y2=0
cc_382 Y N_VGND_M1016_s 0.00173521f $X=7.895 $Y=0.765 $X2=0 $Y2=0
cc_383 Y N_VGND_M1016_s 9.18926e-19 $X=7.96 $Y=0.85 $X2=0 $Y2=0
cc_384 N_Y_c_626_n N_VGND_c_756_n 0.0213178f $X=7.325 $Y=0.72 $X2=0 $Y2=0
cc_385 N_Y_c_626_n N_VGND_c_757_n 0.00850371f $X=7.325 $Y=0.72 $X2=0 $Y2=0
cc_386 N_Y_c_646_n N_VGND_c_758_n 0.0156777f $X=7.41 $Y=0.42 $X2=0 $Y2=0
cc_387 N_Y_c_647_n N_VGND_c_758_n 0.00884855f $X=7.845 $Y=0.72 $X2=0 $Y2=0
cc_388 Y N_VGND_c_758_n 0.0137366f $X=7.895 $Y=0.765 $X2=0 $Y2=0
cc_389 N_Y_c_626_n N_VGND_c_759_n 0.00313948f $X=7.325 $Y=0.72 $X2=0 $Y2=0
cc_390 N_Y_c_646_n N_VGND_c_759_n 0.01143f $X=7.41 $Y=0.42 $X2=0 $Y2=0
cc_391 N_Y_c_647_n N_VGND_c_759_n 0.00244812f $X=7.845 $Y=0.72 $X2=0 $Y2=0
cc_392 N_Y_c_650_n N_VGND_c_762_n 0.00260993f $X=8.265 $Y=0.72 $X2=0 $Y2=0
cc_393 N_Y_c_684_p N_VGND_c_762_n 0.01143f $X=8.35 $Y=0.42 $X2=0 $Y2=0
cc_394 Y N_VGND_c_762_n 5.55499e-19 $X=7.895 $Y=0.765 $X2=0 $Y2=0
cc_395 N_Y_M1007_d N_VGND_c_763_n 0.00253905f $X=4.465 $Y=0.235 $X2=0 $Y2=0
cc_396 N_Y_M1013_d N_VGND_c_763_n 0.00259839f $X=5.395 $Y=0.235 $X2=0 $Y2=0
cc_397 N_Y_M1029_d N_VGND_c_763_n 0.00375565f $X=6.335 $Y=0.235 $X2=0 $Y2=0
cc_398 N_Y_M1014_d N_VGND_c_763_n 0.00309604f $X=7.275 $Y=0.235 $X2=0 $Y2=0
cc_399 N_Y_M1019_d N_VGND_c_763_n 0.00626209f $X=8.215 $Y=0.235 $X2=0 $Y2=0
cc_400 N_Y_c_626_n N_VGND_c_763_n 0.0249903f $X=7.325 $Y=0.72 $X2=0 $Y2=0
cc_401 N_Y_c_646_n N_VGND_c_763_n 0.00643448f $X=7.41 $Y=0.42 $X2=0 $Y2=0
cc_402 N_Y_c_647_n N_VGND_c_763_n 0.00521685f $X=7.845 $Y=0.72 $X2=0 $Y2=0
cc_403 N_Y_c_650_n N_VGND_c_763_n 0.00439883f $X=8.265 $Y=0.72 $X2=0 $Y2=0
cc_404 N_Y_c_684_p N_VGND_c_763_n 0.00643448f $X=8.35 $Y=0.42 $X2=0 $Y2=0
cc_405 Y N_VGND_c_763_n 0.00206408f $X=7.895 $Y=0.765 $X2=0 $Y2=0
cc_406 N_Y_c_626_n N_A_485_47#_M1007_s 0.00407984f $X=7.325 $Y=0.72 $X2=0 $Y2=0
cc_407 N_Y_c_626_n N_A_485_47#_M1027_s 0.00520574f $X=7.325 $Y=0.72 $X2=0 $Y2=0
cc_408 N_Y_M1007_d N_A_485_47#_c_867_n 0.00621528f $X=4.465 $Y=0.235 $X2=0 $Y2=0
cc_409 N_Y_M1013_d N_A_485_47#_c_867_n 0.00414886f $X=5.395 $Y=0.235 $X2=0 $Y2=0
cc_410 N_Y_c_626_n N_A_485_47#_c_867_n 0.0916483f $X=7.325 $Y=0.72 $X2=0 $Y2=0
cc_411 N_A_27_47#_c_704_n N_VGND_M1002_s 0.00407492f $X=1.115 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_412 N_A_27_47#_c_711_n N_VGND_M1023_s 0.00407492f $X=2.055 $Y=0.72 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_711_n N_VGND_c_757_n 0.00313948f $X=2.055 $Y=0.72 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_c_729_p N_VGND_c_757_n 0.0112274f $X=2.14 $Y=0.42 $X2=0 $Y2=0
cc_415 N_A_27_47#_c_702_n N_VGND_c_757_n 0.00245287f $X=4.02 $Y=0.72 $X2=0 $Y2=0
cc_416 N_A_27_47#_c_703_n N_VGND_c_760_n 0.0116326f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_417 N_A_27_47#_c_704_n N_VGND_c_760_n 0.00244812f $X=1.115 $Y=0.72 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_704_n N_VGND_c_761_n 0.00313948f $X=1.115 $Y=0.72 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_710_n N_VGND_c_761_n 0.01143f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_420 N_A_27_47#_c_711_n N_VGND_c_761_n 0.00244812f $X=2.055 $Y=0.72 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_M1002_d N_VGND_c_763_n 0.00430496f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_M1022_d N_VGND_c_763_n 0.00309604f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_M1031_d N_VGND_c_763_n 0.00249348f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_M1018_d N_VGND_c_763_n 0.00259839f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_M1028_d N_VGND_c_763_n 0.00212464f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_c_703_n N_VGND_c_763_n 0.00643448f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_427 N_A_27_47#_c_704_n N_VGND_c_763_n 0.0114934f $X=1.115 $Y=0.72 $X2=0 $Y2=0
cc_428 N_A_27_47#_c_710_n N_VGND_c_763_n 0.00643448f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_429 N_A_27_47#_c_711_n N_VGND_c_763_n 0.0114934f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_430 N_A_27_47#_c_729_p N_VGND_c_763_n 0.00643448f $X=2.14 $Y=0.42 $X2=0 $Y2=0
cc_431 N_A_27_47#_c_702_n N_VGND_c_763_n 0.00746781f $X=4.02 $Y=0.72 $X2=0 $Y2=0
cc_432 N_A_27_47#_c_703_n N_VGND_c_764_n 0.0156777f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_433 N_A_27_47#_c_704_n N_VGND_c_764_n 0.0213178f $X=1.115 $Y=0.72 $X2=0 $Y2=0
cc_434 N_A_27_47#_c_710_n N_VGND_c_765_n 0.0156777f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_435 N_A_27_47#_c_711_n N_VGND_c_765_n 0.0213178f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_436 N_A_27_47#_c_702_n N_A_485_47#_M1010_s 0.00407984f $X=4.02 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_437 N_A_27_47#_c_702_n N_A_485_47#_M1026_s 0.005125f $X=4.02 $Y=0.72 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_M1018_d N_A_485_47#_c_867_n 0.00414886f $X=2.895 $Y=0.235
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_M1028_d N_A_485_47#_c_867_n 0.00498385f $X=3.885 $Y=0.235
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_702_n N_A_485_47#_c_867_n 0.0935441f $X=4.02 $Y=0.72 $X2=0
+ $Y2=0
cc_441 N_VGND_c_763_n N_A_485_47#_M1010_s 0.00258215f $X=8.51 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_442 N_VGND_c_763_n N_A_485_47#_M1026_s 0.00298815f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_443 N_VGND_c_763_n N_A_485_47#_M1007_s 0.00258215f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_444 N_VGND_c_763_n N_A_485_47#_M1027_s 0.00264976f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_c_757_n N_A_485_47#_c_867_n 0.172142f $X=6.725 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_763_n N_A_485_47#_c_867_n 0.1322f $X=8.51 $Y=0 $X2=0 $Y2=0
