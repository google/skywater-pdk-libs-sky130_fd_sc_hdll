* NGSPICE file created from sky130_fd_sc_hdll__dlygate4sd3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__dlygate4sd3_1 A VGND VNB VPB VPWR X
M1000 VPWR a_273_47# a_379_93# VPB phighvt w=420000u l=500000u
+  ad=4.491e+11p pd=4.15e+06u as=1.092e+11p ps=1.36e+06u
M1001 X a_379_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1002 VPWR A a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_273_47# a_27_47# VGND VNB nshort w=420000u l=500000u
+  ad=1.092e+11p pd=1.36e+06u as=3.636e+11p ps=3.51e+06u
M1004 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1005 X a_379_93# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1006 VGND a_273_47# a_379_93# VNB nshort w=420000u l=500000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1007 a_273_47# a_27_47# VPWR VPB phighvt w=420000u l=500000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
.ends

