* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_521_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=2.6e+11p ps=2.1e+06u
M1001 a_119_47# A2_N a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=2.3e+11p ps=2.46e+06u
M1002 a_117_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.7e+11p ps=5.14e+06u
M1003 VGND A2_N a_119_47# VNB nshort w=650000u l=150000u
+  ad=9.425e+11p pd=6.8e+06u as=2.145e+11p ps=1.96e+06u
M1004 Y a_119_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_409_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.4e+11p pd=5.28e+06u as=0p ps=0u
M1006 a_409_297# a_119_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 a_119_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B1 a_521_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B2 a_409_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
