* File: sky130_fd_sc_hdll__and2_4.pxi.spice
* Created: Thu Aug 27 18:56:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND2_4%A N_A_c_55_n N_A_M1004_g N_A_c_56_n N_A_M1002_g A
+ N_A_c_57_n PM_SKY130_FD_SC_HDLL__AND2_4%A
x_PM_SKY130_FD_SC_HDLL__AND2_4%B N_B_c_78_n N_B_M1009_g N_B_c_79_n N_B_M1008_g B
+ N_B_c_80_n B PM_SKY130_FD_SC_HDLL__AND2_4%B
x_PM_SKY130_FD_SC_HDLL__AND2_4%A_27_47# N_A_27_47#_M1002_s N_A_27_47#_M1004_d
+ N_A_27_47#_c_111_n N_A_27_47#_M1001_g N_A_27_47#_c_120_n N_A_27_47#_M1000_g
+ N_A_27_47#_c_112_n N_A_27_47#_M1003_g N_A_27_47#_c_121_n N_A_27_47#_M1005_g
+ N_A_27_47#_c_113_n N_A_27_47#_M1007_g N_A_27_47#_c_122_n N_A_27_47#_M1006_g
+ N_A_27_47#_c_123_n N_A_27_47#_M1011_g N_A_27_47#_c_114_n N_A_27_47#_M1010_g
+ N_A_27_47#_c_115_n N_A_27_47#_c_116_n N_A_27_47#_c_130_n N_A_27_47#_c_131_n
+ N_A_27_47#_c_139_n N_A_27_47#_c_132_n N_A_27_47#_c_117_n N_A_27_47#_c_124_n
+ N_A_27_47#_c_125_n N_A_27_47#_c_118_n N_A_27_47#_c_119_n
+ PM_SKY130_FD_SC_HDLL__AND2_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND2_4%VPWR N_VPWR_M1004_s N_VPWR_M1008_d N_VPWR_M1005_s
+ N_VPWR_M1011_s N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n N_VPWR_c_225_n
+ N_VPWR_c_226_n N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n N_VPWR_c_230_n
+ VPWR N_VPWR_c_231_n N_VPWR_c_221_n N_VPWR_c_233_n N_VPWR_c_234_n
+ PM_SKY130_FD_SC_HDLL__AND2_4%VPWR
x_PM_SKY130_FD_SC_HDLL__AND2_4%X N_X_M1001_s N_X_M1007_s N_X_M1000_d N_X_M1006_d
+ N_X_c_307_n N_X_c_281_n N_X_c_284_n N_X_c_288_n N_X_c_322_p N_X_c_311_n
+ N_X_c_290_n N_X_c_279_n N_X_c_294_n N_X_c_298_n N_X_c_300_n X N_X_c_277_n X
+ PM_SKY130_FD_SC_HDLL__AND2_4%X
x_PM_SKY130_FD_SC_HDLL__AND2_4%VGND N_VGND_M1009_d N_VGND_M1003_d N_VGND_M1010_d
+ N_VGND_c_340_n N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n VGND
+ N_VGND_c_344_n N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n
+ PM_SKY130_FD_SC_HDLL__AND2_4%VGND
cc_1 VNB N_A_c_55_n 0.0333349f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_2 VNB N_A_c_56_n 0.0216244f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_3 VNB N_A_c_57_n 0.0144607f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_4 VNB N_B_c_78_n 0.0174896f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_5 VNB N_B_c_79_n 0.0243152f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_6 VNB N_B_c_80_n 0.0039707f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_7 VNB N_A_27_47#_c_111_n 0.0177885f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_8 VNB N_A_27_47#_c_112_n 0.016944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_113_n 0.0173895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_114_n 0.019214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_115_n 0.00929734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_116_n 0.0141802f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_117_n 0.00132882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_118_n 0.00171227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_119_n 0.0787851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_221_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_X_c_277_n 0.0137701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 0.0250873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_340_n 0.00508483f $X=-0.19 $Y=-0.24 $X2=0.28 $Y2=1.16
cc_20 VNB N_VGND_c_341_n 0.0175594f $X=-0.19 $Y=-0.24 $X2=0.28 $Y2=1.53
cc_21 VNB N_VGND_c_342_n 0.0167346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_343_n 0.0127542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_344_n 0.029709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_345_n 0.0108275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_346_n 0.202584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_347_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_348_n 0.00538815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VPB N_A_c_55_n 0.0327781f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_29 VPB N_A_c_57_n 0.0116013f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_30 VPB N_B_c_79_n 0.0275692f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_31 VPB N_B_c_80_n 0.0036572f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_32 VPB N_A_27_47#_c_120_n 0.0166972f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_33 VPB N_A_27_47#_c_121_n 0.0160009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_47#_c_122_n 0.0162845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_47#_c_123_n 0.0182654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_47#_c_124_n 0.00127583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_c_125_n 0.00920717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_118_n 4.55278e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_119_n 0.0494011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_222_n 0.0103989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_223_n 0.0274522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_224_n 0.0183766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_225_n 0.00449519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_226_n 0.0168506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_227_n 3.32571e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_228_n 0.024116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_229_n 0.0145309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_230_n 0.00583344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_231_n 0.0116899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_221_n 0.0515561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_233_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_234_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_X_c_279_n 0.0190701f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB X 0.0123731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 N_A_c_56_n N_B_c_78_n 0.0383812f $X=0.525 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_56 N_A_c_55_n N_B_c_79_n 0.0619093f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_57 N_A_c_57_n N_B_c_79_n 0.0014365f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_c_55_n N_B_c_80_n 0.00275691f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A_c_57_n N_B_c_80_n 0.0267358f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_c_55_n N_A_27_47#_c_115_n 0.00149931f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_c_57_n N_A_27_47#_c_115_n 0.022552f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_c_56_n N_A_27_47#_c_130_n 0.0143005f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A_c_55_n N_A_27_47#_c_131_n 0.00473012f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A_c_55_n N_A_27_47#_c_132_n 0.00460722f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_c_57_n N_A_27_47#_c_132_n 0.002359f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_c_57_n N_VPWR_M1004_s 0.0034771f $X=0.35 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_67 N_A_c_55_n N_VPWR_c_223_n 0.0128981f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A_c_57_n N_VPWR_c_223_n 0.0154387f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_c_55_n N_VPWR_c_224_n 0.00642146f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_c_55_n N_VPWR_c_221_n 0.0107572f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A_c_56_n N_VGND_c_344_n 0.00422112f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_c_56_n N_VGND_c_346_n 0.00665474f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_73 N_B_c_78_n N_A_27_47#_c_111_n 0.0198481f $X=0.885 $Y=0.995 $X2=0 $Y2=0
cc_74 N_B_c_79_n N_A_27_47#_c_120_n 0.016884f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_75 N_B_c_78_n N_A_27_47#_c_130_n 0.013075f $X=0.885 $Y=0.995 $X2=0 $Y2=0
cc_76 N_B_c_79_n N_A_27_47#_c_130_n 0.00482144f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_77 N_B_c_80_n N_A_27_47#_c_130_n 0.0272969f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B_c_79_n N_A_27_47#_c_139_n 0.0189404f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_79 N_B_c_80_n N_A_27_47#_c_139_n 0.0110616f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B_c_79_n N_A_27_47#_c_132_n 6.3834e-19 $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_81 N_B_c_80_n N_A_27_47#_c_132_n 0.0114768f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B_c_78_n N_A_27_47#_c_117_n 0.00382474f $X=0.885 $Y=0.995 $X2=0 $Y2=0
cc_83 N_B_c_80_n N_A_27_47#_c_117_n 0.00185472f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B_c_79_n N_A_27_47#_c_124_n 0.00501441f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B_c_79_n N_A_27_47#_c_118_n 0.00334719f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B_c_80_n N_A_27_47#_c_118_n 0.0264175f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B_c_79_n N_A_27_47#_c_119_n 0.0151169f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B_c_80_n N_A_27_47#_c_119_n 2.86191e-19 $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B_c_79_n N_VPWR_c_223_n 6.31273e-19 $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B_c_79_n N_VPWR_c_224_n 0.00702461f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B_c_79_n N_VPWR_c_225_n 0.0018504f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_92 N_B_c_79_n N_VPWR_c_221_n 0.0126716f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B_c_78_n N_VGND_c_340_n 0.00627434f $X=0.885 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B_c_78_n N_VGND_c_344_n 0.00422112f $X=0.885 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B_c_78_n N_VGND_c_346_n 0.00615216f $X=0.885 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_139_n N_VPWR_M1008_d 0.00759183f $X=1.25 $Y=1.665 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_124_n N_VPWR_M1008_d 0.00114268f $X=1.355 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_131_n N_VPWR_c_223_n 0.0343774f $X=0.74 $Y=1.96 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_131_n N_VPWR_c_224_n 0.0124822f $X=0.74 $Y=1.96 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_120_n N_VPWR_c_225_n 0.00176848f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_139_n N_VPWR_c_225_n 0.0209938f $X=1.25 $Y=1.665 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_120_n N_VPWR_c_226_n 0.00702461f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_c_121_n N_VPWR_c_226_n 0.00447018f $X=2.015 $Y=1.41 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_120_n N_VPWR_c_227_n 6.3373e-19 $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_121_n N_VPWR_c_227_n 0.0137193f $X=2.015 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_122_n N_VPWR_c_227_n 0.0102323f $X=2.495 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_27_47#_c_123_n N_VPWR_c_227_n 5.80987e-19 $X=2.975 $Y=1.41 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_c_122_n N_VPWR_c_228_n 6.18489e-19 $X=2.495 $Y=1.41 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_c_123_n N_VPWR_c_228_n 0.0146077f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_122_n N_VPWR_c_229_n 0.00642146f $X=2.495 $Y=1.41 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_c_123_n N_VPWR_c_229_n 0.00447018f $X=2.975 $Y=1.41 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_M1004_d N_VPWR_c_221_n 0.00655879f $X=0.59 $Y=1.485 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_120_n N_VPWR_c_221_n 0.0126606f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_121_n N_VPWR_c_221_n 0.00766229f $X=2.015 $Y=1.41 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_c_122_n N_VPWR_c_221_n 0.0107337f $X=2.495 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_123_n N_VPWR_c_221_n 0.00766229f $X=2.975 $Y=1.41 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_c_131_n N_VPWR_c_221_n 0.00684987f $X=0.74 $Y=1.96 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_112_n N_X_c_281_n 0.0115023f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_113_n N_X_c_281_n 0.0114248f $X=2.47 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_119_n N_X_c_281_n 0.00359098f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_121_n N_X_c_284_n 0.0175805f $X=2.015 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_122_n N_X_c_284_n 0.0168709f $X=2.495 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_125_n N_X_c_284_n 0.0480846f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_119_n N_X_c_284_n 0.00161384f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_125_n N_X_c_288_n 0.0156439f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_119_n N_X_c_288_n 0.00136562f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_114_n N_X_c_290_n 0.017501f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_125_n N_X_c_290_n 0.00554628f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_123_n N_X_c_279_n 0.0217949f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_27_47#_c_125_n N_X_c_279_n 0.0056208f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_27_47#_c_130_n N_X_c_294_n 0.0135923f $X=1.25 $Y=0.71 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_117_n N_X_c_294_n 0.0025314f $X=1.355 $Y=1.02 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_125_n N_X_c_294_n 0.0620053f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_27_47#_c_119_n N_X_c_294_n 0.00339319f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_125_n N_X_c_298_n 0.0151856f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_119_n N_X_c_298_n 0.00452326f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_125_n N_X_c_300_n 0.0156439f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_119_n N_X_c_300_n 0.00136936f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_123_n X 0.00433213f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_114_n X 0.01719f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_125_n X 0.015876f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_130_n A_120_47# 0.00271764f $X=1.25 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_143 N_A_27_47#_c_130_n N_VGND_M1009_d 0.0109207f $X=1.25 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_144 N_A_27_47#_c_117_n N_VGND_M1009_d 0.00103313f $X=1.355 $Y=1.02 $X2=-0.19
+ $Y2=-0.24
cc_145 N_A_27_47#_c_111_n N_VGND_c_340_n 0.00320729f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_c_130_n N_VGND_c_340_n 0.0254969f $X=1.25 $Y=0.71 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_111_n N_VGND_c_341_n 0.00558147f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_112_n N_VGND_c_341_n 0.0035176f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_130_n N_VGND_c_341_n 9.77174e-19 $X=1.25 $Y=0.71 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_113_n N_VGND_c_342_n 5.14094e-19 $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_c_114_n N_VGND_c_342_n 0.0102626f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_113_n N_VGND_c_343_n 0.0035176f $X=2.47 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_114_n N_VGND_c_343_n 0.00211056f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_116_n N_VGND_c_344_n 0.021716f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_130_n N_VGND_c_344_n 0.00965588f $X=1.25 $Y=0.71 $X2=0 $Y2=0
cc_156 N_A_27_47#_M1002_s N_VGND_c_346_n 0.00261673f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_111_n N_VGND_c_346_n 0.0104824f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_112_n N_VGND_c_346_n 0.00424616f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_113_n N_VGND_c_346_n 0.00431085f $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_114_n N_VGND_c_346_n 0.0029608f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_116_n N_VGND_c_346_n 0.0125626f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_130_n N_VGND_c_346_n 0.0204516f $X=1.25 $Y=0.71 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_111_n N_VGND_c_348_n 0.00110114f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_112_n N_VGND_c_348_n 0.00856754f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_113_n N_VGND_c_348_n 0.00685368f $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_114_n N_VGND_c_348_n 4.66812e-19 $X=3 $Y=0.995 $X2=0 $Y2=0
cc_167 N_VPWR_c_221_n N_X_M1000_d 0.00621163f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_168 N_VPWR_c_221_n N_X_M1006_d 0.00621163f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_169 N_VPWR_c_226_n N_X_c_307_n 0.0131506f $X=2.04 $Y=2.72 $X2=0 $Y2=0
cc_170 N_VPWR_c_221_n N_X_c_307_n 0.00722976f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_171 N_VPWR_M1005_s N_X_c_284_n 0.00364629f $X=2.105 $Y=1.485 $X2=0 $Y2=0
cc_172 N_VPWR_c_227_n N_X_c_284_n 0.0209288f $X=2.255 $Y=2.02 $X2=0 $Y2=0
cc_173 N_VPWR_c_229_n N_X_c_311_n 0.0131506f $X=3 $Y=2.72 $X2=0 $Y2=0
cc_174 N_VPWR_c_221_n N_X_c_311_n 0.00722976f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_175 N_VPWR_M1011_s N_X_c_279_n 0.0106112f $X=3.065 $Y=1.485 $X2=0 $Y2=0
cc_176 N_VPWR_c_228_n N_X_c_279_n 0.0268973f $X=3.215 $Y=2.02 $X2=0 $Y2=0
cc_177 N_VPWR_M1011_s X 8.15496e-19 $X=3.065 $Y=1.485 $X2=0 $Y2=0
cc_178 N_X_c_281_n N_VGND_M1003_d 0.00421224f $X=2.64 $Y=0.73 $X2=0 $Y2=0
cc_179 N_X_c_290_n N_VGND_M1010_d 0.00825698f $X=3.29 $Y=0.73 $X2=0 $Y2=0
cc_180 N_X_c_277_n N_VGND_M1010_d 0.00163342f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_181 X N_VGND_M1010_d 6.45193e-19 $X=3.43 $Y=0.85 $X2=0 $Y2=0
cc_182 N_X_c_281_n N_VGND_c_341_n 0.00264153f $X=2.64 $Y=0.73 $X2=0 $Y2=0
cc_183 N_X_c_294_n N_VGND_c_341_n 0.00449666f $X=1.87 $Y=0.68 $X2=0 $Y2=0
cc_184 N_X_c_322_p N_VGND_c_342_n 0.0143006f $X=2.735 $Y=0.42 $X2=0 $Y2=0
cc_185 N_X_c_290_n N_VGND_c_342_n 0.0174984f $X=3.29 $Y=0.73 $X2=0 $Y2=0
cc_186 N_X_c_277_n N_VGND_c_342_n 0.0075136f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_187 N_X_c_281_n N_VGND_c_343_n 0.00346656f $X=2.64 $Y=0.73 $X2=0 $Y2=0
cc_188 N_X_c_322_p N_VGND_c_343_n 0.0130838f $X=2.735 $Y=0.42 $X2=0 $Y2=0
cc_189 N_X_c_290_n N_VGND_c_343_n 0.00259276f $X=3.29 $Y=0.73 $X2=0 $Y2=0
cc_190 N_X_c_277_n N_VGND_c_345_n 0.00402329f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_191 N_X_M1001_s N_VGND_c_346_n 0.00648119f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_192 N_X_M1007_s N_VGND_c_346_n 0.00368085f $X=2.545 $Y=0.235 $X2=0 $Y2=0
cc_193 N_X_c_281_n N_VGND_c_346_n 0.0118634f $X=2.64 $Y=0.73 $X2=0 $Y2=0
cc_194 N_X_c_322_p N_VGND_c_346_n 0.00721345f $X=2.735 $Y=0.42 $X2=0 $Y2=0
cc_195 N_X_c_290_n N_VGND_c_346_n 0.00588502f $X=3.29 $Y=0.73 $X2=0 $Y2=0
cc_196 N_X_c_294_n N_VGND_c_346_n 0.00604783f $X=1.87 $Y=0.68 $X2=0 $Y2=0
cc_197 N_X_c_277_n N_VGND_c_346_n 0.00631464f $X=3.43 $Y=0.845 $X2=0 $Y2=0
cc_198 N_X_c_281_n N_VGND_c_348_n 0.0200941f $X=2.64 $Y=0.73 $X2=0 $Y2=0
cc_199 N_X_c_322_p N_VGND_c_348_n 0.0117256f $X=2.735 $Y=0.42 $X2=0 $Y2=0
cc_200 A_120_47# N_VGND_c_346_n 0.00239227f $X=0.6 $Y=0.235 $X2=0.425 $Y2=0.71
