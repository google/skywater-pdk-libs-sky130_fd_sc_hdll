* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__and2_2 A B VGND VNB VPB VPWR X
X0 VGND a_27_75# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A a_27_75# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 a_27_75# A a_123_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 X a_27_75# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_123_75# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_27_75# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 X a_27_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_27_75# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
.ends
