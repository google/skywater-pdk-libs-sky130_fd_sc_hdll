* File: sky130_fd_sc_hdll__sdfxbp_1.spice
* Created: Thu Aug 27 19:27:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdfxbp_1.pex.spice"
.subckt sky130_fd_sc_hdll__sdfxbp_1  VNB VPB CLK SCE D SCD VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* SCD	SCD
* D	D
* SCE	SCE
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_CLK_M1023_g N_A_27_47#_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_211_363#_M1001_d N_A_27_47#_M1001_g N_VGND_M1023_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_SCE_M1017_g N_A_319_47#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.1302 PD=0.86 PS=1.46 NRD=32.856 NRS=7.14 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1025 A_529_47# N_A_319_47#_M1025_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0546 AS=0.0924 PD=0.68 PS=0.86 NRD=21.42 NRS=12.852 M=1 R=2.8 SA=75000.8
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_604_369#_M1010_d N_D_M1010_g A_529_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0546 PD=0.8 PS=0.68 NRD=14.28 NRS=21.42 M=1 R=2.8 SA=75001.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1015 A_717_47# N_SCE_M1015_g N_A_604_369#_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0483 AS=0.0798 PD=0.65 PS=0.8 NRD=17.136 NRS=14.28 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_SCD_M1033_g A_717_47# VNB NSHORT L=0.15 W=0.42 AD=0.1428
+ AS=0.0483 PD=1.52 PS=0.65 NRD=21.42 NRS=17.136 M=1 R=2.8 SA=75002.1 SB=75000.3
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_1001_47#_M1006_d N_A_27_47#_M1006_g N_A_604_369#_M1006_s VNB NSHORT
+ L=0.15 W=0.36 AD=0.0774 AS=0.1008 PD=0.79 PS=1.28 NRD=34.992 NRS=4.992 M=1
+ R=2.4 SA=75000.2 SB=75003.8 A=0.054 P=1.02 MULT=1
MM1029 A_1117_47# N_A_211_363#_M1029_g N_A_1001_47#_M1006_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0634154 AS=0.0774 PD=0.701538 PS=0.79 NRD=40.38 NRS=14.988 M=1
+ R=2.4 SA=75000.8 SB=75003.2 A=0.054 P=1.02 MULT=1
MM1014 N_VGND_M1014_d N_A_1179_183#_M1014_g A_1117_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.139313 AS=0.0739846 PD=1.04604 PS=0.818462 NRD=61.428 NRS=34.608 M=1
+ R=2.8 SA=75001.1 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1003 N_A_1179_183#_M1003_d N_A_1001_47#_M1003_g N_VGND_M1014_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.126592 AS=0.212287 PD=1.2736 PS=1.59396 NRD=4.68 NRS=34.68
+ M=1 R=4.26667 SA=75001.4 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1024 N_A_1464_413#_M1024_d N_A_211_363#_M1024_g N_A_1179_183#_M1003_d VNB
+ NSHORT L=0.15 W=0.36 AD=0.0927 AS=0.071208 PD=0.875 PS=0.7164 NRD=43.332
+ NRS=16.656 M=1 R=2.4 SA=75002.6 SB=75001.4 A=0.054 P=1.02 MULT=1
MM1034 A_1615_47# N_A_27_47#_M1034_g N_A_1464_413#_M1024_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0667385 AS=0.0927 PD=0.715385 PS=0.875 NRD=43.452 NRS=34.992 M=1
+ R=2.4 SA=75003.3 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1020 N_VGND_M1020_d N_A_1653_315#_M1020_g A_1615_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0778615 PD=1.36 PS=0.834615 NRD=0 NRS=37.248 M=1 R=2.8
+ SA=75003.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_1464_413#_M1035_g N_A_1653_315#_M1035_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1032 N_Q_M1032_d N_A_1653_315#_M1032_g N_VGND_M1035_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_1653_315#_M1011_g N_A_2114_47#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0914579 AS=0.1302 PD=0.812523 PS=1.46 NRD=17.856 NRS=12.852
+ M=1 R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1030 N_Q_N_M1030_d N_A_2114_47#_M1030_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.141542 PD=1.82 PS=1.25748 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_CLK_M1007_g N_A_27_47#_M1007_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1028 N_A_211_363#_M1028_d N_A_27_47#_M1028_g N_VPWR_M1007_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1018 N_VPWR_M1018_d N_SCE_M1018_g N_A_319_47#_M1018_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1013 A_503_369# N_SCE_M1013_g N_VPWR_M1018_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.104 AS=0.0928 PD=0.965 PS=0.93 NRD=33.0763 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1016 N_A_604_369#_M1016_d N_D_M1016_g A_503_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.104 PD=0.93 PS=0.965 NRD=1.5366 NRS=33.0763 M=1 R=3.55556
+ SA=90001.2 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1009 A_698_369# N_A_319_47#_M1009_g N_A_604_369#_M1016_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1072 AS=0.0928 PD=0.975 PS=0.93 NRD=34.6129 NRS=1.5366 M=1
+ R=3.55556 SA=90001.6 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1004 N_VPWR_M1004_d N_SCD_M1004_g A_698_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1888 AS=0.1072 PD=1.87 PS=0.975 NRD=9.2196 NRS=34.6129 M=1 R=3.55556
+ SA=90002.1 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1022 N_A_1001_47#_M1022_d N_A_211_363#_M1022_g N_A_604_369#_M1022_s VPB
+ PHIGHVT L=0.18 W=0.42 AD=0.07035 AS=0.1134 PD=0.755 PS=1.38 NRD=14.0658
+ NRS=2.3443 M=1 R=2.33333 SA=90000.2 SB=90003.7 A=0.0756 P=1.2 MULT=1
MM1019 A_1111_413# N_A_27_47#_M1019_g N_A_1001_47#_M1022_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0735 AS=0.07035 PD=0.77 PS=0.755 NRD=56.2829 NRS=11.7215 M=1
+ R=2.33333 SA=90000.7 SB=90003.2 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A_1179_183#_M1000_g A_1111_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.132623 AS=0.0735 PD=0.918974 PS=0.77 NRD=116.072 NRS=56.2829 M=1
+ R=2.33333 SA=90001.2 SB=90002.7 A=0.0756 P=1.2 MULT=1
MM1021 N_A_1179_183#_M1021_d N_A_1001_47#_M1021_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.18 W=0.75 AD=0.147885 AS=0.236827 PD=1.40385 PS=1.64103 NRD=1.3002
+ NRS=1.3002 M=1 R=4.16667 SA=90001.2 SB=90001.2 A=0.135 P=1.86 MULT=1
MM1005 N_A_1464_413#_M1005_d N_A_27_47#_M1005_g N_A_1179_183#_M1021_d VPB
+ PHIGHVT L=0.18 W=0.42 AD=0.0609 AS=0.0828154 PD=0.71 PS=0.786154 NRD=2.3443
+ NRS=28.1316 M=1 R=2.33333 SA=90002.5 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1031 A_1558_413# N_A_211_363#_M1031_g N_A_1464_413#_M1005_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.10185 AS=0.0609 PD=0.905 PS=0.71 NRD=87.9408 NRS=2.3443 M=1
+ R=2.33333 SA=90002.9 SB=90001 A=0.0756 P=1.2 MULT=1
MM1026 N_VPWR_M1026_d N_A_1653_315#_M1026_g A_1558_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1617 AS=0.10185 PD=1.61 PS=0.905 NRD=53.9386 NRS=87.9408 M=1
+ R=2.33333 SA=90003.6 SB=90000.3 A=0.0756 P=1.2 MULT=1
MM1012 N_VPWR_M1012_d N_A_1464_413#_M1012_g N_A_1653_315#_M1012_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1002 N_Q_M1002_d N_A_1653_315#_M1002_g N_VPWR_M1012_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_1653_315#_M1008_g N_A_2114_47#_M1008_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.126595 AS=0.1728 PD=1.05756 PS=1.82 NRD=21.5321 NRS=1.5366
+ M=1 R=3.55556 SA=90000.2 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1027 N_Q_N_M1027_d N_A_2114_47#_M1027_g N_VPWR_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.197805 PD=2.54 PS=1.65244 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX36_noxref VNB VPB NWDIODE A=19.8057 P=27.89
c_115 VNB 0 1.8505e-19 $X=0.145 $Y=-0.085
c_225 VPB 0 1.48877e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__sdfxbp_1.pxi.spice"
*
.ends
*
*
