* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 VPWR A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_503_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_1375_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VPWR A1 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_1375_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND A2 a_1375_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_297# B1 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_511_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_503_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y B1 a_503_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_511_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_1375_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_27_297# B2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_511_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND A2 a_1375_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y A1 a_1375_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VPWR A1 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 Y A1 a_1375_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VGND B2 a_503_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_511_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 VGND B2 a_503_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_503_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 Y B1 a_503_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_503_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_27_297# B2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 a_511_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 a_511_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 a_511_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 a_1375_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 a_27_297# B1 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 a_511_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
