* File: sky130_fd_sc_hdll__o21ba_1.spice
* Created: Thu Aug 27 19:19:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21ba_1.pex.spice"
.subckt sky130_fd_sc_hdll__o21ba_1  VNB VPB B1_N A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_79_199#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121799 AS=0.169 PD=1.19673 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1002 N_A_222_93#_M1002_d N_B1_N_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1302 AS=0.0787009 PD=1.46 PS=0.773271 NRD=12.852 NRS=17.136 M=1
+ R=2.8 SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_460_47#_M1009_d N_A_222_93#_M1009_g N_A_79_199#_M1009_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.10725 AS=0.195 PD=0.98 PS=1.9 NRD=0.912 NRS=6.456 M=1
+ R=4.33333 SA=75000.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_460_47#_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1003 N_A_460_47#_M1003_d N_A1_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2145 AS=0.08775 PD=1.96 PS=0.92 NRD=11.076 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_79_199#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.236408 AS=0.27 PD=1.9507 PS=2.54 NRD=6.8753 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.4 A=0.18 P=2.36 MULT=1
MM1001 N_A_222_93#_M1001_d N_B1_N_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1218 AS=0.0992915 PD=1.42 PS=0.819296 NRD=2.3443 NRS=85.0843 M=1
+ R=2.33333 SA=90000.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1000 N_A_79_199#_M1000_d N_A_222_93#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18
+ W=1 AD=0.15 AS=0.3 PD=1.3 PS=2.6 NRD=2.9353 NRS=6.8753 M=1 R=5.55556
+ SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1008 A_554_297# N_A2_M1008_g N_A_79_199#_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.15 PD=1.29 PS=1.3 NRD=17.7103 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g A_554_297# VPB PHIGHVT L=0.18 W=1 AD=0.29
+ AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=17.7103 M=1 R=5.55556 SA=90001.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_13 A2 A2 PROBETYPE=1
pX12_noxref noxref_14 A1 A1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o21ba_1.pxi.spice"
*
.ends
*
*
