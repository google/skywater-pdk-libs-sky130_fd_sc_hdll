* File: sky130_fd_sc_hdll__ebufn_2.pex.spice
* Created: Wed Sep  2 08:30:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EBUFN_2%A 3 6 7 9 10 11 15
c36 6 0 1.77992e-20 $X=0.495 $Y=1.67
c37 3 0 8.80328e-20 $X=0.47 $Y=0.445
r38 15 18 37.7065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.16
+ $X2=0.565 $Y2=1.325
r39 15 17 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.16
+ $X2=0.565 $Y2=0.995
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r41 11 16 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.645 $Y=1.53
+ $X2=0.645 $Y2=1.16
r42 10 16 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=0.645 $Y=0.85
+ $X2=0.645 $Y2=1.16
r43 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r44 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.67 $X2=0.495
+ $Y2=1.77
r45 6 18 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.495 $Y=1.67
+ $X2=0.495 $Y2=1.325
r46 3 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_2%TE_B 3 6 7 9 10 12 14 15 17 19 20 21 24
r69 27 28 22.0037 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.135 $Y=1.395
+ $X2=1.135 $Y2=1.47
r70 24 27 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.135 $Y=1.16
+ $X2=1.135 $Y2=1.395
r71 24 26 42.7143 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.135 $Y=1.16
+ $X2=1.135 $Y2=1.015
r72 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.135
+ $Y=1.16 $X2=1.135 $Y2=1.16
r73 21 25 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=1.122 $Y=0.85
+ $X2=1.122 $Y2=1.16
r74 17 19 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.53 $Y=1.47
+ $X2=2.53 $Y2=2.015
r75 16 20 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.15 $Y=1.395 $X2=2.06
+ $Y2=1.395
r76 15 17 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.44 $Y=1.395
+ $X2=2.53 $Y2=1.47
r77 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.44 $Y=1.395
+ $X2=2.15 $Y2=1.395
r78 12 20 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.06 $Y=1.47 $X2=2.06
+ $Y2=1.395
r79 12 14 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.06 $Y=1.47
+ $X2=2.06 $Y2=2.015
r80 11 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.3 $Y=1.395
+ $X2=1.135 $Y2=1.395
r81 10 20 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.97 $Y=1.395 $X2=2.06
+ $Y2=1.395
r82 10 11 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.97 $Y=1.395
+ $X2=1.3 $Y2=1.395
r83 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.07 $Y=1.77 $X2=1.07
+ $Y2=2.165
r84 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.07 $Y=1.67 $X2=1.07
+ $Y2=1.77
r85 6 28 66.3154 $w=2e-07 $l=2e-07 $layer=POLY_cond $X=1.07 $Y=1.67 $X2=1.07
+ $Y2=1.47
r86 3 26 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.045 $Y=0.445
+ $X2=1.045 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_2%A_224_47# 1 2 7 9 10 11 14 15 21 24 26 29
+ 34 36 38
c81 38 0 1.36116e-19 $X=2.987 $Y=0.96
c82 34 0 1.77992e-20 $X=1.682 $Y=1.605
c83 15 0 8.80328e-20 $X=1.55 $Y=0.425
c84 11 0 1.57352e-19 $X=2.57 $Y=1.035
r85 32 34 11.4164 $w=3.18e-07 $l=3.17e-07 $layer=LI1_cond $X=1.365 $Y=1.605
+ $X2=1.682 $Y2=1.605
r86 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3 $Y=1.16
+ $X2=3 $Y2=1.16
r87 27 36 1.65465 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=1.83 $Y=1.15 $X2=1.69
+ $Y2=1.15
r88 27 29 53.9343 $w=2.48e-07 $l=1.17e-06 $layer=LI1_cond $X=1.83 $Y=1.15 $X2=3
+ $Y2=1.15
r89 26 34 1.86265 $w=2.65e-07 $l=1.6e-07 $layer=LI1_cond $X=1.682 $Y=1.445
+ $X2=1.682 $Y2=1.605
r90 25 36 4.80568 $w=2.72e-07 $l=1.28938e-07 $layer=LI1_cond $X=1.682 $Y=1.275
+ $X2=1.69 $Y2=1.15
r91 25 26 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=1.682 $Y=1.275
+ $X2=1.682 $Y2=1.445
r92 24 36 4.80568 $w=2.72e-07 $l=1.25e-07 $layer=LI1_cond $X=1.69 $Y=1.025
+ $X2=1.69 $Y2=1.15
r93 23 24 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=1.69 $Y=0.595
+ $X2=1.69 $Y2=1.025
r94 19 32 1.30983 $w=2.9e-07 $l=1.6e-07 $layer=LI1_cond $X=1.365 $Y=1.765
+ $X2=1.365 $Y2=1.605
r95 19 21 18.0814 $w=2.88e-07 $l=4.55e-07 $layer=LI1_cond $X=1.365 $Y=1.765
+ $X2=1.365 $Y2=2.22
r96 15 23 6.89985 $w=3.4e-07 $l=2.29565e-07 $layer=LI1_cond $X=1.55 $Y=0.425
+ $X2=1.69 $Y2=0.595
r97 15 17 8.30437 $w=3.38e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.425
+ $X2=1.305 $Y2=0.425
r98 14 38 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.915 $Y=0.56
+ $X2=2.915 $Y2=0.96
r99 10 30 25.4182 $w=2.95e-07 $l=1.25e-07 $layer=POLY_cond $X=2.987 $Y=1.035
+ $X2=2.987 $Y2=1.16
r100 10 38 29.7108 $w=2.95e-07 $l=7.5e-08 $layer=POLY_cond $X=2.987 $Y=1.035
+ $X2=2.987 $Y2=0.96
r101 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.84 $Y=1.035
+ $X2=2.57 $Y2=1.035
r102 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.495 $Y=0.96
+ $X2=2.57 $Y2=1.035
r103 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.495 $Y=0.96 $X2=2.495
+ $Y2=0.56
r104 2 21 600 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.845 $X2=1.305 $Y2=2.22
r105 1 17 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.235 $X2=1.305 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_2%A_27_47# 1 2 9 11 13 14 16 19 27 29 30 31
+ 38 41
c77 31 0 1.40706e-19 $X=3.57 $Y=1.145
c78 14 0 2.46566e-20 $X=3.995 $Y=1.41
c79 11 0 1.98649e-20 $X=3.525 $Y=1.41
r80 38 39 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=3.995 $Y=1.217
+ $X2=4.02 $Y2=1.217
r81 36 38 33.5118 $w=3.38e-07 $l=2.35e-07 $layer=POLY_cond $X=3.76 $Y=1.217
+ $X2=3.995 $Y2=1.217
r82 34 36 33.5118 $w=3.38e-07 $l=2.35e-07 $layer=POLY_cond $X=3.525 $Y=1.217
+ $X2=3.76 $Y2=1.217
r83 33 34 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=3.5 $Y=1.217
+ $X2=3.525 $Y2=1.217
r84 30 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.16 $X2=3.76 $Y2=1.16
r85 29 31 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=3.765 $Y=1.145
+ $X2=3.57 $Y2=1.145
r86 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.765 $Y=1.145
+ $X2=3.765 $Y2=1.145
r87 27 31 3.94801 $w=1.4e-07 $l=3.19e-06 $layer=MET1_cond $X=0.38 $Y=1.19
+ $X2=3.57 $Y2=1.19
r88 25 45 47.6491 $w=2.58e-07 $l=1.075e-06 $layer=LI1_cond $X=0.215 $Y=1.145
+ $X2=0.215 $Y2=2.22
r89 25 41 31.0273 $w=2.58e-07 $l=7e-07 $layer=LI1_cond $X=0.215 $Y=1.145
+ $X2=0.215 $Y2=0.445
r90 24 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.235 $Y=1.145
+ $X2=0.38 $Y2=1.145
r91 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.235 $Y=1.145
+ $X2=0.235 $Y2=1.145
r92 17 39 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.02 $Y=1.025
+ $X2=4.02 $Y2=1.217
r93 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.02 $Y=1.025
+ $X2=4.02 $Y2=0.56
r94 14 38 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.995 $Y=1.41
+ $X2=3.995 $Y2=1.217
r95 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.995 $Y=1.41
+ $X2=3.995 $Y2=1.985
r96 11 34 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.525 $Y=1.41
+ $X2=3.525 $Y2=1.217
r97 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.525 $Y=1.41
+ $X2=3.525 $Y2=1.985
r98 7 33 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.5 $Y=1.025 $X2=3.5
+ $Y2=1.217
r99 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.5 $Y=1.025 $X2=3.5
+ $Y2=0.56
r100 2 45 600 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.22
r101 1 41 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_2%VPWR 1 2 9 12 15 18 20 36 37 40
r54 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r56 34 37 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.37 $Y2=2.72
r57 33 36 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=4.37 $Y2=2.72
r58 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 31 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r60 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 28 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 27 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r64 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 25 40 11.0851 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=1 $Y=2.72 $X2=0.757
+ $Y2=2.72
r66 25 27 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1 $Y=2.72 $X2=1.15
+ $Y2=2.72
r67 20 40 11.0851 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.757 $Y2=2.72
r68 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 18 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 16 33 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.46 $Y=2.72 $X2=2.53
+ $Y2=2.72
r72 15 30 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.08 $Y=2.72 $X2=2.07
+ $Y2=2.72
r73 14 16 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.27 $Y=2.72 $X2=2.46
+ $Y2=2.72
r74 14 15 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.27 $Y=2.72 $X2=2.08
+ $Y2=2.72
r75 12 14 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.27 $Y=2.36
+ $X2=2.27 $Y2=2.72
r76 7 40 1.99554 $w=4.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.757 $Y=2.635
+ $X2=0.757 $Y2=2.72
r77 7 9 15.1668 $w=4.83e-07 $l=6.15e-07 $layer=LI1_cond $X=0.757 $Y=2.635
+ $X2=0.757 $Y2=2.02
r78 2 12 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.15
+ $Y=1.545 $X2=2.295 $Y2=2.36
r79 1 9 300 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.845 $X2=0.785 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_2%A_340_309# 1 2 3 12 15 16 20 24 25
r46 23 25 9.59153 $w=5.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.215 $Y=2.2
+ $X2=3.375 $Y2=2.2
r47 23 24 18.0543 $w=5.28e-07 $l=5.35e-07 $layer=LI1_cond $X=3.215 $Y=2.2
+ $X2=2.68 $Y2=2.2
r48 18 20 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=4.295 $Y=2.295
+ $X2=4.295 $Y2=1.96
r49 16 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.165 $Y=2.38
+ $X2=4.295 $Y2=2.295
r50 16 25 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.165 $Y=2.38
+ $X2=3.375 $Y2=2.38
r51 15 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.91 $Y=2.02
+ $X2=2.68 $Y2=2.02
r52 10 15 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.805 $Y=2.105
+ $X2=1.91 $Y2=2.02
r53 10 12 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=1.805 $Y=2.105
+ $X2=1.805 $Y2=2.3
r54 3 20 300 $w=1.7e-07 $l=5.51362e-07 $layer=licon1_PDIFF $count=2 $X=4.085
+ $Y=1.485 $X2=4.25 $Y2=1.96
r55 2 23 300 $w=1.7e-07 $l=1.00958e-06 $layer=licon1_PDIFF $count=2 $X=2.62
+ $Y=1.545 $X2=3.215 $Y2=2.3
r56 1 12 600 $w=1.7e-07 $l=8.15107e-07 $layer=licon1_PDIFF $count=1 $X=1.7
+ $Y=1.545 $X2=1.825 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_2%Z 1 2 7 11 13 14 15 16 17 18 19 29 31 36
+ 40 43 49
c58 29 0 1.82009e-19 $X=3.595 $Y=1.605
c59 11 0 1.98649e-20 $X=4.23 $Y=1.535
c60 7 0 2.76821e-19 $X=4.23 $Y=0.745
r61 51 53 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=3.795 $Y=1.605
+ $X2=3.795 $Y2=1.655
r62 49 51 2.01678 $w=3.98e-07 $l=7e-08 $layer=LI1_cond $X=3.795 $Y=1.535
+ $X2=3.795 $Y2=1.605
r63 29 51 2.04652 $w=3.2e-07 $l=2e-07 $layer=LI1_cond $X=3.595 $Y=1.605
+ $X2=3.795 $Y2=1.605
r64 18 19 9.41096 $w=3.98e-07 $l=2.55e-07 $layer=LI1_cond $X=4.345 $Y=1.19
+ $X2=4.345 $Y2=1.445
r65 17 43 3.33465 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.345 $Y=0.745
+ $X2=4.345 $Y2=0.855
r66 17 18 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.345 $Y=0.895
+ $X2=4.345 $Y2=1.19
r67 17 43 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=4.345 $Y=0.895
+ $X2=4.345 $Y2=0.855
r68 16 53 6.19438 $w=3.98e-07 $l=2.15e-07 $layer=LI1_cond $X=3.795 $Y=1.87
+ $X2=3.795 $Y2=1.655
r69 15 29 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=3.255 $Y=1.605
+ $X2=3.595 $Y2=1.605
r70 15 40 9.00346 $w=3.18e-07 $l=2.5e-07 $layer=LI1_cond $X=3.255 $Y=1.605
+ $X2=3.005 $Y2=1.605
r71 14 40 9.29157 $w=3.18e-07 $l=2.58e-07 $layer=LI1_cond $X=2.747 $Y=1.605
+ $X2=3.005 $Y2=1.605
r72 14 36 7.2748 $w=3.18e-07 $l=2.02e-07 $layer=LI1_cond $X=2.747 $Y=1.605
+ $X2=2.545 $Y2=1.605
r73 13 36 10.8042 $w=3.18e-07 $l=3e-07 $layer=LI1_cond $X=2.245 $Y=1.605
+ $X2=2.545 $Y2=1.605
r74 13 31 5.40208 $w=3.18e-07 $l=1.5e-07 $layer=LI1_cond $X=2.245 $Y=1.605
+ $X2=2.095 $Y2=1.605
r75 12 49 5.43236 $w=1.8e-07 $l=2e-07 $layer=LI1_cond $X=3.995 $Y=1.535
+ $X2=3.795 $Y2=1.535
r76 11 19 3.89832 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=4.23 $Y=1.535
+ $X2=4.345 $Y2=1.535
r77 11 12 14.4798 $w=1.78e-07 $l=2.35e-07 $layer=LI1_cond $X=4.23 $Y=1.535
+ $X2=3.995 $Y2=1.535
r78 7 17 3.48622 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=4.23 $Y=0.745
+ $X2=4.345 $Y2=0.745
r79 7 9 24.6204 $w=2.18e-07 $l=4.7e-07 $layer=LI1_cond $X=4.23 $Y=0.745 $X2=3.76
+ $Y2=0.745
r80 2 53 300 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=2 $X=3.615
+ $Y=1.485 $X2=3.76 $Y2=1.655
r81 1 9 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=3.575
+ $Y=0.235 $X2=3.76 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r57 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r58 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r59 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r60 30 33 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=4.37
+ $Y2=0
r61 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r62 29 32 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=4.37
+ $Y2=0
r63 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r64 27 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.68
+ $Y2=0
r65 27 29 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.99
+ $Y2=0
r66 26 40 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r67 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r68 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r69 23 36 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=0.707
+ $Y2=0
r70 23 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=1.15
+ $Y2=0
r71 22 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.49 $Y=0 $X2=2.68
+ $Y2=0
r72 22 25 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=2.49 $Y=0 $X2=1.15
+ $Y2=0
r73 17 36 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.707
+ $Y2=0
r74 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r75 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r76 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r77 11 39 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=0.085
+ $X2=2.68 $Y2=0
r78 11 13 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=2.68 $Y=0.085
+ $X2=2.68 $Y2=0.36
r79 7 36 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0
r80 7 9 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0.36
r81 2 13 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.235 $X2=2.705 $Y2=0.36
r82 1 9 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_2%A_412_47# 1 2 3 10 13 14 18 19 21
r43 19 21 49.9091 $w=1.88e-07 $l=8.55e-07 $layer=LI1_cond $X=3.375 $Y=0.37
+ $X2=4.23 $Y2=0.37
r44 16 18 3.84148 $w=2.83e-07 $l=9.5e-08 $layer=LI1_cond $X=3.232 $Y=0.655
+ $X2=3.232 $Y2=0.56
r45 15 19 7.17723 $w=1.9e-07 $l=1.84483e-07 $layer=LI1_cond $X=3.232 $Y=0.465
+ $X2=3.375 $Y2=0.37
r46 15 18 3.84148 $w=2.83e-07 $l=9.5e-08 $layer=LI1_cond $X=3.232 $Y=0.465
+ $X2=3.232 $Y2=0.56
r47 13 16 7.09239 $w=2e-07 $l=1.85375e-07 $layer=LI1_cond $X=3.09 $Y=0.755
+ $X2=3.232 $Y2=0.655
r48 13 14 42.7 $w=1.98e-07 $l=7.7e-07 $layer=LI1_cond $X=3.09 $Y=0.755 $X2=2.32
+ $Y2=0.755
r49 10 14 7.29955 $w=2e-07 $l=2.03961e-07 $layer=LI1_cond $X=2.16 $Y=0.655
+ $X2=2.32 $Y2=0.755
r50 10 12 3.62188 $w=3.2e-07 $l=9.5e-08 $layer=LI1_cond $X=2.16 $Y=0.655
+ $X2=2.16 $Y2=0.56
r51 3 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.235 $X2=4.23 $Y2=0.38
r52 2 18 182 $w=1.7e-07 $l=4.28515e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.235 $X2=3.23 $Y2=0.56
r53 1 12 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.235 $X2=2.185 $Y2=0.56
.ends

