* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xnor2_2 A B VGND VNB VPB VPWR Y
X0 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_514_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 VGND A a_600_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A a_514_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Y a_27_297# a_600_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 Y B a_514_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VGND B a_600_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_514_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_600_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_600_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_600_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
