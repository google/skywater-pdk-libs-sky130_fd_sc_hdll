* File: sky130_fd_sc_hdll__or3b_4.pxi.spice
* Created: Thu Aug 27 19:24:40 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR3B_4%C_N N_C_N_c_77_n N_C_N_c_78_n N_C_N_M1009_g
+ N_C_N_M1010_g C_N C_N N_C_N_c_76_n PM_SKY130_FD_SC_HDLL__OR3B_4%C_N
x_PM_SKY130_FD_SC_HDLL__OR3B_4%A_186_21# N_A_186_21#_M1002_d N_A_186_21#_M1003_d
+ N_A_186_21#_M1005_d N_A_186_21#_c_106_n N_A_186_21#_M1001_g
+ N_A_186_21#_c_115_n N_A_186_21#_M1000_g N_A_186_21#_c_107_n
+ N_A_186_21#_M1008_g N_A_186_21#_c_116_n N_A_186_21#_M1004_g
+ N_A_186_21#_c_108_n N_A_186_21#_M1012_g N_A_186_21#_c_117_n
+ N_A_186_21#_M1007_g N_A_186_21#_c_118_n N_A_186_21#_M1011_g
+ N_A_186_21#_c_109_n N_A_186_21#_M1013_g N_A_186_21#_c_110_n
+ N_A_186_21#_c_111_n N_A_186_21#_c_112_n N_A_186_21#_c_193_p
+ N_A_186_21#_c_119_n N_A_186_21#_c_113_n N_A_186_21#_c_114_n
+ PM_SKY130_FD_SC_HDLL__OR3B_4%A_186_21#
x_PM_SKY130_FD_SC_HDLL__OR3B_4%A N_A_c_233_n N_A_M1015_g N_A_c_234_n N_A_M1002_g
+ A N_A_c_235_n PM_SKY130_FD_SC_HDLL__OR3B_4%A
x_PM_SKY130_FD_SC_HDLL__OR3B_4%B N_B_c_268_n N_B_M1006_g N_B_c_269_n N_B_M1014_g
+ B B PM_SKY130_FD_SC_HDLL__OR3B_4%B
x_PM_SKY130_FD_SC_HDLL__OR3B_4%A_27_47# N_A_27_47#_M1010_s N_A_27_47#_M1009_s
+ N_A_27_47#_c_296_n N_A_27_47#_M1003_g N_A_27_47#_c_297_n N_A_27_47#_M1005_g
+ N_A_27_47#_c_298_n N_A_27_47#_c_299_n N_A_27_47#_c_300_n N_A_27_47#_c_313_n
+ N_A_27_47#_c_301_n N_A_27_47#_c_329_n N_A_27_47#_c_302_n N_A_27_47#_c_306_n
+ N_A_27_47#_c_338_n PM_SKY130_FD_SC_HDLL__OR3B_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__OR3B_4%VPWR N_VPWR_M1009_d N_VPWR_M1004_d N_VPWR_M1011_d
+ N_VPWR_c_389_n N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n VPWR
+ N_VPWR_c_393_n N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_388_n N_VPWR_c_397_n
+ N_VPWR_c_398_n N_VPWR_c_399_n PM_SKY130_FD_SC_HDLL__OR3B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__OR3B_4%X N_X_M1001_d N_X_M1012_d N_X_M1000_s N_X_M1007_s
+ N_X_c_458_n N_X_c_453_n N_X_c_454_n N_X_c_474_n N_X_c_455_n X X
+ PM_SKY130_FD_SC_HDLL__OR3B_4%X
x_PM_SKY130_FD_SC_HDLL__OR3B_4%VGND N_VGND_M1010_d N_VGND_M1008_s N_VGND_M1013_s
+ N_VGND_M1006_d N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n
+ N_VGND_c_522_n N_VGND_c_523_n N_VGND_c_524_n VGND N_VGND_c_525_n
+ N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n VGND
+ PM_SKY130_FD_SC_HDLL__OR3B_4%VGND
cc_1 VNB N_C_N_M1010_g 0.0359316f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB C_N 0.00882738f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_76_n 0.0413107f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_186_21#_c_106_n 0.0167755f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_186_21#_c_107_n 0.016731f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_6 VNB N_A_186_21#_c_108_n 0.0171691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_186_21#_c_109_n 0.0164255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_186_21#_c_110_n 0.00230632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_186_21#_c_111_n 0.0015978f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_186_21#_c_112_n 0.0106041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_186_21#_c_113_n 0.023569f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_186_21#_c_114_n 0.0763617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_c_233_n 0.0234537f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_14 VNB N_A_c_234_n 0.0169216f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.01
cc_15 VNB N_A_c_235_n 0.00352598f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_16 VNB N_B_c_268_n 0.0171732f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_17 VNB N_B_c_269_n 0.0255339f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.01
cc_18 VNB B 0.00130608f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_19 VNB N_A_27_47#_c_296_n 0.0204077f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_20 VNB N_A_27_47#_c_297_n 0.0273677f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_21 VNB N_A_27_47#_c_298_n 0.0183993f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_22 VNB N_A_27_47#_c_299_n 0.00499741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_300_n 0.00960394f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_24 VNB N_A_27_47#_c_301_n 0.00705029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_302_n 6.47944e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_388_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_453_n 8.7812e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_28 VNB N_X_c_454_n 0.00422882f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_29 VNB N_X_c_455_n 0.00144782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_518_n 0.00470301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_519_n 0.00417622f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_32 VNB N_VGND_c_520_n 0.0161971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_521_n 0.00207171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_522_n 0.0143491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_523_n 0.0211938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_524_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_525_n 0.0226796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_526_n 0.242111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_527_n 0.0232484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_528_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_529_n 0.00649335f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VPB N_C_N_c_77_n 0.0211463f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.625
cc_43 VPB N_C_N_c_78_n 0.0324447f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.725
cc_44 VPB C_N 0.0160532f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_45 VPB N_C_N_c_76_n 0.0101485f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_46 VPB N_A_186_21#_c_115_n 0.0178743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_186_21#_c_116_n 0.0151004f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_48 VPB N_A_186_21#_c_117_n 0.0153796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_186_21#_c_118_n 0.0156001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_186_21#_c_119_n 0.0114264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_186_21#_c_113_n 0.0392722f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_186_21#_c_114_n 0.045425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_c_233_n 0.0248391f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_54 VPB N_A_c_235_n 0.00277287f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_55 VPB N_B_c_269_n 0.0267565f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.01
cc_56 VPB B 0.00120057f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_57 VPB N_A_27_47#_c_297_n 0.0340228f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_58 VPB N_A_27_47#_c_301_n 0.00589909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_302_n 0.00160095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_306_n 0.0187914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_389_n 0.00986749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_390_n 3.18768e-19 $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_63 VPB N_VPWR_c_391_n 0.0132576f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_64 VPB N_VPWR_c_392_n 4.03857e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_393_n 0.0186913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_394_n 0.0133964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_395_n 0.047693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_388_n 0.0523854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_397_n 0.00571014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_398_n 0.00502934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_399_n 0.00516238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_X_c_453_n 8.38654e-19 $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_73 VPB X 0.00445537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 N_C_N_M1010_g N_A_186_21#_c_106_n 0.0155923f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_75 N_C_N_c_77_n N_A_186_21#_c_115_n 0.00844727f $X=0.495 $Y=1.625 $X2=0 $Y2=0
cc_76 N_C_N_c_78_n N_A_186_21#_c_115_n 0.015879f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_77 N_C_N_c_76_n N_A_186_21#_c_114_n 0.0155923f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_78 N_C_N_M1010_g N_A_27_47#_c_298_n 0.00442001f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_79 N_C_N_M1010_g N_A_27_47#_c_299_n 0.0180861f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_80 C_N N_A_27_47#_c_299_n 0.00618246f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_81 N_C_N_c_76_n N_A_27_47#_c_299_n 0.00301897f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_82 C_N N_A_27_47#_c_300_n 0.0227094f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_83 N_C_N_c_76_n N_A_27_47#_c_300_n 0.00599978f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_84 N_C_N_c_78_n N_A_27_47#_c_313_n 0.0183148f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_85 C_N N_A_27_47#_c_313_n 0.00421277f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_86 N_C_N_c_78_n N_A_27_47#_c_301_n 0.00209021f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_87 N_C_N_M1010_g N_A_27_47#_c_301_n 0.0117652f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_88 C_N N_A_27_47#_c_301_n 0.0350078f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_89 N_C_N_c_78_n N_A_27_47#_c_306_n 0.00472318f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_90 C_N N_A_27_47#_c_306_n 0.0226231f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_91 N_C_N_c_76_n N_A_27_47#_c_306_n 8.96314e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_92 N_C_N_c_78_n N_VPWR_c_389_n 0.00396865f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_93 N_C_N_c_78_n N_VPWR_c_393_n 0.00453698f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_94 N_C_N_c_78_n N_VPWR_c_388_n 0.00602858f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_95 N_C_N_M1010_g N_X_c_458_n 5.80679e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_96 N_C_N_M1010_g N_VGND_c_518_n 0.00496578f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_97 N_C_N_M1010_g N_VGND_c_526_n 0.00723476f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_98 N_C_N_M1010_g N_VGND_c_527_n 0.00439206f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_186_21#_c_118_n N_A_c_233_n 0.0361781f $X=2.44 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_100 N_A_186_21#_c_110_n N_A_c_233_n 0.00115955f $X=2.445 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_101 N_A_186_21#_c_111_n N_A_c_233_n 4.63303e-19 $X=2.53 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_102 N_A_186_21#_c_112_n N_A_c_233_n 0.00250198f $X=4.25 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_186_21#_c_114_n N_A_c_233_n 0.0251002f $X=2.44 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_104 N_A_186_21#_c_109_n N_A_c_234_n 0.0200143f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_186_21#_c_111_n N_A_c_234_n 0.00325439f $X=2.53 $Y=1.075 $X2=0 $Y2=0
cc_106 N_A_186_21#_c_112_n N_A_c_234_n 0.0100712f $X=4.25 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_186_21#_c_118_n N_A_c_235_n 0.00125594f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A_186_21#_c_110_n N_A_c_235_n 0.0133948f $X=2.445 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_186_21#_c_111_n N_A_c_235_n 0.00557906f $X=2.53 $Y=1.075 $X2=0 $Y2=0
cc_110 N_A_186_21#_c_112_n N_A_c_235_n 0.0199018f $X=4.25 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_186_21#_c_114_n N_A_c_235_n 0.00258036f $X=2.44 $Y=1.202 $X2=0 $Y2=0
cc_112 N_A_186_21#_c_112_n N_B_c_268_n 0.0115681f $X=4.25 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_113 N_A_186_21#_c_112_n N_B_c_269_n 0.00201602f $X=4.25 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_186_21#_c_119_n N_B_c_269_n 0.0011699f $X=4.25 $Y=2.317 $X2=0 $Y2=0
cc_115 N_A_186_21#_c_112_n B 0.0164428f $X=4.25 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_186_21#_c_112_n N_A_27_47#_c_296_n 0.0115968f $X=4.25 $Y=0.74 $X2=0
+ $Y2=0
cc_117 N_A_186_21#_c_113_n N_A_27_47#_c_296_n 0.00431115f $X=4.352 $Y=2.21 $X2=0
+ $Y2=0
cc_118 N_A_186_21#_c_112_n N_A_27_47#_c_297_n 0.00415219f $X=4.25 $Y=0.74 $X2=0
+ $Y2=0
cc_119 N_A_186_21#_c_119_n N_A_27_47#_c_297_n 0.00926795f $X=4.25 $Y=2.317 $X2=0
+ $Y2=0
cc_120 N_A_186_21#_c_113_n N_A_27_47#_c_297_n 0.016414f $X=4.352 $Y=2.21 $X2=0
+ $Y2=0
cc_121 N_A_186_21#_c_106_n N_A_27_47#_c_299_n 0.00139637f $X=1.005 $Y=0.995
+ $X2=0 $Y2=0
cc_122 N_A_186_21#_c_106_n N_A_27_47#_c_301_n 0.00424215f $X=1.005 $Y=0.995
+ $X2=0 $Y2=0
cc_123 N_A_186_21#_c_115_n N_A_27_47#_c_301_n 0.00460406f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_124 N_A_186_21#_c_115_n N_A_27_47#_c_329_n 0.0159914f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_125 N_A_186_21#_c_116_n N_A_27_47#_c_329_n 0.0130372f $X=1.5 $Y=1.41 $X2=0
+ $Y2=0
cc_126 N_A_186_21#_c_117_n N_A_27_47#_c_329_n 0.0135685f $X=1.97 $Y=1.41 $X2=0
+ $Y2=0
cc_127 N_A_186_21#_c_118_n N_A_27_47#_c_329_n 0.0144997f $X=2.44 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A_186_21#_c_110_n N_A_27_47#_c_329_n 0.00461594f $X=2.445 $Y=1.16 $X2=0
+ $Y2=0
cc_129 N_A_186_21#_c_119_n N_A_27_47#_c_329_n 0.00955595f $X=4.25 $Y=2.317 $X2=0
+ $Y2=0
cc_130 N_A_186_21#_c_114_n N_A_27_47#_c_329_n 4.99213e-19 $X=2.44 $Y=1.202 $X2=0
+ $Y2=0
cc_131 N_A_186_21#_c_112_n N_A_27_47#_c_302_n 0.0108516f $X=4.25 $Y=0.74 $X2=0
+ $Y2=0
cc_132 N_A_186_21#_c_113_n N_A_27_47#_c_302_n 0.0418182f $X=4.352 $Y=2.21 $X2=0
+ $Y2=0
cc_133 N_A_186_21#_c_115_n N_A_27_47#_c_338_n 0.00166683f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_134 N_A_186_21#_c_115_n N_VPWR_c_389_n 0.01012f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_186_21#_c_116_n N_VPWR_c_389_n 0.00119371f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_186_21#_c_115_n N_VPWR_c_390_n 0.00132887f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_137 N_A_186_21#_c_116_n N_VPWR_c_390_n 0.0120673f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_186_21#_c_117_n N_VPWR_c_390_n 0.00900567f $X=1.97 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_186_21#_c_118_n N_VPWR_c_390_n 0.0011914f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_186_21#_c_117_n N_VPWR_c_391_n 0.00459627f $X=1.97 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_186_21#_c_118_n N_VPWR_c_391_n 0.00301372f $X=2.44 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_186_21#_c_117_n N_VPWR_c_392_n 0.00134018f $X=1.97 $Y=1.41 $X2=0
+ $Y2=0
cc_143 N_A_186_21#_c_118_n N_VPWR_c_392_n 0.012303f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_186_21#_c_115_n N_VPWR_c_394_n 0.00459627f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_145 N_A_186_21#_c_116_n N_VPWR_c_394_n 0.00315759f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_186_21#_c_119_n N_VPWR_c_395_n 0.0295899f $X=4.25 $Y=2.317 $X2=0
+ $Y2=0
cc_147 N_A_186_21#_M1005_d N_VPWR_c_388_n 0.00219934f $X=4 $Y=1.485 $X2=0 $Y2=0
cc_148 N_A_186_21#_c_115_n N_VPWR_c_388_n 0.00530041f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_149 N_A_186_21#_c_116_n N_VPWR_c_388_n 0.0038373f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_186_21#_c_117_n N_VPWR_c_388_n 0.00530041f $X=1.97 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_A_186_21#_c_118_n N_VPWR_c_388_n 0.00369099f $X=2.44 $Y=1.41 $X2=0
+ $Y2=0
cc_152 N_A_186_21#_c_119_n N_VPWR_c_388_n 0.0209375f $X=4.25 $Y=2.317 $X2=0
+ $Y2=0
cc_153 N_A_186_21#_c_106_n N_X_c_458_n 0.008232f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_186_21#_c_107_n N_X_c_458_n 0.0067113f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_186_21#_c_108_n N_X_c_458_n 5.41213e-19 $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_186_21#_c_106_n N_X_c_453_n 0.00203472f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_186_21#_c_115_n N_X_c_453_n 0.00739447f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_186_21#_c_107_n N_X_c_453_n 0.00213918f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_186_21#_c_110_n N_X_c_453_n 0.0131834f $X=2.445 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_186_21#_c_114_n N_X_c_453_n 0.0300086f $X=2.44 $Y=1.202 $X2=0 $Y2=0
cc_161 N_A_186_21#_c_107_n N_X_c_454_n 0.00883787f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_186_21#_c_108_n N_X_c_454_n 0.0119201f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_186_21#_c_109_n N_X_c_454_n 0.00139449f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_186_21#_c_110_n N_X_c_454_n 0.0582825f $X=2.445 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_186_21#_c_111_n N_X_c_454_n 0.0054731f $X=2.53 $Y=1.075 $X2=0 $Y2=0
cc_166 N_A_186_21#_c_193_p N_X_c_454_n 0.00679992f $X=2.615 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_186_21#_c_114_n N_X_c_454_n 0.00677781f $X=2.44 $Y=1.202 $X2=0 $Y2=0
cc_168 N_A_186_21#_c_107_n N_X_c_474_n 5.22855e-19 $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_186_21#_c_108_n N_X_c_474_n 0.00745779f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_186_21#_c_109_n N_X_c_474_n 0.00632002f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_186_21#_c_193_p N_X_c_474_n 0.00552965f $X=2.615 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_186_21#_c_106_n N_X_c_455_n 0.00259026f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_186_21#_c_107_n N_X_c_455_n 0.00140811f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_186_21#_c_114_n N_X_c_455_n 0.00124443f $X=2.44 $Y=1.202 $X2=0 $Y2=0
cc_175 N_A_186_21#_c_116_n X 0.0144287f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_186_21#_c_117_n X 0.0141219f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_186_21#_c_118_n X 0.0080627f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_186_21#_c_110_n X 0.0714913f $X=2.445 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_186_21#_c_114_n X 0.0202908f $X=2.44 $Y=1.202 $X2=0 $Y2=0
cc_180 N_A_186_21#_c_111_n N_VGND_M1013_s 7.2386e-19 $X=2.53 $Y=1.075 $X2=0
+ $Y2=0
cc_181 N_A_186_21#_c_112_n N_VGND_M1013_s 0.00762369f $X=4.25 $Y=0.74 $X2=0
+ $Y2=0
cc_182 N_A_186_21#_c_112_n N_VGND_M1006_d 0.00978829f $X=4.25 $Y=0.74 $X2=0
+ $Y2=0
cc_183 N_A_186_21#_c_106_n N_VGND_c_518_n 0.00419567f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_186_21#_c_107_n N_VGND_c_519_n 0.00428959f $X=1.475 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_186_21#_c_108_n N_VGND_c_519_n 0.00150539f $X=1.945 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_186_21#_c_108_n N_VGND_c_520_n 0.0043257f $X=1.945 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_186_21#_c_109_n N_VGND_c_520_n 0.00256701f $X=2.465 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_186_21#_c_193_p N_VGND_c_520_n 2.45707e-19 $X=2.615 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_186_21#_c_108_n N_VGND_c_521_n 5.00598e-19 $X=1.945 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A_186_21#_c_109_n N_VGND_c_521_n 0.0103593f $X=2.465 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_186_21#_c_112_n N_VGND_c_521_n 0.0143992f $X=4.25 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_186_21#_c_193_p N_VGND_c_521_n 0.00769258f $X=2.615 $Y=0.74 $X2=0
+ $Y2=0
cc_193 N_A_186_21#_c_112_n N_VGND_c_522_n 0.00805556f $X=4.25 $Y=0.74 $X2=0
+ $Y2=0
cc_194 N_A_186_21#_c_106_n N_VGND_c_523_n 0.00483491f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_186_21#_c_107_n N_VGND_c_523_n 0.00425617f $X=1.475 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_186_21#_c_112_n N_VGND_c_525_n 0.0102709f $X=4.25 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_186_21#_M1002_d N_VGND_c_526_n 0.00323135f $X=3.01 $Y=0.235 $X2=0
+ $Y2=0
cc_198 N_A_186_21#_M1003_d N_VGND_c_526_n 0.00373163f $X=3.96 $Y=0.235 $X2=0
+ $Y2=0
cc_199 N_A_186_21#_c_106_n N_VGND_c_526_n 0.00843259f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_186_21#_c_107_n N_VGND_c_526_n 0.00611453f $X=1.475 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_186_21#_c_108_n N_VGND_c_526_n 0.00619129f $X=1.945 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_186_21#_c_109_n N_VGND_c_526_n 0.00469928f $X=2.465 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_186_21#_c_112_n N_VGND_c_526_n 0.0339878f $X=4.25 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_186_21#_c_193_p N_VGND_c_526_n 0.00110938f $X=2.615 $Y=0.74 $X2=0
+ $Y2=0
cc_205 N_A_186_21#_c_112_n N_VGND_c_529_n 0.0245057f $X=4.25 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_c_234_n N_B_c_268_n 0.0260613f $X=2.935 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_207 N_A_c_233_n N_B_c_269_n 0.0790523f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_c_235_n N_B_c_269_n 0.00455145f $X=2.885 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_c_233_n B 7.4085e-19 $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_c_235_n B 0.0443909f $X=2.885 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_c_233_n N_A_27_47#_c_329_n 0.0144125f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_c_235_n N_A_27_47#_c_329_n 0.0179965f $X=2.885 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_c_233_n N_VPWR_c_392_n 0.0105202f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_c_233_n N_VPWR_c_395_n 0.0044524f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_c_233_n N_VPWR_c_388_n 0.00518028f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_c_233_n X 2.99822e-19 $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_c_235_n X 0.00783529f $X=2.885 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_c_235_n A_600_297# 0.00261226f $X=2.885 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_219 N_A_c_234_n N_VGND_c_521_n 0.00162962f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_c_234_n N_VGND_c_522_n 0.00428022f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_c_234_n N_VGND_c_526_n 0.00585784f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_c_234_n N_VGND_c_529_n 0.00120258f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_223 N_B_c_268_n N_A_27_47#_c_296_n 0.0177944f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B_c_269_n N_A_27_47#_c_297_n 0.0668347f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_225 B N_A_27_47#_c_297_n 0.00373847f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_226 N_B_c_269_n N_A_27_47#_c_329_n 0.0162978f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_227 B N_A_27_47#_c_329_n 0.0140478f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_228 N_B_c_269_n N_A_27_47#_c_302_n 0.00244642f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_229 B N_A_27_47#_c_302_n 0.0331895f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_230 N_B_c_269_n N_VPWR_c_392_n 0.00224847f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_231 N_B_c_269_n N_VPWR_c_395_n 0.00517927f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_232 N_B_c_269_n N_VPWR_c_388_n 0.00716671f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_233 B A_694_297# 0.0027975f $X=3.36 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_234 N_B_c_268_n N_VGND_c_522_n 0.00342417f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B_c_268_n N_VGND_c_526_n 0.00405449f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B_c_268_n N_VGND_c_529_n 0.00917505f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_301_n N_VPWR_M1009_d 0.00451385f $X=0.73 $Y=1.81 $X2=-0.19
+ $Y2=-0.24
cc_238 N_A_27_47#_c_329_n N_VPWR_M1009_d 0.00324693f $X=3.86 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_239 N_A_27_47#_c_338_n N_VPWR_M1009_d 0.00255548f $X=0.73 $Y=1.925 $X2=-0.19
+ $Y2=-0.24
cc_240 N_A_27_47#_c_329_n N_VPWR_M1004_d 0.00350347f $X=3.86 $Y=1.955 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_329_n N_VPWR_M1011_d 0.00774223f $X=3.86 $Y=1.955 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_329_n N_VPWR_c_389_n 0.00655922f $X=3.86 $Y=1.955 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_338_n N_VPWR_c_389_n 0.0144404f $X=0.73 $Y=1.925 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_329_n N_VPWR_c_390_n 0.0198977f $X=3.86 $Y=1.955 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_329_n N_VPWR_c_391_n 0.00768508f $X=3.86 $Y=1.955 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_329_n N_VPWR_c_392_n 0.0206216f $X=3.86 $Y=1.955 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_313_n N_VPWR_c_393_n 0.00337107f $X=0.645 $Y=1.925 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_306_n N_VPWR_c_393_n 0.00669761f $X=0.26 $Y=1.975 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_329_n N_VPWR_c_394_n 0.00775894f $X=3.86 $Y=1.955 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_297_n N_VPWR_c_395_n 0.00461156f $X=3.91 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_329_n N_VPWR_c_395_n 0.0142087f $X=3.86 $Y=1.955 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_297_n N_VPWR_c_388_n 0.00753486f $X=3.91 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_313_n N_VPWR_c_388_n 0.00706969f $X=0.645 $Y=1.925 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_329_n N_VPWR_c_388_n 0.0581071f $X=3.86 $Y=1.955 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_306_n N_VPWR_c_388_n 0.00838075f $X=0.26 $Y=1.975 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_338_n N_VPWR_c_388_n 7.87123e-19 $X=0.73 $Y=1.925 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_329_n N_X_M1000_s 0.00490491f $X=3.86 $Y=1.955 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_329_n N_X_M1007_s 0.00491654f $X=3.86 $Y=1.955 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_298_n N_X_c_458_n 0.00453622f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_301_n N_X_c_453_n 0.0540184f $X=0.73 $Y=1.81 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_329_n N_X_c_453_n 0.0158614f $X=3.86 $Y=1.955 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_299_n N_X_c_455_n 0.0133878f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_329_n X 0.0630657f $X=3.86 $Y=1.955 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_329_n A_600_297# 0.00849733f $X=3.86 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_265 N_A_27_47#_c_329_n A_694_297# 0.0114452f $X=3.86 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_266 N_A_27_47#_c_299_n N_VGND_M1010_d 0.00324145f $X=0.645 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_267 N_A_27_47#_c_298_n N_VGND_c_518_n 0.0128022f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_299_n N_VGND_c_518_n 0.0124847f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_296_n N_VGND_c_525_n 0.00342417f $X=3.885 $Y=0.995 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_M1010_s N_VGND_c_526_n 0.00302988f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_296_n N_VGND_c_526_n 0.00518989f $X=3.885 $Y=0.995 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_298_n N_VGND_c_526_n 0.00973659f $X=0.26 $Y=0.455 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_299_n N_VGND_c_526_n 0.00840262f $X=0.645 $Y=0.82 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_298_n N_VGND_c_527_n 0.01476f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_299_n N_VGND_c_527_n 0.00460418f $X=0.645 $Y=0.82 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_296_n N_VGND_c_529_n 0.0168594f $X=3.885 $Y=0.995 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_388_n N_X_M1000_s 0.00357693f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_c_388_n N_X_M1007_s 0.00357693f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_M1004_d X 0.00190556f $X=1.59 $Y=1.485 $X2=0 $Y2=0
cc_280 N_VPWR_c_388_n A_600_297# 0.00357693f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_281 N_VPWR_c_388_n A_694_297# 0.00431699f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_282 N_X_c_454_n N_VGND_M1008_s 0.00251598f $X=2.005 $Y=0.82 $X2=0 $Y2=0
cc_283 N_X_c_458_n N_VGND_c_518_n 0.0210691f $X=1.265 $Y=0.395 $X2=0 $Y2=0
cc_284 N_X_c_458_n N_VGND_c_519_n 0.0172733f $X=1.265 $Y=0.395 $X2=0 $Y2=0
cc_285 N_X_c_454_n N_VGND_c_519_n 0.0127122f $X=2.005 $Y=0.82 $X2=0 $Y2=0
cc_286 N_X_c_454_n N_VGND_c_520_n 0.00213422f $X=2.005 $Y=0.82 $X2=0 $Y2=0
cc_287 N_X_c_474_n N_VGND_c_520_n 0.0142956f $X=2.155 $Y=0.42 $X2=0 $Y2=0
cc_288 N_X_c_474_n N_VGND_c_521_n 0.0144215f $X=2.155 $Y=0.42 $X2=0 $Y2=0
cc_289 N_X_c_458_n N_VGND_c_523_n 0.0210662f $X=1.265 $Y=0.395 $X2=0 $Y2=0
cc_290 N_X_c_454_n N_VGND_c_523_n 0.00260082f $X=2.005 $Y=0.82 $X2=0 $Y2=0
cc_291 N_X_M1001_d N_VGND_c_526_n 0.00257127f $X=1.08 $Y=0.235 $X2=0 $Y2=0
cc_292 N_X_M1012_d N_VGND_c_526_n 0.00823216f $X=2.02 $Y=0.235 $X2=0 $Y2=0
cc_293 N_X_c_458_n N_VGND_c_526_n 0.0152475f $X=1.265 $Y=0.395 $X2=0 $Y2=0
cc_294 N_X_c_454_n N_VGND_c_526_n 0.00992881f $X=2.005 $Y=0.82 $X2=0 $Y2=0
cc_295 N_X_c_474_n N_VGND_c_526_n 0.00882622f $X=2.155 $Y=0.42 $X2=0 $Y2=0
