* File: sky130_fd_sc_hdll__dlrtn_1.spice
* Created: Thu Aug 27 19:05:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__dlrtn_1.pex.spice"
.subckt sky130_fd_sc_hdll__dlrtn_1  VNB VPB GATE_N D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* GATE_N	GATE_N
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_GATE_N_M1014_g N_A_27_363#_M1014_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_203_47#_M1002_d N_A_27_363#_M1002_g N_VGND_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_D_M1007_g N_A_319_369#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.1092 PD=0.715 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1018 A_500_47# N_A_319_369#_M1018_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.06195 PD=0.850769 PS=0.715 NRD=38.568 NRS=5.712 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1010 N_A_604_47#_M1010_d N_A_27_363#_M1010_g A_500_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0684 AS=0.0684 PD=0.729231 PS=0.729231 NRD=14.988 NRS=45 M=1 R=2.4
+ SA=75001.1 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1005 A_708_47# N_A_203_47#_M1005_g N_A_604_47#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0798 PD=0.63 PS=0.850769 NRD=14.28 NRS=12.852 M=1 R=2.8
+ SA=75001.5 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_750_21#_M1000_g A_708_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 A_981_47# N_A_604_47#_M1013_g N_A_750_21#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.082875 AS=0.169 PD=0.905 PS=1.82 NRD=13.38 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_RESET_B_M1009_g A_981_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.082875 PD=0.985 PS=0.905 NRD=6.456 NRS=13.38 M=1 R=4.33333
+ SA=75000.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1011 N_Q_M1011_d N_A_750_21#_M1011_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.108875 PD=1.82 PS=0.985 NRD=0 NRS=3.684 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_GATE_N_M1001_g N_A_27_363#_M1001_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1016 N_A_203_47#_M1016_d N_A_27_363#_M1016_g N_VPWR_M1001_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1008 N_VPWR_M1008_d N_D_M1008_g N_A_319_369#_M1008_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90002.8 A=0.1152 P=1.64 MULT=1
MM1004 A_503_369# N_A_319_369#_M1004_g N_VPWR_M1008_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.122023 AS=0.0928 PD=1.18943 PS=0.93 NRD=41.7443 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90002.4 A=0.1152 P=1.64 MULT=1
MM1017 N_A_604_47#_M1017_d N_A_203_47#_M1017_g A_503_369# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.0800774 PD=0.71 PS=0.780566 NRD=2.3443 NRS=63.631 M=1
+ R=2.33333 SA=90001.2 SB=90003 A=0.0756 P=1.2 MULT=1
MM1015 A_702_413# N_A_27_363#_M1015_g N_A_604_47#_M1017_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.063 AS=0.0609 PD=0.72 PS=0.71 NRD=44.5417 NRS=2.3443 M=1 R=2.33333
+ SA=90001.6 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1003 N_VPWR_M1003_d N_A_750_21#_M1003_g A_702_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.138955 AS=0.063 PD=1.02042 PS=0.72 NRD=2.3443 NRS=44.5417 M=1 R=2.33333
+ SA=90002.1 SB=90002 A=0.0756 P=1.2 MULT=1
MM1019 N_A_750_21#_M1019_d N_A_604_47#_M1019_g N_VPWR_M1003_d VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.330845 PD=1.29 PS=2.42958 NRD=0.9653 NRS=5.8903 M=1
+ R=5.55556 SA=90001.4 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_RESET_B_M1012_g N_A_750_21#_M1019_d VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.9 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1006 N_Q_M1006_d N_A_750_21#_M1006_g N_VPWR_M1012_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
c_131 VPB 0 1.5379e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__dlrtn_1.pxi.spice"
*
.ends
*
*
