* File: sky130_fd_sc_hdll__a22o_1.spice
* Created: Wed Sep  2 08:18:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a22o_1.pex.spice"
.subckt sky130_fd_sc_hdll__a22o_1  VNB VPB B2 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1009 A_119_47# N_B2_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.2015 PD=0.92 PS=1.92 NRD=14.76 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_297#_M1002_d N_B1_M1002_g A_119_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0.912 NRS=14.76 M=1 R=4.33333
+ SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 A_411_47# N_A1_M1004_g N_A_27_297#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.221 PD=1.02 PS=1.98 NRD=23.988 NRS=13.836 M=1 R=4.33333
+ SA=75000.3 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_411_47# VNB NSHORT L=0.15 W=0.65 AD=0.117
+ AS=0.12025 PD=1.01 PS=1.02 NRD=6.456 NRS=23.988 M=1 R=4.33333 SA=75000.8
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_27_297#_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.26 AS=0.117 PD=2.1 PS=1.01 NRD=24.912 NRS=8.304 M=1 R=4.33333 SA=75001.3
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1003 N_A_117_297#_M1003_d N_B2_M1003_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1000 N_A_27_297#_M1000_d N_B1_M1000_g N_A_117_297#_M1003_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_A_117_297#_M1008_d N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.17 AS=0.27 PD=1.34 PS=2.54 NRD=5.8903 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_117_297#_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.165 AS=0.17 PD=1.33 PS=1.34 NRD=8.8453 NRS=5.8903 M=1 R=5.55556
+ SA=90000.7 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1007 N_X_M1007_d N_A_27_297#_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.41 AS=0.165 PD=2.82 PS=1.33 NRD=28.565 NRS=0.9653 M=1 R=5.55556
+ SA=90001.2 SB=90000.3 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hdll__a22o_1.pxi.spice"
*
.ends
*
*
