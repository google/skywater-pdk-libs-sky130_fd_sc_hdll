* File: sky130_fd_sc_hdll__nor4_6.spice
* Created: Wed Sep  2 08:41:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor4_6.pex.spice"
.subckt sky130_fd_sc_hdll__nor4_6  VNB VPB A B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65 AD=0.2145
+ AS=0.08775 PD=1.96 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.3 SB=75011.5
+ A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75011.1 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1011_d N_A_M1019_g N_Y_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75010.6 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A_M1021_g N_Y_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75010.2 A=0.0975 P=1.6 MULT=1
MM1026 N_VGND_M1021_d N_A_M1026_g N_Y_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75009.7 A=0.0975 P=1.6 MULT=1
MM1034 N_VGND_M1034_d N_A_M1034_g N_Y_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75009.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1034_d N_B_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75008.7 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_B_M1008_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75008.3 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1008_d N_B_M1012_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75007.8 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1022_d N_B_M1022_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75007.4 A=0.0975 P=1.6 MULT=1
MM1036 N_VGND_M1022_d N_B_M1036_g N_Y_M1036_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005
+ SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1046 N_VGND_M1046_d N_B_M1046_g N_Y_M1036_s VNB NSHORT L=0.15 W=0.65
+ AD=0.28925 AS=0.08775 PD=1.54 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.4
+ SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1046_d N_C_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.28925 AS=0.08775 PD=1.54 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006.4
+ SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_C_M1013_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006.8
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1028 N_VGND_M1013_d N_C_M1028_g N_Y_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75007.4
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1038 N_VGND_M1038_d N_C_M1038_g N_Y_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75007.8
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1039 N_VGND_M1038_d N_C_M1039_g N_Y_M1039_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75008.3
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1044 N_VGND_M1044_d N_C_M1044_g N_Y_M1039_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75008.7
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_D_M1004_g N_VGND_M1044_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75009.2
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1004_d N_D_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75009.7
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1025 N_Y_M1025_d N_D_M1025_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75010.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1032 N_Y_M1025_d N_D_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75010.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1041 N_Y_M1041_d N_D_M1041_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75011.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1047 N_Y_M1041_d N_D_M1047_g N_VGND_M1047_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.221 PD=0.92 PS=1.98 NRD=0 NRS=10.152 M=1 R=4.33333 SA=75011.5
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_27_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90005.3 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1000_d N_A_M1005_g N_A_27_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_A_27_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1014_d N_A_M1020_g N_A_27_297#_M1020_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90003.9 A=0.18 P=2.36 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_A_27_297#_M1020_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1042 N_VPWR_M1030_d N_A_M1042_g N_A_27_297#_M1042_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90003 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1042_s N_B_M1009_g N_A_685_297#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1017 N_A_27_297#_M1017_d N_B_M1017_g N_A_685_297#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1024 N_A_27_297#_M1017_d N_B_M1024_g N_A_685_297#_M1024_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1033 N_A_27_297#_M1033_d N_B_M1033_g N_A_685_297#_M1024_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1035 N_A_27_297#_M1033_d N_B_M1035_g N_A_685_297#_M1035_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.9 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1040 N_A_27_297#_M1040_d N_B_M1040_g N_A_685_297#_M1035_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.4 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_1263_297#_M1001_d N_C_M1001_g N_A_685_297#_M1001_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90005.4 A=0.18 P=2.36 MULT=1
MM1007 N_A_1263_297#_M1007_d N_C_M1007_g N_A_685_297#_M1001_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1015 N_A_1263_297#_M1007_d N_C_M1015_g N_A_685_297#_M1015_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1016 N_A_1263_297#_M1016_d N_C_M1016_g N_A_685_297#_M1015_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90004 A=0.18 P=2.36 MULT=1
MM1043 N_A_1263_297#_M1016_d N_C_M1043_g N_A_685_297#_M1043_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1045 N_A_1263_297#_M1045_d N_C_M1045_g N_A_685_297#_M1043_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90003 A=0.18 P=2.36 MULT=1
MM1002 N_Y_M1002_d N_D_M1002_g N_A_1263_297#_M1045_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1018 N_Y_M1002_d N_D_M1018_g N_A_1263_297#_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1027 N_Y_M1027_d N_D_M1027_g N_A_1263_297#_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.9 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1029 N_Y_M1027_d N_D_M1029_g N_A_1263_297#_M1029_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1031 N_Y_M1031_d N_D_M1031_g N_A_1263_297#_M1029_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.9 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1037 N_Y_M1031_d N_D_M1037_g N_A_1263_297#_M1037_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.3 PD=1.29 PS=2.6 NRD=0.9653 NRS=2.9353 M=1 R=5.55556 SA=90005.3
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX48_noxref VNB VPB NWDIODE A=20.544 P=28.81
*
.include "sky130_fd_sc_hdll__nor4_6.pxi.spice"
*
.ends
*
*
