* File: sky130_fd_sc_hdll__muxb16to1_1.pex.spice
* Created: Thu Aug 27 19:11:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[0] 1 3 4 6 8 13 15
c29 4 0 5.33021e-20 $X=0.495 $Y=1.41
r30 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.69 $Y=0.51
+ $X2=0.645 $Y2=0.51
r31 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.5 $Y=1.19
+ $X2=0.645 $Y2=1.19
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.5
+ $Y=1.16 $X2=0.5 $Y2=1.16
r33 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.645 $Y=1.055
+ $X2=0.645 $Y2=1.19
r34 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.645 $Y=0.625
+ $X2=0.645 $Y2=0.51
r35 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.645 $Y=0.625
+ $X2=0.645 $Y2=1.055
r36 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.5 $Y2=1.16
r37 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r38 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.5 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[8] 1 3 4 6 8 13 15
c31 1 0 5.33021e-20 $X=0.47 $Y=4.445
r32 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.69 $Y=4.93
+ $X2=0.645 $Y2=4.93
r33 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.5 $Y=4.25
+ $X2=0.645 $Y2=4.25
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.5
+ $Y=4.28 $X2=0.5 $Y2=4.28
r35 8 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.645 $Y=4.815
+ $X2=0.645 $Y2=4.93
r36 7 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.645 $Y=4.385
+ $X2=0.645 $Y2=4.25
r37 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.645 $Y=4.385
+ $X2=0.645 $Y2=4.815
r38 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.495 $Y=4.03
+ $X2=0.5 $Y2=4.28
r39 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=4.03
+ $X2=0.495 $Y2=3.455
r40 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=0.47 $Y=4.445
+ $X2=0.5 $Y2=4.28
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=4.445 $X2=0.47
+ $Y2=4.88
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_184_265# 1 2 9 11 12 15 22 26
r58 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=1.545 $Y=1.405
+ $X2=1.775 $Y2=1.63
r59 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=1.325 $Y=1.34
+ $X2=1.02 $Y2=1.34
r60 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=1.325 $Y=1.405
+ $X2=1.545 $Y2=1.405
r61 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.34 $X2=1.325 $Y2=1.34
r62 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.775 $Y=2.31
+ $X2=1.775 $Y2=1.635
r63 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.545 $Y=1.175
+ $X2=1.545 $Y2=1.405
r64 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=1.545 $Y=0.755
+ $X2=1.775 $Y2=0.542
r65 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.545 $Y=0.755
+ $X2=1.545 $Y2=1.175
r66 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.02 $Y=1.475
+ $X2=1.02 $Y2=1.34
r67 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.02 $Y=1.475 $X2=1.02
+ $Y2=2.075
r68 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.485 $X2=1.775 $Y2=1.63
r69 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.485 $X2=1.775 $Y2=2.31
r70 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=0.235 $X2=1.775 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_184_793# 1 2 9 12 13 15 26
r56 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=1.325 $Y=4.1
+ $X2=1.02 $Y2=4.1
r57 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=1.325 $Y=4.035
+ $X2=1.545 $Y2=4.035
r58 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=4.1 $X2=1.325 $Y2=4.1
r59 13 20 9.67586 $w=2.9e-07 $l=3.25269e-07 $layer=LI1_cond $X=1.775 $Y=3.805
+ $X2=1.545 $Y2=4.035
r60 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.775 $Y=3.805
+ $X2=1.775 $Y2=3.13
r61 12 25 8.93631 $w=3.14e-07 $l=3.18842e-07 $layer=LI1_cond $X=1.545 $Y=4.685
+ $X2=1.775 $Y2=4.897
r62 11 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.545 $Y=4.265
+ $X2=1.545 $Y2=4.035
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.545 $Y=4.265
+ $X2=1.545 $Y2=4.685
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.02 $Y=3.965
+ $X2=1.02 $Y2=4.1
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.02 $Y=3.965 $X2=1.02
+ $Y2=3.365
r66 2 13 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=2.955 $X2=1.775 $Y2=3.81
r67 2 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=2.955 $X2=1.775 $Y2=3.13
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=4.685 $X2=1.775 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[0] 1 3 4 5 6 8 9 11 12 17
r49 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.975
+ $Y=1.03 $X2=1.975 $Y2=1.03
r50 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=1.975 $Y=0.905
+ $X2=1.975 $Y2=1.03
r51 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.005 $Y=1.19
+ $X2=2.005 $Y2=1.03
r52 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.01 $Y=0.83
+ $X2=1.975 $Y2=0.905
r53 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.01 $Y=0.83
+ $X2=2.01 $Y2=0.495
r54 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=2.01 $Y=1.41
+ $X2=1.975 $Y2=1.03
r55 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.01 $Y=1.41 $X2=2.01
+ $Y2=1.985
r56 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.84 $Y=0.905
+ $X2=1.975 $Y2=0.905
r57 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.84 $Y=0.905 $X2=1.02
+ $Y2=0.905
r58 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.945 $Y=0.83
+ $X2=1.02 $Y2=0.905
r59 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.945 $Y=0.83
+ $X2=0.945 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[8] 1 3 4 5 6 8 9 11 12
r48 15 17 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=1.975 $Y=4.41
+ $X2=1.975 $Y2=4.535
r49 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.975
+ $Y=4.41 $X2=1.975 $Y2=4.41
r50 12 16 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.005 $Y=4.25
+ $X2=2.005 $Y2=4.41
r51 9 17 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.01 $Y=4.61
+ $X2=1.975 $Y2=4.535
r52 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.01 $Y=4.61
+ $X2=2.01 $Y2=4.945
r53 6 15 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=2.01 $Y=4.03
+ $X2=1.975 $Y2=4.41
r54 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.01 $Y=4.03 $X2=2.01
+ $Y2=3.455
r55 4 17 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.84 $Y=4.535
+ $X2=1.975 $Y2=4.535
r56 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.84 $Y=4.535 $X2=1.02
+ $Y2=4.535
r57 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.945 $Y=4.61
+ $X2=1.02 $Y2=4.535
r58 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.945 $Y=4.61
+ $X2=0.945 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[1] 1 3 4 6 7 9 11 12 17
r46 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.03 $X2=2.625 $Y2=1.03
r47 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=2.625 $Y=0.905
+ $X2=2.625 $Y2=1.03
r48 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.595 $Y=1.19
+ $X2=2.595 $Y2=1.03
r49 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.655 $Y=0.83
+ $X2=3.655 $Y2=0.495
r50 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.76 $Y=0.905
+ $X2=2.625 $Y2=0.905
r51 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.58 $Y=0.905
+ $X2=3.655 $Y2=0.83
r52 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.58 $Y=0.905 $X2=2.76
+ $Y2=0.905
r53 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.59 $Y=0.83
+ $X2=2.625 $Y2=0.905
r54 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.59 $Y=0.83 $X2=2.59
+ $Y2=0.495
r55 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=2.59 $Y=1.41
+ $X2=2.625 $Y2=1.03
r56 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.59 $Y=1.41 $X2=2.59
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[9] 1 3 4 6 7 9 11 12
r47 15 17 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=2.625 $Y=4.41
+ $X2=2.625 $Y2=4.535
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=4.41 $X2=2.625 $Y2=4.41
r49 12 16 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.595 $Y=4.25
+ $X2=2.595 $Y2=4.41
r50 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.655 $Y=4.61
+ $X2=3.655 $Y2=4.945
r51 8 17 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.76 $Y=4.535
+ $X2=2.625 $Y2=4.535
r52 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.58 $Y=4.535
+ $X2=3.655 $Y2=4.61
r53 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.58 $Y=4.535 $X2=2.76
+ $Y2=4.535
r54 4 17 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.59 $Y=4.61
+ $X2=2.625 $Y2=4.535
r55 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.59 $Y=4.61 $X2=2.59
+ $Y2=4.945
r56 1 15 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=2.59 $Y=4.03
+ $X2=2.625 $Y2=4.41
r57 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.59 $Y=4.03 $X2=2.59
+ $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_533_47# 1 2 9 13 16 19 22 24
r57 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=3.275 $Y=1.34
+ $X2=3.58 $Y2=1.34
r58 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.275
+ $Y=1.34 $X2=3.275 $Y2=1.34
r59 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=3.055 $Y=1.405
+ $X2=3.275 $Y2=1.405
r60 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=2.825 $Y=1.63
+ $X2=3.055 $Y2=1.405
r61 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.055 $Y=1.175
+ $X2=3.055 $Y2=1.405
r62 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=3.055 $Y=0.755
+ $X2=2.825 $Y2=0.542
r63 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.055 $Y=0.755
+ $X2=3.055 $Y2=1.175
r64 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.825 $Y=2.31
+ $X2=2.825 $Y2=1.635
r65 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=3.58 $Y=1.475
+ $X2=3.58 $Y2=1.34
r66 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=3.58 $Y=1.475 $X2=3.58
+ $Y2=2.075
r67 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.485 $X2=2.825 $Y2=1.63
r68 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.485 $X2=2.825 $Y2=2.31
r69 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.825 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_533_937# 1 2 9 13 16 19 22 24
r59 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=3.275 $Y=4.1
+ $X2=3.58 $Y2=4.1
r60 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.275
+ $Y=4.1 $X2=3.275 $Y2=4.1
r61 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=3.055 $Y=4.035
+ $X2=3.275 $Y2=4.035
r62 16 24 8.93631 $w=3.14e-07 $l=3.18842e-07 $layer=LI1_cond $X=3.055 $Y=4.685
+ $X2=2.825 $Y2=4.897
r63 15 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.055 $Y=4.265
+ $X2=3.055 $Y2=4.035
r64 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.055 $Y=4.265
+ $X2=3.055 $Y2=4.685
r65 11 19 9.67586 $w=2.9e-07 $l=3.25269e-07 $layer=LI1_cond $X=2.825 $Y=3.805
+ $X2=3.055 $Y2=4.035
r66 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.825 $Y=3.805
+ $X2=2.825 $Y2=3.13
r67 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=3.58 $Y=3.965
+ $X2=3.58 $Y2=4.1
r68 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=3.58 $Y=3.965 $X2=3.58
+ $Y2=3.365
r69 2 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=2.955 $X2=2.825 $Y2=3.81
r70 2 13 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=2.955 $X2=2.825 $Y2=3.13
r71 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=4.685 $X2=2.825 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[1] 1 3 4 6 8 12 15 21
c38 8 0 1.78369e-19 $X=3.955 $Y=1.055
c39 1 0 2.31671e-19 $X=4.105 $Y=1.41
r40 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.91 $Y=0.51
+ $X2=3.955 $Y2=0.51
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.1
+ $Y=1.16 $X2=4.1 $Y2=1.16
r42 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.955 $Y=1.19
+ $X2=4.1 $Y2=1.19
r43 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.955 $Y=1.055
+ $X2=3.955 $Y2=1.19
r44 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.955 $Y=0.625
+ $X2=3.955 $Y2=0.51
r45 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.955 $Y=0.625
+ $X2=3.955 $Y2=1.055
r46 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.13 $Y=0.995
+ $X2=4.1 $Y2=1.16
r47 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.13 $Y=0.995 $X2=4.13
+ $Y2=0.56
r48 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=4.105 $Y=1.41
+ $X2=4.1 $Y2=1.16
r49 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.105 $Y=1.41
+ $X2=4.105 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[9] 1 3 4 6 8 12 15 21
c41 8 0 1.78369e-19 $X=3.955 $Y=4.815
c42 4 0 2.31671e-19 $X=4.13 $Y=4.445
r43 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.91 $Y=4.93
+ $X2=3.955 $Y2=4.93
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.1
+ $Y=4.28 $X2=4.1 $Y2=4.28
r45 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.955 $Y=4.25
+ $X2=4.1 $Y2=4.25
r46 8 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.955 $Y=4.815
+ $X2=3.955 $Y2=4.93
r47 7 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.955 $Y=4.385
+ $X2=3.955 $Y2=4.25
r48 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.955 $Y=4.385
+ $X2=3.955 $Y2=4.815
r49 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.13 $Y=4.445
+ $X2=4.1 $Y2=4.28
r50 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.13 $Y=4.445 $X2=4.13
+ $Y2=4.88
r51 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=4.105 $Y=4.03
+ $X2=4.1 $Y2=4.28
r52 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.105 $Y=4.03
+ $X2=4.105 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[2] 1 3 4 6 8 13 15
c38 8 0 1.78369e-19 $X=4.785 $Y=1.055
c39 4 0 2.31671e-19 $X=4.635 $Y=1.41
r40 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.83 $Y=0.51
+ $X2=4.785 $Y2=0.51
r41 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.64 $Y=1.19
+ $X2=4.785 $Y2=1.19
r42 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.64
+ $Y=1.16 $X2=4.64 $Y2=1.16
r43 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.785 $Y=1.055
+ $X2=4.785 $Y2=1.19
r44 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.785 $Y=0.625
+ $X2=4.785 $Y2=0.51
r45 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.785 $Y=0.625
+ $X2=4.785 $Y2=1.055
r46 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=4.635 $Y=1.41
+ $X2=4.64 $Y2=1.16
r47 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.635 $Y=1.41
+ $X2=4.635 $Y2=1.985
r48 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.61 $Y=0.995
+ $X2=4.64 $Y2=1.16
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.61 $Y=0.995 $X2=4.61
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[10] 1 3 4 6 8 13 15
c41 8 0 1.78369e-19 $X=4.785 $Y=4.815
c42 1 0 2.31671e-19 $X=4.61 $Y=4.445
r43 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.83 $Y=4.93
+ $X2=4.785 $Y2=4.93
r44 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.64 $Y=4.25
+ $X2=4.785 $Y2=4.25
r45 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.64
+ $Y=4.28 $X2=4.64 $Y2=4.28
r46 8 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.785 $Y=4.815
+ $X2=4.785 $Y2=4.93
r47 7 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.785 $Y=4.385
+ $X2=4.785 $Y2=4.25
r48 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.785 $Y=4.385
+ $X2=4.785 $Y2=4.815
r49 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=4.635 $Y=4.03
+ $X2=4.64 $Y2=4.28
r50 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.635 $Y=4.03
+ $X2=4.635 $Y2=3.455
r51 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.61 $Y=4.445
+ $X2=4.64 $Y2=4.28
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.61 $Y=4.445 $X2=4.61
+ $Y2=4.88
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1012_265# 1 2 9 11 12 15 22 26
r58 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=5.685 $Y=1.405
+ $X2=5.915 $Y2=1.63
r59 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=5.465 $Y=1.34
+ $X2=5.16 $Y2=1.34
r60 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=5.465 $Y=1.405
+ $X2=5.685 $Y2=1.405
r61 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.465
+ $Y=1.34 $X2=5.465 $Y2=1.34
r62 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.915 $Y=2.31
+ $X2=5.915 $Y2=1.635
r63 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.685 $Y=1.175
+ $X2=5.685 $Y2=1.405
r64 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=5.685 $Y=0.755
+ $X2=5.915 $Y2=0.542
r65 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.685 $Y=0.755
+ $X2=5.685 $Y2=1.175
r66 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.16 $Y=1.475
+ $X2=5.16 $Y2=1.34
r67 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=5.16 $Y=1.475 $X2=5.16
+ $Y2=2.075
r68 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.485 $X2=5.915 $Y2=1.63
r69 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.485 $X2=5.915 $Y2=2.31
r70 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=5.79
+ $Y=0.235 $X2=5.915 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1012_793# 1 2 9 12 13 15 26
r56 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=5.465 $Y=4.1
+ $X2=5.16 $Y2=4.1
r57 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=5.465 $Y=4.035
+ $X2=5.685 $Y2=4.035
r58 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.465
+ $Y=4.1 $X2=5.465 $Y2=4.1
r59 13 20 9.67586 $w=2.9e-07 $l=3.25269e-07 $layer=LI1_cond $X=5.915 $Y=3.805
+ $X2=5.685 $Y2=4.035
r60 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.915 $Y=3.805
+ $X2=5.915 $Y2=3.13
r61 12 25 8.93631 $w=3.14e-07 $l=3.18842e-07 $layer=LI1_cond $X=5.685 $Y=4.685
+ $X2=5.915 $Y2=4.897
r62 11 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.685 $Y=4.265
+ $X2=5.685 $Y2=4.035
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.685 $Y=4.265
+ $X2=5.685 $Y2=4.685
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.16 $Y=3.965
+ $X2=5.16 $Y2=4.1
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=5.16 $Y=3.965 $X2=5.16
+ $Y2=3.365
r66 2 13 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=2.955 $X2=5.915 $Y2=3.81
r67 2 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=2.955 $X2=5.915 $Y2=3.13
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=5.79
+ $Y=4.685 $X2=5.915 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[2] 1 3 4 5 6 8 9 11 12 17
r49 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.115
+ $Y=1.03 $X2=6.115 $Y2=1.03
r50 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=6.115 $Y=0.905
+ $X2=6.115 $Y2=1.03
r51 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=6.145 $Y=1.19
+ $X2=6.145 $Y2=1.03
r52 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.15 $Y=0.83
+ $X2=6.115 $Y2=0.905
r53 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.15 $Y=0.83
+ $X2=6.15 $Y2=0.495
r54 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=6.15 $Y=1.41
+ $X2=6.115 $Y2=1.03
r55 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.15 $Y=1.41 $X2=6.15
+ $Y2=1.985
r56 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.98 $Y=0.905
+ $X2=6.115 $Y2=0.905
r57 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.98 $Y=0.905 $X2=5.16
+ $Y2=0.905
r58 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.085 $Y=0.83
+ $X2=5.16 $Y2=0.905
r59 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.085 $Y=0.83
+ $X2=5.085 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[10] 1 3 4 5 6 8 9 11 12
r48 15 17 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=6.115 $Y=4.41
+ $X2=6.115 $Y2=4.535
r49 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.115
+ $Y=4.41 $X2=6.115 $Y2=4.41
r50 12 16 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=6.145 $Y=4.25
+ $X2=6.145 $Y2=4.41
r51 9 17 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.15 $Y=4.61
+ $X2=6.115 $Y2=4.535
r52 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.15 $Y=4.61
+ $X2=6.15 $Y2=4.945
r53 6 15 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=6.15 $Y=4.03
+ $X2=6.115 $Y2=4.41
r54 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.15 $Y=4.03 $X2=6.15
+ $Y2=3.455
r55 4 17 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.98 $Y=4.535
+ $X2=6.115 $Y2=4.535
r56 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.98 $Y=4.535 $X2=5.16
+ $Y2=4.535
r57 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.085 $Y=4.61
+ $X2=5.16 $Y2=4.535
r58 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.085 $Y=4.61
+ $X2=5.085 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[3] 1 3 4 6 7 9 11 12 17
r46 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.765
+ $Y=1.03 $X2=6.765 $Y2=1.03
r47 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=6.765 $Y=0.905
+ $X2=6.765 $Y2=1.03
r48 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=6.735 $Y=1.19
+ $X2=6.735 $Y2=1.03
r49 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.795 $Y=0.83
+ $X2=7.795 $Y2=0.495
r50 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.9 $Y=0.905
+ $X2=6.765 $Y2=0.905
r51 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.72 $Y=0.905
+ $X2=7.795 $Y2=0.83
r52 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.72 $Y=0.905 $X2=6.9
+ $Y2=0.905
r53 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.73 $Y=0.83
+ $X2=6.765 $Y2=0.905
r54 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.73 $Y=0.83 $X2=6.73
+ $Y2=0.495
r55 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=6.73 $Y=1.41
+ $X2=6.765 $Y2=1.03
r56 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.73 $Y=1.41 $X2=6.73
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[11] 1 3 4 6 7 9 11 12
r47 15 17 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=6.765 $Y=4.41
+ $X2=6.765 $Y2=4.535
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.765
+ $Y=4.41 $X2=6.765 $Y2=4.41
r49 12 16 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=6.735 $Y=4.25
+ $X2=6.735 $Y2=4.41
r50 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.795 $Y=4.61
+ $X2=7.795 $Y2=4.945
r51 8 17 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.9 $Y=4.535
+ $X2=6.765 $Y2=4.535
r52 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.72 $Y=4.535
+ $X2=7.795 $Y2=4.61
r53 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.72 $Y=4.535 $X2=6.9
+ $Y2=4.535
r54 4 17 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.73 $Y=4.61
+ $X2=6.765 $Y2=4.535
r55 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.73 $Y=4.61 $X2=6.73
+ $Y2=4.945
r56 1 15 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=6.73 $Y=4.03
+ $X2=6.765 $Y2=4.41
r57 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.73 $Y=4.03 $X2=6.73
+ $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1361_47# 1 2 9 13 16 19 22 24
r57 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=7.415 $Y=1.34
+ $X2=7.72 $Y2=1.34
r58 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.415
+ $Y=1.34 $X2=7.415 $Y2=1.34
r59 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=7.195 $Y=1.405
+ $X2=7.415 $Y2=1.405
r60 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=6.965 $Y=1.63
+ $X2=7.195 $Y2=1.405
r61 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.195 $Y=1.175
+ $X2=7.195 $Y2=1.405
r62 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=7.195 $Y=0.755
+ $X2=6.965 $Y2=0.542
r63 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.195 $Y=0.755
+ $X2=7.195 $Y2=1.175
r64 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.965 $Y=2.31
+ $X2=6.965 $Y2=1.635
r65 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.72 $Y=1.475
+ $X2=7.72 $Y2=1.34
r66 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=7.72 $Y=1.475 $X2=7.72
+ $Y2=2.075
r67 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.485 $X2=6.965 $Y2=1.63
r68 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.485 $X2=6.965 $Y2=2.31
r69 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.235 $X2=6.965 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1361_937# 1 2 9 13 16 19 22 24
r59 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=7.415 $Y=4.1
+ $X2=7.72 $Y2=4.1
r60 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.415
+ $Y=4.1 $X2=7.415 $Y2=4.1
r61 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=7.195 $Y=4.035
+ $X2=7.415 $Y2=4.035
r62 16 24 8.93631 $w=3.14e-07 $l=3.18842e-07 $layer=LI1_cond $X=7.195 $Y=4.685
+ $X2=6.965 $Y2=4.897
r63 15 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.195 $Y=4.265
+ $X2=7.195 $Y2=4.035
r64 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.195 $Y=4.265
+ $X2=7.195 $Y2=4.685
r65 11 19 9.67586 $w=2.9e-07 $l=3.25269e-07 $layer=LI1_cond $X=6.965 $Y=3.805
+ $X2=7.195 $Y2=4.035
r66 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.965 $Y=3.805
+ $X2=6.965 $Y2=3.13
r67 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.72 $Y=3.965
+ $X2=7.72 $Y2=4.1
r68 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=7.72 $Y=3.965 $X2=7.72
+ $Y2=3.365
r69 2 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=2.955 $X2=6.965 $Y2=3.81
r70 2 13 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=2.955 $X2=6.965 $Y2=3.13
r71 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=4.685 $X2=6.965 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[3] 1 3 4 6 8 12 15 21
c38 8 0 1.78369e-19 $X=8.095 $Y=1.055
c39 1 0 2.31671e-19 $X=8.245 $Y=1.41
r40 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.05 $Y=0.51
+ $X2=8.095 $Y2=0.51
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.24
+ $Y=1.16 $X2=8.24 $Y2=1.16
r42 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.095 $Y=1.19
+ $X2=8.24 $Y2=1.19
r43 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.095 $Y=1.055
+ $X2=8.095 $Y2=1.19
r44 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.095 $Y=0.625
+ $X2=8.095 $Y2=0.51
r45 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.095 $Y=0.625
+ $X2=8.095 $Y2=1.055
r46 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=8.27 $Y=0.995
+ $X2=8.24 $Y2=1.16
r47 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.27 $Y=0.995 $X2=8.27
+ $Y2=0.56
r48 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=8.245 $Y=1.41
+ $X2=8.24 $Y2=1.16
r49 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.245 $Y=1.41
+ $X2=8.245 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[11] 1 3 4 6 8 12 15 21
c41 8 0 1.78369e-19 $X=8.095 $Y=4.815
c42 4 0 2.31671e-19 $X=8.27 $Y=4.445
r43 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.05 $Y=4.93
+ $X2=8.095 $Y2=4.93
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.24
+ $Y=4.28 $X2=8.24 $Y2=4.28
r45 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.095 $Y=4.25
+ $X2=8.24 $Y2=4.25
r46 8 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.095 $Y=4.815
+ $X2=8.095 $Y2=4.93
r47 7 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.095 $Y=4.385
+ $X2=8.095 $Y2=4.25
r48 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.095 $Y=4.385
+ $X2=8.095 $Y2=4.815
r49 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=8.27 $Y=4.445
+ $X2=8.24 $Y2=4.28
r50 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.27 $Y=4.445 $X2=8.27
+ $Y2=4.88
r51 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=8.245 $Y=4.03
+ $X2=8.24 $Y2=4.28
r52 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.245 $Y=4.03
+ $X2=8.245 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[4] 1 3 4 6 8 13 15
c38 8 0 1.78369e-19 $X=8.925 $Y=1.055
c39 4 0 2.31671e-19 $X=8.775 $Y=1.41
r40 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.97 $Y=0.51
+ $X2=8.925 $Y2=0.51
r41 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.78 $Y=1.19
+ $X2=8.925 $Y2=1.19
r42 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.78
+ $Y=1.16 $X2=8.78 $Y2=1.16
r43 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.925 $Y=1.055
+ $X2=8.925 $Y2=1.19
r44 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.925 $Y=0.625
+ $X2=8.925 $Y2=0.51
r45 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.925 $Y=0.625
+ $X2=8.925 $Y2=1.055
r46 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=8.775 $Y=1.41
+ $X2=8.78 $Y2=1.16
r47 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.775 $Y=1.41
+ $X2=8.775 $Y2=1.985
r48 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=8.75 $Y=0.995
+ $X2=8.78 $Y2=1.16
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.75 $Y=0.995 $X2=8.75
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[12] 1 3 4 6 8 13 15
c41 8 0 1.78369e-19 $X=8.925 $Y=4.815
c42 1 0 2.31671e-19 $X=8.75 $Y=4.445
r43 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.97 $Y=4.93
+ $X2=8.925 $Y2=4.93
r44 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.78 $Y=4.25
+ $X2=8.925 $Y2=4.25
r45 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.78
+ $Y=4.28 $X2=8.78 $Y2=4.28
r46 8 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.925 $Y=4.815
+ $X2=8.925 $Y2=4.93
r47 7 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.925 $Y=4.385
+ $X2=8.925 $Y2=4.25
r48 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.925 $Y=4.385
+ $X2=8.925 $Y2=4.815
r49 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=8.775 $Y=4.03
+ $X2=8.78 $Y2=4.28
r50 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.775 $Y=4.03
+ $X2=8.775 $Y2=3.455
r51 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=8.75 $Y=4.445
+ $X2=8.78 $Y2=4.28
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.75 $Y=4.445 $X2=8.75
+ $Y2=4.88
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1840_265# 1 2 9 11 12 15 22 26
r58 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=9.825 $Y=1.405
+ $X2=10.055 $Y2=1.63
r59 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=9.605 $Y=1.34
+ $X2=9.3 $Y2=1.34
r60 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=9.605 $Y=1.405
+ $X2=9.825 $Y2=1.405
r61 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.605
+ $Y=1.34 $X2=9.605 $Y2=1.34
r62 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.055 $Y=2.31
+ $X2=10.055 $Y2=1.635
r63 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=9.825 $Y=1.175
+ $X2=9.825 $Y2=1.405
r64 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=9.825 $Y=0.755
+ $X2=10.055 $Y2=0.542
r65 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.825 $Y=0.755
+ $X2=9.825 $Y2=1.175
r66 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=9.3 $Y=1.475 $X2=9.3
+ $Y2=1.34
r67 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=9.3 $Y=1.475 $X2=9.3
+ $Y2=2.075
r68 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=1.485 $X2=10.055 $Y2=1.63
r69 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=1.485 $X2=10.055 $Y2=2.31
r70 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=9.93
+ $Y=0.235 $X2=10.055 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_1840_793# 1 2 9 12 13 15 26
r56 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=9.605 $Y=4.1
+ $X2=9.3 $Y2=4.1
r57 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=9.605 $Y=4.035
+ $X2=9.825 $Y2=4.035
r58 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.605
+ $Y=4.1 $X2=9.605 $Y2=4.1
r59 13 20 9.67586 $w=2.9e-07 $l=3.25269e-07 $layer=LI1_cond $X=10.055 $Y=3.805
+ $X2=9.825 $Y2=4.035
r60 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.055 $Y=3.805
+ $X2=10.055 $Y2=3.13
r61 12 25 8.93631 $w=3.14e-07 $l=3.18842e-07 $layer=LI1_cond $X=9.825 $Y=4.685
+ $X2=10.055 $Y2=4.897
r62 11 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=9.825 $Y=4.265
+ $X2=9.825 $Y2=4.035
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.825 $Y=4.265
+ $X2=9.825 $Y2=4.685
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=9.3 $Y=3.965 $X2=9.3
+ $Y2=4.1
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=9.3 $Y=3.965 $X2=9.3
+ $Y2=3.365
r66 2 13 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=2.955 $X2=10.055 $Y2=3.81
r67 2 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=2.955 $X2=10.055 $Y2=3.13
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=9.93
+ $Y=4.685 $X2=10.055 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[4] 1 3 4 5 6 8 9 11 12 17
r49 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.255
+ $Y=1.03 $X2=10.255 $Y2=1.03
r50 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=10.255 $Y=0.905
+ $X2=10.255 $Y2=1.03
r51 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=10.285 $Y=1.19
+ $X2=10.285 $Y2=1.03
r52 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=10.29 $Y=0.83
+ $X2=10.255 $Y2=0.905
r53 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.29 $Y=0.83
+ $X2=10.29 $Y2=0.495
r54 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=10.29 $Y=1.41
+ $X2=10.255 $Y2=1.03
r55 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.29 $Y=1.41
+ $X2=10.29 $Y2=1.985
r56 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.12 $Y=0.905
+ $X2=10.255 $Y2=0.905
r57 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=10.12 $Y=0.905 $X2=9.3
+ $Y2=0.905
r58 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.225 $Y=0.83
+ $X2=9.3 $Y2=0.905
r59 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.225 $Y=0.83
+ $X2=9.225 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[12] 1 3 4 5 6 8 9 11 12
r48 15 17 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=10.255 $Y=4.41
+ $X2=10.255 $Y2=4.535
r49 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.255
+ $Y=4.41 $X2=10.255 $Y2=4.41
r50 12 16 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=10.285 $Y=4.25
+ $X2=10.285 $Y2=4.41
r51 9 17 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=10.29 $Y=4.61
+ $X2=10.255 $Y2=4.535
r52 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.29 $Y=4.61
+ $X2=10.29 $Y2=4.945
r53 6 15 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=10.29 $Y=4.03
+ $X2=10.255 $Y2=4.41
r54 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.29 $Y=4.03
+ $X2=10.29 $Y2=3.455
r55 4 17 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.12 $Y=4.535
+ $X2=10.255 $Y2=4.535
r56 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=10.12 $Y=4.535 $X2=9.3
+ $Y2=4.535
r57 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.225 $Y=4.61
+ $X2=9.3 $Y2=4.535
r58 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.225 $Y=4.61
+ $X2=9.225 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[5] 1 3 4 6 7 9 11 12 17
r46 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.905
+ $Y=1.03 $X2=10.905 $Y2=1.03
r47 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=10.905 $Y=0.905
+ $X2=10.905 $Y2=1.03
r48 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=10.875 $Y=1.19
+ $X2=10.875 $Y2=1.03
r49 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=11.935 $Y=0.83
+ $X2=11.935 $Y2=0.495
r50 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.04 $Y=0.905
+ $X2=10.905 $Y2=0.905
r51 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.86 $Y=0.905
+ $X2=11.935 $Y2=0.83
r52 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=11.86 $Y=0.905
+ $X2=11.04 $Y2=0.905
r53 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=10.87 $Y=0.83
+ $X2=10.905 $Y2=0.905
r54 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.87 $Y=0.83
+ $X2=10.87 $Y2=0.495
r55 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=10.87 $Y=1.41
+ $X2=10.905 $Y2=1.03
r56 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.87 $Y=1.41
+ $X2=10.87 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[13] 1 3 4 6 7 9 11 12
r47 15 17 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=10.905 $Y=4.41
+ $X2=10.905 $Y2=4.535
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.905
+ $Y=4.41 $X2=10.905 $Y2=4.41
r49 12 16 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=10.875 $Y=4.25
+ $X2=10.875 $Y2=4.41
r50 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=11.935 $Y=4.61
+ $X2=11.935 $Y2=4.945
r51 8 17 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.04 $Y=4.535
+ $X2=10.905 $Y2=4.535
r52 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.86 $Y=4.535
+ $X2=11.935 $Y2=4.61
r53 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=11.86 $Y=4.535
+ $X2=11.04 $Y2=4.535
r54 4 17 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=10.87 $Y=4.61
+ $X2=10.905 $Y2=4.535
r55 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.87 $Y=4.61
+ $X2=10.87 $Y2=4.945
r56 1 15 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=10.87 $Y=4.03
+ $X2=10.905 $Y2=4.41
r57 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.87 $Y=4.03
+ $X2=10.87 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2189_47# 1 2 9 13 16 19 22 24
r57 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=11.555 $Y=1.34
+ $X2=11.86 $Y2=1.34
r58 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.555
+ $Y=1.34 $X2=11.555 $Y2=1.34
r59 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=11.335 $Y=1.405
+ $X2=11.555 $Y2=1.405
r60 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=11.105 $Y=1.63
+ $X2=11.335 $Y2=1.405
r61 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=11.335 $Y=1.175
+ $X2=11.335 $Y2=1.405
r62 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=11.335 $Y=0.755
+ $X2=11.105 $Y2=0.542
r63 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=11.335 $Y=0.755
+ $X2=11.335 $Y2=1.175
r64 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=11.105 $Y=2.31
+ $X2=11.105 $Y2=1.635
r65 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.86 $Y=1.475
+ $X2=11.86 $Y2=1.34
r66 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=11.86 $Y=1.475 $X2=11.86
+ $Y2=2.075
r67 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.96
+ $Y=1.485 $X2=11.105 $Y2=1.63
r68 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.96
+ $Y=1.485 $X2=11.105 $Y2=2.31
r69 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=10.945
+ $Y=0.235 $X2=11.105 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2189_937# 1 2 9 13 16 19 22 24
r59 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=11.555 $Y=4.1
+ $X2=11.86 $Y2=4.1
r60 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.555
+ $Y=4.1 $X2=11.555 $Y2=4.1
r61 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=11.335 $Y=4.035
+ $X2=11.555 $Y2=4.035
r62 16 24 8.93631 $w=3.14e-07 $l=3.18842e-07 $layer=LI1_cond $X=11.335 $Y=4.685
+ $X2=11.105 $Y2=4.897
r63 15 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=11.335 $Y=4.265
+ $X2=11.335 $Y2=4.035
r64 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=11.335 $Y=4.265
+ $X2=11.335 $Y2=4.685
r65 11 19 9.67586 $w=2.9e-07 $l=3.25269e-07 $layer=LI1_cond $X=11.105 $Y=3.805
+ $X2=11.335 $Y2=4.035
r66 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=11.105 $Y=3.805
+ $X2=11.105 $Y2=3.13
r67 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.86 $Y=3.965
+ $X2=11.86 $Y2=4.1
r68 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=11.86 $Y=3.965 $X2=11.86
+ $Y2=3.365
r69 2 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.96
+ $Y=2.955 $X2=11.105 $Y2=3.81
r70 2 13 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.96
+ $Y=2.955 $X2=11.105 $Y2=3.13
r71 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=10.945
+ $Y=4.685 $X2=11.105 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[5] 1 3 4 6 8 12 15 21
c38 8 0 1.78369e-19 $X=12.235 $Y=1.055
c39 1 0 2.31671e-19 $X=12.385 $Y=1.41
r40 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=12.19 $Y=0.51
+ $X2=12.235 $Y2=0.51
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.38
+ $Y=1.16 $X2=12.38 $Y2=1.16
r42 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=12.235 $Y=1.19
+ $X2=12.38 $Y2=1.19
r43 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.235 $Y=1.055
+ $X2=12.235 $Y2=1.19
r44 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=12.235 $Y=0.625
+ $X2=12.235 $Y2=0.51
r45 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=12.235 $Y=0.625
+ $X2=12.235 $Y2=1.055
r46 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=12.41 $Y=0.995
+ $X2=12.38 $Y2=1.16
r47 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.41 $Y=0.995
+ $X2=12.41 $Y2=0.56
r48 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=12.385 $Y=1.41
+ $X2=12.38 $Y2=1.16
r49 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.385 $Y=1.41
+ $X2=12.385 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[13] 1 3 4 6 8 12 15 21
c41 8 0 1.78369e-19 $X=12.235 $Y=4.815
c42 4 0 2.31671e-19 $X=12.41 $Y=4.445
r43 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=12.19 $Y=4.93
+ $X2=12.235 $Y2=4.93
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.38
+ $Y=4.28 $X2=12.38 $Y2=4.28
r45 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=12.235 $Y=4.25
+ $X2=12.38 $Y2=4.25
r46 8 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=12.235 $Y=4.815
+ $X2=12.235 $Y2=4.93
r47 7 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.235 $Y=4.385
+ $X2=12.235 $Y2=4.25
r48 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=12.235 $Y=4.385
+ $X2=12.235 $Y2=4.815
r49 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=12.41 $Y=4.445
+ $X2=12.38 $Y2=4.28
r50 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.41 $Y=4.445
+ $X2=12.41 $Y2=4.88
r51 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=12.385 $Y=4.03
+ $X2=12.38 $Y2=4.28
r52 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.385 $Y=4.03
+ $X2=12.385 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[6] 1 3 4 6 8 13 15
c38 8 0 1.78369e-19 $X=13.065 $Y=1.055
c39 4 0 2.31671e-19 $X=12.915 $Y=1.41
r40 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=13.11 $Y=0.51
+ $X2=13.065 $Y2=0.51
r41 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=12.92 $Y=1.19
+ $X2=13.065 $Y2=1.19
r42 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.92
+ $Y=1.16 $X2=12.92 $Y2=1.16
r43 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.065 $Y=1.055
+ $X2=13.065 $Y2=1.19
r44 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=13.065 $Y=0.625
+ $X2=13.065 $Y2=0.51
r45 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.065 $Y=0.625
+ $X2=13.065 $Y2=1.055
r46 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=12.915 $Y=1.41
+ $X2=12.92 $Y2=1.16
r47 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.915 $Y=1.41
+ $X2=12.915 $Y2=1.985
r48 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=12.89 $Y=0.995
+ $X2=12.92 $Y2=1.16
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.89 $Y=0.995
+ $X2=12.89 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[14] 1 3 4 6 8 13 15
c41 8 0 1.78369e-19 $X=13.065 $Y=4.815
c42 1 0 2.31671e-19 $X=12.89 $Y=4.445
r43 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=13.11 $Y=4.93
+ $X2=13.065 $Y2=4.93
r44 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=12.92 $Y=4.25
+ $X2=13.065 $Y2=4.25
r45 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.92
+ $Y=4.28 $X2=12.92 $Y2=4.28
r46 8 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=13.065 $Y=4.815
+ $X2=13.065 $Y2=4.93
r47 7 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.065 $Y=4.385
+ $X2=13.065 $Y2=4.25
r48 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.065 $Y=4.385
+ $X2=13.065 $Y2=4.815
r49 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=12.915 $Y=4.03
+ $X2=12.92 $Y2=4.28
r50 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.915 $Y=4.03
+ $X2=12.915 $Y2=3.455
r51 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=12.89 $Y=4.445
+ $X2=12.92 $Y2=4.28
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.89 $Y=4.445
+ $X2=12.89 $Y2=4.88
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2668_265# 1 2 9 11 12 15 22 26
r58 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=13.965 $Y=1.405
+ $X2=14.195 $Y2=1.63
r59 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=13.745 $Y=1.34
+ $X2=13.44 $Y2=1.34
r60 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=13.745 $Y=1.405
+ $X2=13.965 $Y2=1.405
r61 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.745
+ $Y=1.34 $X2=13.745 $Y2=1.34
r62 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=14.195 $Y=2.31
+ $X2=14.195 $Y2=1.635
r63 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=13.965 $Y=1.175
+ $X2=13.965 $Y2=1.405
r64 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=13.965 $Y=0.755
+ $X2=14.195 $Y2=0.542
r65 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=13.965 $Y=0.755
+ $X2=13.965 $Y2=1.175
r66 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.44 $Y=1.475
+ $X2=13.44 $Y2=1.34
r67 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=13.44 $Y=1.475 $X2=13.44
+ $Y2=2.075
r68 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=14.07
+ $Y=1.485 $X2=14.195 $Y2=1.63
r69 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=14.07
+ $Y=1.485 $X2=14.195 $Y2=2.31
r70 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=14.07
+ $Y=0.235 $X2=14.195 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_2668_793# 1 2 9 12 13 15 26
r56 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=13.745 $Y=4.1
+ $X2=13.44 $Y2=4.1
r57 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=13.745 $Y=4.035
+ $X2=13.965 $Y2=4.035
r58 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.745
+ $Y=4.1 $X2=13.745 $Y2=4.1
r59 13 20 9.67586 $w=2.9e-07 $l=3.25269e-07 $layer=LI1_cond $X=14.195 $Y=3.805
+ $X2=13.965 $Y2=4.035
r60 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=14.195 $Y=3.805
+ $X2=14.195 $Y2=3.13
r61 12 25 8.93631 $w=3.14e-07 $l=3.18842e-07 $layer=LI1_cond $X=13.965 $Y=4.685
+ $X2=14.195 $Y2=4.897
r62 11 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=13.965 $Y=4.265
+ $X2=13.965 $Y2=4.035
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=13.965 $Y=4.265
+ $X2=13.965 $Y2=4.685
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.44 $Y=3.965
+ $X2=13.44 $Y2=4.1
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=13.44 $Y=3.965 $X2=13.44
+ $Y2=3.365
r66 2 13 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=14.07
+ $Y=2.955 $X2=14.195 $Y2=3.81
r67 2 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=14.07
+ $Y=2.955 $X2=14.195 $Y2=3.13
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=14.07
+ $Y=4.685 $X2=14.195 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[6] 1 3 4 5 6 8 9 11 12 17
r49 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.395
+ $Y=1.03 $X2=14.395 $Y2=1.03
r50 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=14.395 $Y=0.905
+ $X2=14.395 $Y2=1.03
r51 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=14.425 $Y=1.19
+ $X2=14.425 $Y2=1.03
r52 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=14.43 $Y=0.83
+ $X2=14.395 $Y2=0.905
r53 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=14.43 $Y=0.83
+ $X2=14.43 $Y2=0.495
r54 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=14.43 $Y=1.41
+ $X2=14.395 $Y2=1.03
r55 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.43 $Y=1.41
+ $X2=14.43 $Y2=1.985
r56 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.26 $Y=0.905
+ $X2=14.395 $Y2=0.905
r57 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=14.26 $Y=0.905
+ $X2=13.44 $Y2=0.905
r58 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.365 $Y=0.83
+ $X2=13.44 $Y2=0.905
r59 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=13.365 $Y=0.83
+ $X2=13.365 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[14] 1 3 4 5 6 8 9 11 12
r48 15 17 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=14.395 $Y=4.41
+ $X2=14.395 $Y2=4.535
r49 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.395
+ $Y=4.41 $X2=14.395 $Y2=4.41
r50 12 16 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=14.425 $Y=4.25
+ $X2=14.425 $Y2=4.41
r51 9 17 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=14.43 $Y=4.61
+ $X2=14.395 $Y2=4.535
r52 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=14.43 $Y=4.61
+ $X2=14.43 $Y2=4.945
r53 6 15 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=14.43 $Y=4.03
+ $X2=14.395 $Y2=4.41
r54 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.43 $Y=4.03
+ $X2=14.43 $Y2=3.455
r55 4 17 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.26 $Y=4.535
+ $X2=14.395 $Y2=4.535
r56 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=14.26 $Y=4.535
+ $X2=13.44 $Y2=4.535
r57 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.365 $Y=4.61
+ $X2=13.44 $Y2=4.535
r58 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=13.365 $Y=4.61
+ $X2=13.365 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[7] 1 3 4 6 7 9 11 12 17
r46 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.045
+ $Y=1.03 $X2=15.045 $Y2=1.03
r47 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=15.045 $Y=0.905
+ $X2=15.045 $Y2=1.03
r48 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=15.015 $Y=1.19
+ $X2=15.015 $Y2=1.03
r49 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.075 $Y=0.83
+ $X2=16.075 $Y2=0.495
r50 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=15.18 $Y=0.905
+ $X2=15.045 $Y2=0.905
r51 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16 $Y=0.905
+ $X2=16.075 $Y2=0.83
r52 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=16 $Y=0.905 $X2=15.18
+ $Y2=0.905
r53 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=15.01 $Y=0.83
+ $X2=15.045 $Y2=0.905
r54 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.01 $Y=0.83
+ $X2=15.01 $Y2=0.495
r55 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=15.01 $Y=1.41
+ $X2=15.045 $Y2=1.03
r56 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.01 $Y=1.41
+ $X2=15.01 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%S[15] 1 3 4 6 7 9 11 12
r47 15 17 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=15.045 $Y=4.41
+ $X2=15.045 $Y2=4.535
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.045
+ $Y=4.41 $X2=15.045 $Y2=4.41
r49 12 16 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=15.015 $Y=4.25
+ $X2=15.015 $Y2=4.41
r50 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.075 $Y=4.61
+ $X2=16.075 $Y2=4.945
r51 8 17 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=15.18 $Y=4.535
+ $X2=15.045 $Y2=4.535
r52 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16 $Y=4.535
+ $X2=16.075 $Y2=4.61
r53 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=16 $Y=4.535 $X2=15.18
+ $Y2=4.535
r54 4 17 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=15.01 $Y=4.61
+ $X2=15.045 $Y2=4.535
r55 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.01 $Y=4.61
+ $X2=15.01 $Y2=4.945
r56 1 15 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=15.01 $Y=4.03
+ $X2=15.045 $Y2=4.41
r57 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.01 $Y=4.03
+ $X2=15.01 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_3017_47# 1 2 9 13 16 19 22 24
r57 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=15.695 $Y=1.34
+ $X2=16 $Y2=1.34
r58 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.695
+ $Y=1.34 $X2=15.695 $Y2=1.34
r59 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=15.475 $Y=1.405
+ $X2=15.695 $Y2=1.405
r60 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=15.245 $Y=1.63
+ $X2=15.475 $Y2=1.405
r61 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=15.475 $Y=1.175
+ $X2=15.475 $Y2=1.405
r62 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=15.475 $Y=0.755
+ $X2=15.245 $Y2=0.542
r63 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=15.475 $Y=0.755
+ $X2=15.475 $Y2=1.175
r64 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=15.245 $Y=2.31
+ $X2=15.245 $Y2=1.635
r65 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=16 $Y=1.475 $X2=16
+ $Y2=1.34
r66 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=16 $Y=1.475 $X2=16
+ $Y2=2.075
r67 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=15.1
+ $Y=1.485 $X2=15.245 $Y2=1.63
r68 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=15.1
+ $Y=1.485 $X2=15.245 $Y2=2.31
r69 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=15.085
+ $Y=0.235 $X2=15.245 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%A_3017_937# 1 2 9 13 16 19 22 24
r59 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=15.695 $Y=4.1
+ $X2=16 $Y2=4.1
r60 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.695
+ $Y=4.1 $X2=15.695 $Y2=4.1
r61 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=15.475 $Y=4.035
+ $X2=15.695 $Y2=4.035
r62 16 24 8.93631 $w=3.14e-07 $l=3.18842e-07 $layer=LI1_cond $X=15.475 $Y=4.685
+ $X2=15.245 $Y2=4.897
r63 15 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=15.475 $Y=4.265
+ $X2=15.475 $Y2=4.035
r64 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=15.475 $Y=4.265
+ $X2=15.475 $Y2=4.685
r65 11 19 9.67586 $w=2.9e-07 $l=3.25269e-07 $layer=LI1_cond $X=15.245 $Y=3.805
+ $X2=15.475 $Y2=4.035
r66 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=15.245 $Y=3.805
+ $X2=15.245 $Y2=3.13
r67 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=16 $Y=3.965 $X2=16
+ $Y2=4.1
r68 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=16 $Y=3.965 $X2=16
+ $Y2=3.365
r69 2 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=15.1
+ $Y=2.955 $X2=15.245 $Y2=3.81
r70 2 13 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=15.1
+ $Y=2.955 $X2=15.245 $Y2=3.13
r71 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=15.085
+ $Y=4.685 $X2=15.245 $Y2=4.945
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[7] 1 3 4 6 8 12 15 21
c29 1 0 5.33021e-20 $X=16.525 $Y=1.41
r30 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=16.33 $Y=0.51
+ $X2=16.375 $Y2=0.51
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.52
+ $Y=1.16 $X2=16.52 $Y2=1.16
r32 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=16.375 $Y=1.19
+ $X2=16.52 $Y2=1.19
r33 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.375 $Y=1.055
+ $X2=16.375 $Y2=1.19
r34 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=16.375 $Y=0.625
+ $X2=16.375 $Y2=0.51
r35 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=16.375 $Y=0.625
+ $X2=16.375 $Y2=1.055
r36 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=16.55 $Y=0.995
+ $X2=16.52 $Y2=1.16
r37 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=16.55 $Y=0.995
+ $X2=16.55 $Y2=0.56
r38 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=16.525 $Y=1.41
+ $X2=16.52 $Y2=1.16
r39 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.525 $Y=1.41
+ $X2=16.525 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%D[15] 1 3 4 6 8 12 15 21
c31 4 0 5.33021e-20 $X=16.55 $Y=4.445
r32 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=16.33 $Y=4.93
+ $X2=16.375 $Y2=4.93
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.52
+ $Y=4.28 $X2=16.52 $Y2=4.28
r34 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=16.375 $Y=4.25
+ $X2=16.52 $Y2=4.25
r35 8 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=16.375 $Y=4.815
+ $X2=16.375 $Y2=4.93
r36 7 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.375 $Y=4.385
+ $X2=16.375 $Y2=4.25
r37 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=16.375 $Y=4.385
+ $X2=16.375 $Y2=4.815
r38 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=16.55 $Y=4.445
+ $X2=16.52 $Y2=4.28
r39 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=16.55 $Y=4.445
+ $X2=16.55 $Y2=4.88
r40 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=16.525 $Y=4.03
+ $X2=16.52 $Y2=4.28
r41 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.525 $Y=4.03
+ $X2=16.525 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 57 63 69 75 81 87 93 99 105 111 117 123 129 135 141 147 153 159
+ 164 165 167 168 170 171 173 174 175 176 177 178 179 187 195 198 205 213 216
+ 223 231 234 241 249 252 258 270
r491 254 255 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.33 $Y=2.72
+ $X2=16.33 $Y2=2.72
r492 252 270 3.80956 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=16.595 $Y=2.72
+ $X2=16.807 $Y2=2.72
r493 252 254 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=16.595 $Y=2.72
+ $X2=16.33 $Y2=2.72
r494 250 255 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=16.33 $Y2=2.72
r495 249 250 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.41 $Y=2.72
+ $X2=15.41 $Y2=2.72
r496 246 250 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=15.41 $Y2=2.72
r497 245 246 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=2.72
+ $X2=14.49 $Y2=2.72
r498 242 246 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=14.49 $Y2=2.72
r499 241 242 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r500 239 267 13.9941 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.845 $Y=2.72
+ $X2=12.65 $Y2=2.72
r501 239 241 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=12.845 $Y=2.72
+ $X2=13.11 $Y2=2.72
r502 236 237 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r503 234 267 13.9941 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.455 $Y=2.72
+ $X2=12.65 $Y2=2.72
r504 234 236 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=12.455 $Y=2.72
+ $X2=12.19 $Y2=2.72
r505 232 237 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=12.19 $Y2=2.72
r506 231 232 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r507 228 232 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r508 227 228 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r509 224 228 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=10.35 $Y2=2.72
r510 223 224 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r511 221 264 13.9941 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=8.705 $Y=2.72
+ $X2=8.51 $Y2=2.72
r512 221 223 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.705 $Y=2.72
+ $X2=8.97 $Y2=2.72
r513 218 219 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r514 216 264 13.9941 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=8.315 $Y=2.72
+ $X2=8.51 $Y2=2.72
r515 216 218 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.315 $Y=2.72
+ $X2=8.05 $Y2=2.72
r516 214 219 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r517 213 214 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r518 210 214 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r519 209 210 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r520 206 210 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=6.21 $Y2=2.72
r521 205 206 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r522 203 261 13.9941 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.37 $Y2=2.72
r523 203 205 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.83 $Y2=2.72
r524 200 201 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r525 198 261 13.9941 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.175 $Y=2.72
+ $X2=4.37 $Y2=2.72
r526 198 200 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.175 $Y=2.72
+ $X2=3.91 $Y2=2.72
r527 196 201 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r528 195 196 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r529 192 196 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r530 191 192 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r531 188 192 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r532 187 188 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r533 185 258 3.80956 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r534 185 187 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r535 179 255 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=16.79 $Y=2.72
+ $X2=16.33 $Y2=2.72
r536 179 270 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.79 $Y=2.72
+ $X2=16.79 $Y2=2.72
r537 178 242 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r538 178 237 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r539 178 267 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r540 177 224 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r541 177 219 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r542 177 264 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r543 176 206 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r544 176 201 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r545 176 261 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r546 175 188 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r547 175 258 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r548 173 245 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.555 $Y=2.72
+ $X2=14.49 $Y2=2.72
r549 173 174 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.555 $Y=2.72
+ $X2=14.72 $Y2=2.72
r550 172 249 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=14.885 $Y=2.72
+ $X2=15.41 $Y2=2.72
r551 172 174 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.885 $Y=2.72
+ $X2=14.72 $Y2=2.72
r552 170 227 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.35 $Y2=2.72
r553 170 171 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.58 $Y2=2.72
r554 169 231 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=10.745 $Y=2.72
+ $X2=11.27 $Y2=2.72
r555 169 171 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.745 $Y=2.72
+ $X2=10.58 $Y2=2.72
r556 167 209 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.275 $Y=2.72
+ $X2=6.21 $Y2=2.72
r557 167 168 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=2.72
+ $X2=6.44 $Y2=2.72
r558 166 213 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=7.13 $Y2=2.72
r559 166 168 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=6.44 $Y2=2.72
r560 164 191 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.07 $Y2=2.72
r561 164 165 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.3 $Y2=2.72
r562 163 195 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.99 $Y2=2.72
r563 163 165 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.3 $Y2=2.72
r564 159 161 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=16.76 $Y=3.1
+ $X2=16.76 $Y2=3.78
r565 157 270 2.88756 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=16.76 $Y=2.805
+ $X2=16.807 $Y2=2.72
r566 157 159 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=16.76 $Y=2.805
+ $X2=16.76 $Y2=3.1
r567 153 156 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=16.76 $Y=1.66
+ $X2=16.76 $Y2=2.34
r568 151 270 2.88756 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=16.76 $Y=2.635
+ $X2=16.807 $Y2=2.72
r569 151 156 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=16.76 $Y=2.635
+ $X2=16.76 $Y2=2.34
r570 147 149 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=14.72 $Y=3.13
+ $X2=14.72 $Y2=3.81
r571 145 174 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.72 $Y=2.805
+ $X2=14.72 $Y2=2.72
r572 145 147 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=14.72 $Y=2.805
+ $X2=14.72 $Y2=3.13
r573 141 144 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=14.72 $Y=1.63
+ $X2=14.72 $Y2=2.31
r574 139 174 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.72 $Y=2.635
+ $X2=14.72 $Y2=2.72
r575 139 144 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=14.72 $Y=2.635
+ $X2=14.72 $Y2=2.31
r576 135 137 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=12.65 $Y=3.1
+ $X2=12.65 $Y2=3.78
r577 133 267 2.65897 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.65 $Y=2.805
+ $X2=12.65 $Y2=2.72
r578 133 135 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=12.65 $Y=2.805
+ $X2=12.65 $Y2=3.1
r579 129 132 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=12.65 $Y=1.66
+ $X2=12.65 $Y2=2.34
r580 127 267 2.65897 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.65 $Y=2.635
+ $X2=12.65 $Y2=2.72
r581 127 132 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=12.65 $Y=2.635
+ $X2=12.65 $Y2=2.34
r582 123 125 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.58 $Y=3.13
+ $X2=10.58 $Y2=3.81
r583 121 171 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.58 $Y=2.805
+ $X2=10.58 $Y2=2.72
r584 121 123 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=10.58 $Y=2.805
+ $X2=10.58 $Y2=3.13
r585 117 120 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.58 $Y=1.63
+ $X2=10.58 $Y2=2.31
r586 115 171 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.58 $Y=2.635
+ $X2=10.58 $Y2=2.72
r587 115 120 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=10.58 $Y=2.635
+ $X2=10.58 $Y2=2.31
r588 111 113 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=8.51 $Y=3.1
+ $X2=8.51 $Y2=3.78
r589 109 264 2.65897 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.51 $Y=2.805
+ $X2=8.51 $Y2=2.72
r590 109 111 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=8.51 $Y=2.805
+ $X2=8.51 $Y2=3.1
r591 105 108 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=8.51 $Y=1.66
+ $X2=8.51 $Y2=2.34
r592 103 264 2.65897 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.51 $Y=2.635
+ $X2=8.51 $Y2=2.72
r593 103 108 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=8.51 $Y=2.635
+ $X2=8.51 $Y2=2.34
r594 99 101 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.44 $Y=3.13
+ $X2=6.44 $Y2=3.81
r595 97 168 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=2.805
+ $X2=6.44 $Y2=2.72
r596 97 99 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.44 $Y=2.805
+ $X2=6.44 $Y2=3.13
r597 93 96 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.44 $Y=1.63
+ $X2=6.44 $Y2=2.31
r598 91 168 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=2.635
+ $X2=6.44 $Y2=2.72
r599 91 96 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.44 $Y=2.635
+ $X2=6.44 $Y2=2.31
r600 87 89 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=4.37 $Y=3.1
+ $X2=4.37 $Y2=3.78
r601 85 261 2.65897 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=2.805
+ $X2=4.37 $Y2=2.72
r602 85 87 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=4.37 $Y=2.805
+ $X2=4.37 $Y2=3.1
r603 81 84 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=4.37 $Y=1.66
+ $X2=4.37 $Y2=2.34
r604 79 261 2.65897 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=2.635
+ $X2=4.37 $Y2=2.72
r605 79 84 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=4.37 $Y=2.635
+ $X2=4.37 $Y2=2.34
r606 75 77 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.3 $Y=3.13 $X2=2.3
+ $Y2=3.81
r607 73 165 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.805
+ $X2=2.3 $Y2=2.72
r608 73 75 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.3 $Y=2.805
+ $X2=2.3 $Y2=3.13
r609 69 72 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.3 $Y=1.63 $X2=2.3
+ $Y2=2.31
r610 67 165 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.635
+ $X2=2.3 $Y2=2.72
r611 67 72 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.3 $Y=2.635
+ $X2=2.3 $Y2=2.31
r612 63 65 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.1
+ $X2=0.26 $Y2=3.78
r613 61 258 2.88756 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.805
+ $X2=0.212 $Y2=2.72
r614 61 63 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.805
+ $X2=0.26 $Y2=3.1
r615 57 60 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r616 55 258 2.88756 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r617 55 60 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r618 18 161 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=16.615
+ $Y=2.955 $X2=16.76 $Y2=3.78
r619 18 159 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=16.615
+ $Y=2.955 $X2=16.76 $Y2=3.1
r620 17 156 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=16.615
+ $Y=1.485 $X2=16.76 $Y2=2.34
r621 17 153 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=16.615
+ $Y=1.485 $X2=16.76 $Y2=1.66
r622 16 149 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=2.955 $X2=14.72 $Y2=3.81
r623 16 147 400 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=2.955 $X2=14.72 $Y2=3.13
r624 15 144 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=1.485 $X2=14.72 $Y2=2.31
r625 15 141 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=1.485 $X2=14.72 $Y2=1.63
r626 14 137 400 $w=1.7e-07 $l=9.08295e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=2.955 $X2=12.65 $Y2=3.78
r627 14 135 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=2.955 $X2=12.65 $Y2=3.1
r628 13 132 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.65 $Y2=2.34
r629 13 129 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.65 $Y2=1.66
r630 12 125 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=10.38
+ $Y=2.955 $X2=10.58 $Y2=3.81
r631 12 123 400 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=10.38
+ $Y=2.955 $X2=10.58 $Y2=3.13
r632 11 120 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=10.38
+ $Y=1.485 $X2=10.58 $Y2=2.31
r633 11 117 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=10.38
+ $Y=1.485 $X2=10.58 $Y2=1.63
r634 10 113 400 $w=1.7e-07 $l=9.08295e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=2.955 $X2=8.51 $Y2=3.78
r635 10 111 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=2.955 $X2=8.51 $Y2=3.1
r636 9 108 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=1.485 $X2=8.51 $Y2=2.34
r637 9 105 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=1.485 $X2=8.51 $Y2=1.66
r638 8 101 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=2.955 $X2=6.44 $Y2=3.81
r639 8 99 400 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=2.955 $X2=6.44 $Y2=3.13
r640 7 96 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.485 $X2=6.44 $Y2=2.31
r641 7 93 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.485 $X2=6.44 $Y2=1.63
r642 6 89 400 $w=1.7e-07 $l=9.08295e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=2.955 $X2=4.37 $Y2=3.78
r643 6 87 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=2.955 $X2=4.37 $Y2=3.1
r644 5 84 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.485 $X2=4.37 $Y2=2.34
r645 5 81 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.485 $X2=4.37 $Y2=1.66
r646 4 77 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=2.955 $X2=2.3 $Y2=3.81
r647 4 75 400 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=2.955 $X2=2.3 $Y2=3.13
r648 3 72 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.485 $X2=2.3 $Y2=2.31
r649 3 69 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.485 $X2=2.3 $Y2=1.63
r650 2 65 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.955 $X2=0.26 $Y2=3.78
r651 2 63 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.955 $X2=0.26 $Y2=3.1
r652 1 60 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r653 1 57 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%Z 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 98 100 101 103 105 107 112
+ 116 120 122 127 131 134 136 138 140 141 143 145 147 152 156 160 162 167 171
+ 174 176 178 180 181 183 185 187 192 196 200 202 207 211 214 216 218 220 221
+ 223 225 227 232 236 240 242 247 251 254 256 265 267 268 269 271 272 275 279
+ 289 291 292 293 295 296 299 303 313 315 316 317 319 320 323 327 337 339 340
+ 341 343 344 347 351 353 354 355 356 357 358 359 360 361 362 363 364 365 366
+ 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385
+ 386 387 388 389 390 391 392 393 394 395 396 415 420 425 430 435 440 445 450
+ 455 460 465 470 475 480 485 490
c1026 351 0 5.33021e-20 $X=16.035 $Y=4.52
c1027 347 0 5.33021e-20 $X=16.035 $Y=0.92
c1028 327 0 5.33021e-20 $X=11.895 $Y=4.52
c1029 323 0 5.33021e-20 $X=11.895 $Y=0.92
c1030 303 0 5.33021e-20 $X=7.755 $Y=4.52
c1031 299 0 5.33021e-20 $X=7.755 $Y=0.92
c1032 279 0 5.33021e-20 $X=3.615 $Y=4.52
c1033 275 0 5.33021e-20 $X=3.615 $Y=0.92
c1034 225 0 5.33021e-20 $X=13.587 $Y=4.605
c1035 221 0 5.33021e-20 $X=13.587 $Y=0.835
c1036 185 0 5.33021e-20 $X=9.447 $Y=4.605
c1037 181 0 5.33021e-20 $X=9.447 $Y=0.835
c1038 145 0 5.33021e-20 $X=5.307 $Y=4.605
c1039 141 0 5.33021e-20 $X=5.307 $Y=0.835
c1040 105 0 5.33021e-20 $X=1.167 $Y=4.605
c1041 101 0 5.33021e-20 $X=1.167 $Y=0.835
r1042 490 492 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=15.87 $Y=3.57
+ $X2=16.035 $Y2=3.57
r1043 485 487 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=15.87 $Y=1.87
+ $X2=16.035 $Y2=1.87
r1044 478 480 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=3.57
+ $X2=13.57 $Y2=3.57
r1045 473 475 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=1.87
+ $X2=13.57 $Y2=1.87
r1046 470 472 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=11.73 $Y=3.57
+ $X2=11.895 $Y2=3.57
r1047 465 467 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=11.73 $Y=1.87
+ $X2=11.895 $Y2=1.87
r1048 458 460 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=9.265 $Y=3.57
+ $X2=9.43 $Y2=3.57
r1049 453 455 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=9.265 $Y=1.87
+ $X2=9.43 $Y2=1.87
r1050 450 452 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=7.59 $Y=3.57
+ $X2=7.755 $Y2=3.57
r1051 445 447 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=7.59 $Y=1.87
+ $X2=7.755 $Y2=1.87
r1052 438 440 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=3.57
+ $X2=5.29 $Y2=3.57
r1053 433 435 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=1.87
+ $X2=5.29 $Y2=1.87
r1054 430 432 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=3.57
+ $X2=3.615 $Y2=3.57
r1055 425 427 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=1.87
+ $X2=3.615 $Y2=1.87
r1056 418 420 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.57
+ $X2=1.15 $Y2=3.57
r1057 413 415 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=1.87
+ $X2=1.15 $Y2=1.87
r1058 396 490 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.87 $Y=3.57
+ $X2=15.87 $Y2=3.57
r1059 395 485 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.87 $Y=1.87
+ $X2=15.87 $Y2=1.87
r1060 394 480 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=3.57
+ $X2=13.57 $Y2=3.57
r1061 393 475 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=1.87
+ $X2=13.57 $Y2=1.87
r1062 392 470 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=3.57
+ $X2=11.73 $Y2=3.57
r1063 391 465 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=1.87
+ $X2=11.73 $Y2=1.87
r1064 390 460 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=3.57
+ $X2=9.43 $Y2=3.57
r1065 389 455 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=1.87
+ $X2=9.43 $Y2=1.87
r1066 388 450 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=3.57
+ $X2=7.59 $Y2=3.57
r1067 387 445 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=1.87
+ $X2=7.59 $Y2=1.87
r1068 386 440 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=3.57
+ $X2=5.29 $Y2=3.57
r1069 385 435 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r1070 384 430 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=3.57
+ $X2=3.45 $Y2=3.57
r1071 383 425 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=1.87
+ $X2=3.45 $Y2=1.87
r1072 382 420 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=3.57
+ $X2=1.15 $Y2=3.57
r1073 381 415 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.87
+ $X2=1.15 $Y2=1.87
r1074 380 394 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.715 $Y=3.57
+ $X2=13.57 $Y2=3.57
r1075 379 396 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.725 $Y=3.57
+ $X2=15.87 $Y2=3.57
r1076 379 380 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=15.725 $Y=3.57
+ $X2=13.715 $Y2=3.57
r1077 378 393 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.715 $Y=1.87
+ $X2=13.57 $Y2=1.87
r1078 377 395 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.725 $Y=1.87
+ $X2=15.87 $Y2=1.87
r1079 377 378 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=15.725 $Y=1.87
+ $X2=13.715 $Y2=1.87
r1080 376 392 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.875 $Y=3.57
+ $X2=11.73 $Y2=3.57
r1081 375 394 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.425 $Y=3.57
+ $X2=13.57 $Y2=3.57
r1082 375 376 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=13.425 $Y=3.57
+ $X2=11.875 $Y2=3.57
r1083 374 391 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.875 $Y=1.87
+ $X2=11.73 $Y2=1.87
r1084 373 393 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.425 $Y=1.87
+ $X2=13.57 $Y2=1.87
r1085 373 374 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=13.425 $Y=1.87
+ $X2=11.875 $Y2=1.87
r1086 372 390 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.575 $Y=3.57
+ $X2=9.43 $Y2=3.57
r1087 371 392 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.585 $Y=3.57
+ $X2=11.73 $Y2=3.57
r1088 371 372 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=11.585 $Y=3.57
+ $X2=9.575 $Y2=3.57
r1089 370 389 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.575 $Y=1.87
+ $X2=9.43 $Y2=1.87
r1090 369 391 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.585 $Y=1.87
+ $X2=11.73 $Y2=1.87
r1091 369 370 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=11.585 $Y=1.87
+ $X2=9.575 $Y2=1.87
r1092 368 388 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.735 $Y=3.57
+ $X2=7.59 $Y2=3.57
r1093 367 390 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.285 $Y=3.57
+ $X2=9.43 $Y2=3.57
r1094 367 368 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=9.285 $Y=3.57
+ $X2=7.735 $Y2=3.57
r1095 366 387 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.735 $Y=1.87
+ $X2=7.59 $Y2=1.87
r1096 365 389 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.285 $Y=1.87
+ $X2=9.43 $Y2=1.87
r1097 365 366 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=9.285 $Y=1.87
+ $X2=7.735 $Y2=1.87
r1098 364 386 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=3.57
+ $X2=5.29 $Y2=3.57
r1099 363 388 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=3.57
+ $X2=7.59 $Y2=3.57
r1100 363 364 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=7.445 $Y=3.57
+ $X2=5.435 $Y2=3.57
r1101 362 385 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=1.87
+ $X2=5.29 $Y2=1.87
r1102 361 387 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=1.87
+ $X2=7.59 $Y2=1.87
r1103 361 362 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=7.445 $Y=1.87
+ $X2=5.435 $Y2=1.87
r1104 360 384 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.595 $Y=3.57
+ $X2=3.45 $Y2=3.57
r1105 359 386 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=3.57
+ $X2=5.29 $Y2=3.57
r1106 359 360 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=5.145 $Y=3.57
+ $X2=3.595 $Y2=3.57
r1107 358 383 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.595 $Y=1.87
+ $X2=3.45 $Y2=1.87
r1108 357 385 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r1109 357 358 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=3.595 $Y2=1.87
r1110 356 382 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=3.57
+ $X2=1.15 $Y2=3.57
r1111 355 384 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.305 $Y=3.57
+ $X2=3.45 $Y2=3.57
r1112 355 356 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=3.305 $Y=3.57
+ $X2=1.295 $Y2=3.57
r1113 354 381 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.87
+ $X2=1.15 $Y2=1.87
r1114 353 383 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.305 $Y=1.87
+ $X2=3.45 $Y2=1.87
r1115 353 354 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=3.305 $Y=1.87
+ $X2=1.295 $Y2=1.87
r1116 343 344 6.00906 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=15.765 $Y=3.1
+ $X2=15.765 $Y2=2.975
r1117 341 344 27.592 $w=2.03e-07 $l=5.1e-07 $layer=LI1_cond $X=15.827 $Y=2.465
+ $X2=15.827 $Y2=2.975
r1118 339 340 6.00906 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=13.675 $Y=3.1
+ $X2=13.675 $Y2=2.975
r1119 337 340 27.592 $w=2.03e-07 $l=5.1e-07 $layer=LI1_cond $X=13.612 $Y=2.465
+ $X2=13.612 $Y2=2.975
r1120 319 320 6.00906 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=11.625 $Y=3.1
+ $X2=11.625 $Y2=2.975
r1121 317 320 27.592 $w=2.03e-07 $l=5.1e-07 $layer=LI1_cond $X=11.687 $Y=2.465
+ $X2=11.687 $Y2=2.975
r1122 315 316 6.00906 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=9.535 $Y=3.1
+ $X2=9.535 $Y2=2.975
r1123 313 316 27.592 $w=2.03e-07 $l=5.1e-07 $layer=LI1_cond $X=9.472 $Y=2.465
+ $X2=9.472 $Y2=2.975
r1124 295 296 6.00906 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=7.485 $Y=3.1
+ $X2=7.485 $Y2=2.975
r1125 293 296 27.592 $w=2.03e-07 $l=5.1e-07 $layer=LI1_cond $X=7.547 $Y=2.465
+ $X2=7.547 $Y2=2.975
r1126 291 292 6.00906 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=5.395 $Y=3.1
+ $X2=5.395 $Y2=2.975
r1127 289 292 27.592 $w=2.03e-07 $l=5.1e-07 $layer=LI1_cond $X=5.332 $Y=2.465
+ $X2=5.332 $Y2=2.975
r1128 271 272 6.00906 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=3.1
+ $X2=3.345 $Y2=2.975
r1129 269 272 27.592 $w=2.03e-07 $l=5.1e-07 $layer=LI1_cond $X=3.407 $Y=2.465
+ $X2=3.407 $Y2=2.975
r1130 267 268 6.00906 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.255 $Y=3.1
+ $X2=1.255 $Y2=2.975
r1131 265 268 27.592 $w=2.03e-07 $l=5.1e-07 $layer=LI1_cond $X=1.192 $Y=2.465
+ $X2=1.192 $Y2=2.975
r1132 256 351 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.035 $Y=4.435
+ $X2=16.035 $Y2=4.52
r1133 255 492 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=16.035 $Y=3.685
+ $X2=16.035 $Y2=3.57
r1134 255 256 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=16.035 $Y=3.685
+ $X2=16.035 $Y2=4.435
r1135 254 487 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=16.035 $Y=1.755
+ $X2=16.035 $Y2=1.87
r1136 253 347 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.035 $Y=1.005
+ $X2=16.035 $Y2=0.92
r1137 253 254 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=16.035 $Y=1.005
+ $X2=16.035 $Y2=1.755
r1138 249 351 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=15.852 $Y=4.52
+ $X2=16.035 $Y2=4.52
r1139 249 251 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=15.852 $Y=4.605
+ $X2=15.852 $Y2=4.945
r1140 245 347 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=15.852 $Y=0.92
+ $X2=16.035 $Y2=0.92
r1141 245 247 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=15.852 $Y=0.835
+ $X2=15.852 $Y2=0.495
r1142 242 490 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=15.765 $Y=3.57
+ $X2=15.87 $Y2=3.57
r1143 241 343 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=15.765 $Y=3.14
+ $X2=15.765 $Y2=3.1
r1144 241 242 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=15.765 $Y=3.14
+ $X2=15.765 $Y2=3.455
r1145 238 341 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=15.765 $Y=2.3
+ $X2=15.765 $Y2=2.465
r1146 238 240 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=15.765 $Y=2.3
+ $X2=15.765 $Y2=2
r1147 237 485 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=15.765 $Y=1.87
+ $X2=15.87 $Y2=1.87
r1148 237 240 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=15.765 $Y=1.985
+ $X2=15.765 $Y2=2
r1149 236 480 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=13.675 $Y=3.57
+ $X2=13.57 $Y2=3.57
r1150 235 339 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=13.675 $Y=3.14
+ $X2=13.675 $Y2=3.1
r1151 235 236 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=13.675 $Y=3.14
+ $X2=13.675 $Y2=3.455
r1152 230 337 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.675 $Y=2.3
+ $X2=13.675 $Y2=2.465
r1153 230 232 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=13.675 $Y=2.3
+ $X2=13.675 $Y2=2
r1154 229 475 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=13.675 $Y=1.87
+ $X2=13.57 $Y2=1.87
r1155 229 232 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=13.675 $Y=1.985
+ $X2=13.675 $Y2=2
r1156 225 333 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=13.587 $Y=4.52
+ $X2=13.405 $Y2=4.52
r1157 225 227 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=13.587 $Y=4.605
+ $X2=13.587 $Y2=4.945
r1158 221 329 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=13.587 $Y=0.92
+ $X2=13.405 $Y2=0.92
r1159 221 223 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=13.587 $Y=0.835
+ $X2=13.587 $Y2=0.495
r1160 220 333 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.405 $Y=4.435
+ $X2=13.405 $Y2=4.52
r1161 219 478 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=13.405 $Y=3.685
+ $X2=13.405 $Y2=3.57
r1162 219 220 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=13.405 $Y=3.685
+ $X2=13.405 $Y2=4.435
r1163 218 473 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=13.405 $Y=1.755
+ $X2=13.405 $Y2=1.87
r1164 217 329 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.405 $Y=1.005
+ $X2=13.405 $Y2=0.92
r1165 217 218 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=13.405 $Y=1.005
+ $X2=13.405 $Y2=1.755
r1166 216 327 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.895 $Y=4.435
+ $X2=11.895 $Y2=4.52
r1167 215 472 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=11.895 $Y=3.685
+ $X2=11.895 $Y2=3.57
r1168 215 216 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=11.895 $Y=3.685
+ $X2=11.895 $Y2=4.435
r1169 214 467 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=11.895 $Y=1.755
+ $X2=11.895 $Y2=1.87
r1170 213 323 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.895 $Y=1.005
+ $X2=11.895 $Y2=0.92
r1171 213 214 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=11.895 $Y=1.005
+ $X2=11.895 $Y2=1.755
r1172 209 327 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=11.712 $Y=4.52
+ $X2=11.895 $Y2=4.52
r1173 209 211 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=11.712 $Y=4.605
+ $X2=11.712 $Y2=4.945
r1174 205 323 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=11.712 $Y=0.92
+ $X2=11.895 $Y2=0.92
r1175 205 207 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=11.712 $Y=0.835
+ $X2=11.712 $Y2=0.495
r1176 202 470 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=11.625 $Y=3.57
+ $X2=11.73 $Y2=3.57
r1177 201 319 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=11.625 $Y=3.14
+ $X2=11.625 $Y2=3.1
r1178 201 202 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=11.625 $Y=3.14
+ $X2=11.625 $Y2=3.455
r1179 198 317 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.625 $Y=2.3
+ $X2=11.625 $Y2=2.465
r1180 198 200 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=11.625 $Y=2.3
+ $X2=11.625 $Y2=2
r1181 197 465 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=11.625 $Y=1.87
+ $X2=11.73 $Y2=1.87
r1182 197 200 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.625 $Y=1.985
+ $X2=11.625 $Y2=2
r1183 196 460 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=9.535 $Y=3.57
+ $X2=9.43 $Y2=3.57
r1184 195 315 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=9.535 $Y=3.14
+ $X2=9.535 $Y2=3.1
r1185 195 196 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=9.535 $Y=3.14
+ $X2=9.535 $Y2=3.455
r1186 190 313 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.535 $Y=2.3
+ $X2=9.535 $Y2=2.465
r1187 190 192 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=9.535 $Y=2.3
+ $X2=9.535 $Y2=2
r1188 189 455 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=9.535 $Y=1.87
+ $X2=9.43 $Y2=1.87
r1189 189 192 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=9.535 $Y=1.985
+ $X2=9.535 $Y2=2
r1190 185 309 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=9.447 $Y=4.52
+ $X2=9.265 $Y2=4.52
r1191 185 187 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=9.447 $Y=4.605
+ $X2=9.447 $Y2=4.945
r1192 181 305 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=9.447 $Y=0.92
+ $X2=9.265 $Y2=0.92
r1193 181 183 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=9.447 $Y=0.835
+ $X2=9.447 $Y2=0.495
r1194 180 309 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=4.435
+ $X2=9.265 $Y2=4.52
r1195 179 458 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.265 $Y=3.685
+ $X2=9.265 $Y2=3.57
r1196 179 180 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=9.265 $Y=3.685
+ $X2=9.265 $Y2=4.435
r1197 178 453 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.265 $Y=1.755
+ $X2=9.265 $Y2=1.87
r1198 177 305 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=1.005
+ $X2=9.265 $Y2=0.92
r1199 177 178 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=9.265 $Y=1.005
+ $X2=9.265 $Y2=1.755
r1200 176 303 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.755 $Y=4.435
+ $X2=7.755 $Y2=4.52
r1201 175 452 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.755 $Y=3.685
+ $X2=7.755 $Y2=3.57
r1202 175 176 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=7.755 $Y=3.685
+ $X2=7.755 $Y2=4.435
r1203 174 447 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.755 $Y=1.755
+ $X2=7.755 $Y2=1.87
r1204 173 299 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.755 $Y=1.005
+ $X2=7.755 $Y2=0.92
r1205 173 174 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=7.755 $Y=1.005
+ $X2=7.755 $Y2=1.755
r1206 169 303 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=7.572 $Y=4.52
+ $X2=7.755 $Y2=4.52
r1207 169 171 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=7.572 $Y=4.605
+ $X2=7.572 $Y2=4.945
r1208 165 299 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=7.572 $Y=0.92
+ $X2=7.755 $Y2=0.92
r1209 165 167 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=7.572 $Y=0.835
+ $X2=7.572 $Y2=0.495
r1210 162 450 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=7.485 $Y=3.57
+ $X2=7.59 $Y2=3.57
r1211 161 295 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=7.485 $Y=3.14
+ $X2=7.485 $Y2=3.1
r1212 161 162 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=7.485 $Y=3.14
+ $X2=7.485 $Y2=3.455
r1213 158 293 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=2.3
+ $X2=7.485 $Y2=2.465
r1214 158 160 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=7.485 $Y=2.3
+ $X2=7.485 $Y2=2
r1215 157 445 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=7.485 $Y=1.87
+ $X2=7.59 $Y2=1.87
r1216 157 160 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.485 $Y=1.985
+ $X2=7.485 $Y2=2
r1217 156 440 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=3.57
+ $X2=5.29 $Y2=3.57
r1218 155 291 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=5.395 $Y=3.14
+ $X2=5.395 $Y2=3.1
r1219 155 156 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.395 $Y=3.14
+ $X2=5.395 $Y2=3.455
r1220 150 289 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.395 $Y=2.3
+ $X2=5.395 $Y2=2.465
r1221 150 152 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=5.395 $Y=2.3
+ $X2=5.395 $Y2=2
r1222 149 435 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=1.87
+ $X2=5.29 $Y2=1.87
r1223 149 152 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.395 $Y=1.985
+ $X2=5.395 $Y2=2
r1224 145 285 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=5.307 $Y=4.52
+ $X2=5.125 $Y2=4.52
r1225 145 147 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=5.307 $Y=4.605
+ $X2=5.307 $Y2=4.945
r1226 141 281 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=5.307 $Y=0.92
+ $X2=5.125 $Y2=0.92
r1227 141 143 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=5.307 $Y=0.835
+ $X2=5.307 $Y2=0.495
r1228 140 285 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=4.435
+ $X2=5.125 $Y2=4.52
r1229 139 438 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.125 $Y=3.685
+ $X2=5.125 $Y2=3.57
r1230 139 140 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.125 $Y=3.685
+ $X2=5.125 $Y2=4.435
r1231 138 433 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.125 $Y=1.755
+ $X2=5.125 $Y2=1.87
r1232 137 281 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=1.005
+ $X2=5.125 $Y2=0.92
r1233 137 138 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.125 $Y=1.005
+ $X2=5.125 $Y2=1.755
r1234 136 279 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=4.435
+ $X2=3.615 $Y2=4.52
r1235 135 432 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.615 $Y=3.685
+ $X2=3.615 $Y2=3.57
r1236 135 136 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.615 $Y=3.685
+ $X2=3.615 $Y2=4.435
r1237 134 427 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.615 $Y=1.755
+ $X2=3.615 $Y2=1.87
r1238 133 275 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=1.005
+ $X2=3.615 $Y2=0.92
r1239 133 134 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.615 $Y=1.005
+ $X2=3.615 $Y2=1.755
r1240 129 279 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=3.432 $Y=4.52
+ $X2=3.615 $Y2=4.52
r1241 129 131 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=3.432 $Y=4.605
+ $X2=3.432 $Y2=4.945
r1242 125 275 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=3.432 $Y=0.92
+ $X2=3.615 $Y2=0.92
r1243 125 127 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=3.432 $Y=0.835
+ $X2=3.432 $Y2=0.495
r1244 122 430 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=3.345 $Y=3.57
+ $X2=3.45 $Y2=3.57
r1245 121 271 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=3.345 $Y=3.14
+ $X2=3.345 $Y2=3.1
r1246 121 122 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.345 $Y=3.14
+ $X2=3.345 $Y2=3.455
r1247 118 269 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=2.3
+ $X2=3.345 $Y2=2.465
r1248 118 120 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.345 $Y=2.3
+ $X2=3.345 $Y2=2
r1249 117 425 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=3.345 $Y=1.87
+ $X2=3.45 $Y2=1.87
r1250 117 120 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.345 $Y=1.985
+ $X2=3.345 $Y2=2
r1251 116 420 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=1.255 $Y=3.57
+ $X2=1.15 $Y2=3.57
r1252 115 267 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=1.255 $Y=3.14
+ $X2=1.255 $Y2=3.1
r1253 115 116 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.255 $Y=3.14
+ $X2=1.255 $Y2=3.455
r1254 110 265 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=2.3
+ $X2=1.255 $Y2=2.465
r1255 110 112 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.255 $Y=2.3
+ $X2=1.255 $Y2=2
r1256 109 415 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=1.255 $Y=1.87
+ $X2=1.15 $Y2=1.87
r1257 109 112 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.255 $Y=1.985
+ $X2=1.255 $Y2=2
r1258 105 261 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=1.167 $Y=4.52
+ $X2=0.985 $Y2=4.52
r1259 105 107 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=1.167 $Y=4.605
+ $X2=1.167 $Y2=4.945
r1260 101 257 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=1.167 $Y=0.92
+ $X2=0.985 $Y2=0.92
r1261 101 103 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=1.167 $Y=0.835
+ $X2=1.167 $Y2=0.495
r1262 100 261 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=4.435
+ $X2=0.985 $Y2=4.52
r1263 99 418 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.985 $Y=3.685
+ $X2=0.985 $Y2=3.57
r1264 99 100 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.985 $Y=3.685
+ $X2=0.985 $Y2=4.435
r1265 98 413 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.985 $Y=1.755
+ $X2=0.985 $Y2=1.87
r1266 97 257 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=1.005
+ $X2=0.985 $Y2=0.92
r1267 97 98 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.985 $Y=1.005
+ $X2=0.985 $Y2=1.755
r1268 32 343 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=15.64
+ $Y=2.955 $X2=15.765 $Y2=3.1
r1269 31 240 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=15.64
+ $Y=1.665 $X2=15.765 $Y2=2
r1270 30 339 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=13.53
+ $Y=2.955 $X2=13.675 $Y2=3.1
r1271 29 232 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=13.53
+ $Y=1.665 $X2=13.675 $Y2=2
r1272 28 319 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=11.5
+ $Y=2.955 $X2=11.625 $Y2=3.1
r1273 27 200 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=11.5
+ $Y=1.665 $X2=11.625 $Y2=2
r1274 26 315 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.39
+ $Y=2.955 $X2=9.535 $Y2=3.1
r1275 25 192 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=9.39
+ $Y=1.665 $X2=9.535 $Y2=2
r1276 24 295 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=7.36
+ $Y=2.955 $X2=7.485 $Y2=3.1
r1277 23 160 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=7.36
+ $Y=1.665 $X2=7.485 $Y2=2
r1278 22 291 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.25
+ $Y=2.955 $X2=5.395 $Y2=3.1
r1279 21 152 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=5.25
+ $Y=1.665 $X2=5.395 $Y2=2
r1280 20 271 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=2.955 $X2=3.345 $Y2=3.1
r1281 19 120 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=1.665 $X2=3.345 $Y2=2
r1282 18 267 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=2.955 $X2=1.255 $Y2=3.1
r1283 17 112 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.665 $X2=1.255 $Y2=2
r1284 16 251 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=15.74
+ $Y=4.685 $X2=15.865 $Y2=4.945
r1285 15 247 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=15.74
+ $Y=0.235 $X2=15.865 $Y2=0.495
r1286 14 227 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=13.44
+ $Y=4.685 $X2=13.575 $Y2=4.945
r1287 13 223 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=13.44
+ $Y=0.235 $X2=13.575 $Y2=0.495
r1288 12 211 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=11.6
+ $Y=4.685 $X2=11.725 $Y2=4.945
r1289 11 207 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=11.6
+ $Y=0.235 $X2=11.725 $Y2=0.495
r1290 10 187 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.3
+ $Y=4.685 $X2=9.435 $Y2=4.945
r1291 9 183 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.3
+ $Y=0.235 $X2=9.435 $Y2=0.495
r1292 8 171 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=4.685 $X2=7.585 $Y2=4.945
r1293 7 167 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.585 $Y2=0.495
r1294 6 147 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=5.16
+ $Y=4.685 $X2=5.295 $Y2=4.945
r1295 5 143 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=5.16
+ $Y=0.235 $X2=5.295 $Y2=0.495
r1296 4 131 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=4.685 $X2=3.445 $Y2=4.945
r1297 3 127 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.235 $X2=3.445 $Y2=0.495
r1298 2 107 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=4.685 $X2=1.155 $Y2=4.945
r1299 1 103 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_1%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 55 57 59 61 65 69 73 77 81 85 89 93 97 101 105 109 113 117 119 121
+ 123 125 128 129 131 132 134 135 137 138 140 141 143 144 146 147 149 150 151
+ 152 153 154 155 156 157 158 159 160 185 192 213 220 241 248 269 276 290 293
+ 296 299 302 305
r408 281 282 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.33 $Y=5.44
+ $X2=16.33 $Y2=5.44
r409 279 282 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=14.95 $Y=5.44
+ $X2=16.33 $Y2=5.44
r410 278 281 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=14.95 $Y=5.44
+ $X2=16.33 $Y2=5.44
r411 278 279 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=5.44
+ $X2=14.95 $Y2=5.44
r412 276 311 4.07647 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=16.63 $Y=5.44
+ $X2=16.825 $Y2=5.44
r413 276 281 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=16.63 $Y=5.44
+ $X2=16.33 $Y2=5.44
r414 274 275 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.33 $Y=0
+ $X2=16.33 $Y2=0
r415 272 275 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=14.95 $Y=0
+ $X2=16.33 $Y2=0
r416 271 274 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=14.95 $Y=0
+ $X2=16.33 $Y2=0
r417 271 272 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r418 269 308 4.07647 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=16.63 $Y=0
+ $X2=16.825 $Y2=0
r419 269 274 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=16.63 $Y=0
+ $X2=16.33 $Y2=0
r420 268 279 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=5.44
+ $X2=14.95 $Y2=5.44
r421 267 268 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=5.44
+ $X2=14.49 $Y2=5.44
r422 265 268 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=13.11 $Y=5.44
+ $X2=14.49 $Y2=5.44
r423 264 267 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=13.11 $Y=5.44
+ $X2=14.49 $Y2=5.44
r424 264 265 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=5.44
+ $X2=13.11 $Y2=5.44
r425 262 305 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.81 $Y=5.44
+ $X2=12.65 $Y2=5.44
r426 262 264 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.81 $Y=5.44
+ $X2=13.11 $Y2=5.44
r427 261 272 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.95 $Y2=0
r428 260 261 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r429 258 261 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=14.49 $Y2=0
r430 257 260 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=13.11 $Y=0
+ $X2=14.49 $Y2=0
r431 257 258 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r432 255 302 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.81 $Y=0
+ $X2=12.65 $Y2=0
r433 255 257 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.81 $Y=0
+ $X2=13.11 $Y2=0
r434 253 254 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=5.44
+ $X2=12.19 $Y2=5.44
r435 251 254 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=10.81 $Y=5.44
+ $X2=12.19 $Y2=5.44
r436 250 253 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=10.81 $Y=5.44
+ $X2=12.19 $Y2=5.44
r437 250 251 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=5.44
+ $X2=10.81 $Y2=5.44
r438 248 305 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.49 $Y=5.44
+ $X2=12.65 $Y2=5.44
r439 248 253 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.49 $Y=5.44
+ $X2=12.19 $Y2=5.44
r440 246 247 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r441 244 247 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=12.19 $Y2=0
r442 243 246 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=10.81 $Y=0
+ $X2=12.19 $Y2=0
r443 243 244 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r444 241 302 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.49 $Y=0
+ $X2=12.65 $Y2=0
r445 241 246 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.49 $Y=0
+ $X2=12.19 $Y2=0
r446 240 251 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=5.44
+ $X2=10.81 $Y2=5.44
r447 239 240 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=5.44
+ $X2=10.35 $Y2=5.44
r448 237 240 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.97 $Y=5.44
+ $X2=10.35 $Y2=5.44
r449 236 239 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=8.97 $Y=5.44
+ $X2=10.35 $Y2=5.44
r450 236 237 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=5.44
+ $X2=8.97 $Y2=5.44
r451 234 299 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.67 $Y=5.44
+ $X2=8.51 $Y2=5.44
r452 234 236 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.67 $Y=5.44
+ $X2=8.97 $Y2=5.44
r453 233 244 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r454 232 233 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r455 230 233 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=10.35 $Y2=0
r456 229 232 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=8.97 $Y=0
+ $X2=10.35 $Y2=0
r457 229 230 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r458 227 296 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.67 $Y=0 $X2=8.51
+ $Y2=0
r459 227 229 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.67 $Y=0 $X2=8.97
+ $Y2=0
r460 225 226 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=5.44
+ $X2=8.05 $Y2=5.44
r461 223 226 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=5.44
+ $X2=8.05 $Y2=5.44
r462 222 225 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.67 $Y=5.44
+ $X2=8.05 $Y2=5.44
r463 222 223 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=5.44
+ $X2=6.67 $Y2=5.44
r464 220 299 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.35 $Y=5.44
+ $X2=8.51 $Y2=5.44
r465 220 225 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.35 $Y=5.44
+ $X2=8.05 $Y2=5.44
r466 218 219 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r467 216 219 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=8.05 $Y2=0
r468 215 218 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=8.05 $Y2=0
r469 215 216 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r470 213 296 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.35 $Y=0 $X2=8.51
+ $Y2=0
r471 213 218 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.35 $Y=0 $X2=8.05
+ $Y2=0
r472 212 223 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=5.44
+ $X2=6.67 $Y2=5.44
r473 211 212 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=5.44
+ $X2=6.21 $Y2=5.44
r474 209 212 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=5.44
+ $X2=6.21 $Y2=5.44
r475 208 211 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=5.44
+ $X2=6.21 $Y2=5.44
r476 208 209 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=5.44
+ $X2=4.83 $Y2=5.44
r477 206 293 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.53 $Y=5.44
+ $X2=4.37 $Y2=5.44
r478 206 208 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.53 $Y=5.44
+ $X2=4.83 $Y2=5.44
r479 205 216 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=6.67 $Y2=0
r480 204 205 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r481 202 205 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.21 $Y2=0
r482 201 204 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=6.21 $Y2=0
r483 201 202 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r484 199 290 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.37
+ $Y2=0
r485 199 201 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.83
+ $Y2=0
r486 197 198 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=5.44
+ $X2=3.91 $Y2=5.44
r487 195 198 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=5.44
+ $X2=3.91 $Y2=5.44
r488 194 197 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=5.44
+ $X2=3.91 $Y2=5.44
r489 194 195 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=5.44
+ $X2=2.53 $Y2=5.44
r490 192 293 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.21 $Y=5.44
+ $X2=4.37 $Y2=5.44
r491 192 197 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.21 $Y=5.44
+ $X2=3.91 $Y2=5.44
r492 190 191 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r493 188 191 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r494 187 190 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r495 187 188 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r496 185 290 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.37
+ $Y2=0
r497 185 190 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=3.91
+ $Y2=0
r498 184 195 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=5.44
+ $X2=2.53 $Y2=5.44
r499 183 184 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=5.44
+ $X2=2.07 $Y2=5.44
r500 181 184 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=5.44
+ $X2=2.07 $Y2=5.44
r501 180 183 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=5.44
+ $X2=2.07 $Y2=5.44
r502 180 181 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=5.44
+ $X2=0.69 $Y2=5.44
r503 178 287 4.07647 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=5.44
+ $X2=0.195 $Y2=5.44
r504 178 180 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=5.44
+ $X2=0.69 $Y2=5.44
r505 177 188 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.53 $Y2=0
r506 176 177 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r507 174 177 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r508 173 176 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r509 173 174 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r510 171 284 4.07647 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0
+ $X2=0.195 $Y2=0
r511 171 173 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.69
+ $Y2=0
r512 160 282 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=16.79 $Y=5.44
+ $X2=16.33 $Y2=5.44
r513 160 311 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.79 $Y=5.44
+ $X2=16.79 $Y2=5.44
r514 159 275 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=16.79 $Y=0
+ $X2=16.33 $Y2=0
r515 159 308 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.79 $Y=0
+ $X2=16.79 $Y2=0
r516 158 265 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=5.44
+ $X2=13.11 $Y2=5.44
r517 158 254 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=5.44
+ $X2=12.19 $Y2=5.44
r518 158 305 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=5.44
+ $X2=12.65 $Y2=5.44
r519 157 258 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r520 157 247 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r521 157 302 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r522 156 237 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=5.44
+ $X2=8.97 $Y2=5.44
r523 156 226 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=5.44
+ $X2=8.05 $Y2=5.44
r524 156 299 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=5.44
+ $X2=8.51 $Y2=5.44
r525 155 230 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.97 $Y2=0
r526 155 219 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r527 155 296 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r528 154 209 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=5.44
+ $X2=4.83 $Y2=5.44
r529 154 198 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=5.44
+ $X2=3.91 $Y2=5.44
r530 154 293 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=5.44
+ $X2=4.37 $Y2=5.44
r531 153 202 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r532 153 191 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=3.91 $Y2=0
r533 153 290 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r534 152 181 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=5.44
+ $X2=0.69 $Y2=5.44
r535 152 287 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=5.44
+ $X2=0.23 $Y2=5.44
r536 151 174 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r537 151 284 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r538 149 267 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.555 $Y=5.44
+ $X2=14.49 $Y2=5.44
r539 149 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.555 $Y=5.44
+ $X2=14.72 $Y2=5.44
r540 148 278 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.885 $Y=5.44
+ $X2=14.95 $Y2=5.44
r541 148 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.885 $Y=5.44
+ $X2=14.72 $Y2=5.44
r542 146 260 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.555 $Y=0
+ $X2=14.49 $Y2=0
r543 146 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.555 $Y=0
+ $X2=14.72 $Y2=0
r544 145 271 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.885 $Y=0
+ $X2=14.95 $Y2=0
r545 145 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.885 $Y=0
+ $X2=14.72 $Y2=0
r546 143 239 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.415 $Y=5.44
+ $X2=10.35 $Y2=5.44
r547 143 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=5.44
+ $X2=10.58 $Y2=5.44
r548 142 250 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.745 $Y=5.44
+ $X2=10.81 $Y2=5.44
r549 142 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.745 $Y=5.44
+ $X2=10.58 $Y2=5.44
r550 140 232 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.415 $Y=0
+ $X2=10.35 $Y2=0
r551 140 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=0
+ $X2=10.58 $Y2=0
r552 139 243 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.745 $Y=0
+ $X2=10.81 $Y2=0
r553 139 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.745 $Y=0
+ $X2=10.58 $Y2=0
r554 137 211 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.275 $Y=5.44
+ $X2=6.21 $Y2=5.44
r555 137 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=5.44
+ $X2=6.44 $Y2=5.44
r556 136 222 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=5.44
+ $X2=6.67 $Y2=5.44
r557 136 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=5.44
+ $X2=6.44 $Y2=5.44
r558 134 204 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.275 $Y=0
+ $X2=6.21 $Y2=0
r559 134 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=0
+ $X2=6.44 $Y2=0
r560 133 215 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=0
+ $X2=6.67 $Y2=0
r561 133 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=0
+ $X2=6.44 $Y2=0
r562 131 183 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=5.44
+ $X2=2.07 $Y2=5.44
r563 131 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=5.44
+ $X2=2.3 $Y2=5.44
r564 130 194 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.465 $Y=5.44
+ $X2=2.53 $Y2=5.44
r565 130 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=5.44
+ $X2=2.3 $Y2=5.44
r566 128 176 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=0
+ $X2=2.07 $Y2=0
r567 128 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0
+ $X2=2.3 $Y2=0
r568 127 187 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.465 $Y=0
+ $X2=2.53 $Y2=0
r569 127 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0
+ $X2=2.3 $Y2=0
r570 123 311 3.13575 $w=2.6e-07 $l=1.12916e-07 $layer=LI1_cond $X=16.76 $Y=5.355
+ $X2=16.825 $Y2=5.44
r571 123 125 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=16.76 $Y=5.355
+ $X2=16.76 $Y2=4.72
r572 119 308 3.13575 $w=2.6e-07 $l=1.12916e-07 $layer=LI1_cond $X=16.76 $Y=0.085
+ $X2=16.825 $Y2=0
r573 119 121 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=16.76 $Y=0.085
+ $X2=16.76 $Y2=0.38
r574 115 150 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.72 $Y=5.355
+ $X2=14.72 $Y2=5.44
r575 115 117 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=14.72 $Y=5.355
+ $X2=14.72 $Y2=4.945
r576 111 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.72 $Y=0.085
+ $X2=14.72 $Y2=0
r577 111 113 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=14.72 $Y=0.085
+ $X2=14.72 $Y2=0.495
r578 107 305 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=12.65 $Y=5.355
+ $X2=12.65 $Y2=5.44
r579 107 109 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=12.65 $Y=5.355
+ $X2=12.65 $Y2=4.72
r580 103 302 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=12.65 $Y=0.085
+ $X2=12.65 $Y2=0
r581 103 105 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=12.65 $Y=0.085
+ $X2=12.65 $Y2=0.38
r582 99 144 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.58 $Y=5.355
+ $X2=10.58 $Y2=5.44
r583 99 101 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.58 $Y=5.355
+ $X2=10.58 $Y2=4.945
r584 95 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.58 $Y=0.085
+ $X2=10.58 $Y2=0
r585 95 97 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.58 $Y=0.085
+ $X2=10.58 $Y2=0.495
r586 91 299 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.51 $Y=5.355
+ $X2=8.51 $Y2=5.44
r587 91 93 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=8.51 $Y=5.355
+ $X2=8.51 $Y2=4.72
r588 87 296 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.51 $Y=0.085
+ $X2=8.51 $Y2=0
r589 87 89 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=8.51 $Y=0.085
+ $X2=8.51 $Y2=0.38
r590 83 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=5.355
+ $X2=6.44 $Y2=5.44
r591 83 85 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.44 $Y=5.355
+ $X2=6.44 $Y2=4.945
r592 79 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0
r593 79 81 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0.495
r594 75 293 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=5.355
+ $X2=4.37 $Y2=5.44
r595 75 77 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=4.37 $Y=5.355
+ $X2=4.37 $Y2=4.72
r596 71 290 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0
r597 71 73 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0.38
r598 67 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=5.355
+ $X2=2.3 $Y2=5.44
r599 67 69 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.3 $Y=5.355
+ $X2=2.3 $Y2=4.945
r600 63 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=0.085
+ $X2=2.3 $Y2=0
r601 63 65 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.3 $Y=0.085
+ $X2=2.3 $Y2=0.495
r602 59 287 3.13575 $w=2.6e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.26 $Y=5.355
+ $X2=0.195 $Y2=5.44
r603 59 61 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=5.355
+ $X2=0.26 $Y2=4.72
r604 55 284 3.13575 $w=2.6e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.195 $Y2=0
r605 55 57 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r606 18 125 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=16.625
+ $Y=4.555 $X2=16.76 $Y2=4.72
r607 17 121 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=16.625
+ $Y=0.235 $X2=16.76 $Y2=0.38
r608 16 117 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=14.505
+ $Y=4.685 $X2=14.72 $Y2=4.945
r609 15 113 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=14.505
+ $Y=0.235 $X2=14.72 $Y2=0.495
r610 14 109 91 $w=1.7e-07 $l=2.33345e-07 $layer=licon1_NDIFF $count=2 $X=12.485
+ $Y=4.555 $X2=12.65 $Y2=4.72
r611 13 105 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=12.485
+ $Y=0.235 $X2=12.65 $Y2=0.38
r612 12 101 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=10.365
+ $Y=4.685 $X2=10.58 $Y2=4.945
r613 11 97 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=10.365
+ $Y=0.235 $X2=10.58 $Y2=0.495
r614 10 93 91 $w=1.7e-07 $l=2.33345e-07 $layer=licon1_NDIFF $count=2 $X=8.345
+ $Y=4.555 $X2=8.51 $Y2=4.72
r615 9 89 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=8.345
+ $Y=0.235 $X2=8.51 $Y2=0.38
r616 8 85 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=6.225
+ $Y=4.685 $X2=6.44 $Y2=4.945
r617 7 81 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=6.225
+ $Y=0.235 $X2=6.44 $Y2=0.495
r618 6 77 91 $w=1.7e-07 $l=2.33345e-07 $layer=licon1_NDIFF $count=2 $X=4.205
+ $Y=4.555 $X2=4.37 $Y2=4.72
r619 5 73 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=4.205
+ $Y=0.235 $X2=4.37 $Y2=0.38
r620 4 69 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=4.685 $X2=2.3 $Y2=4.945
r621 3 65 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.235 $X2=2.3 $Y2=0.495
r622 2 61 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=4.555 $X2=0.26 $Y2=4.72
r623 1 57 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

