* File: sky130_fd_sc_hdll__a221oi_2.pxi.spice
* Created: Wed Sep  2 08:18:09 2020
* 
x_PM_SKY130_FD_SC_HDLL__A221OI_2%C1 N_C1_c_90_n N_C1_M1004_g N_C1_c_86_n
+ N_C1_M1007_g N_C1_c_91_n N_C1_M1018_g N_C1_c_87_n N_C1_M1016_g C1 C1
+ N_C1_c_89_n PM_SKY130_FD_SC_HDLL__A221OI_2%C1
x_PM_SKY130_FD_SC_HDLL__A221OI_2%B2 N_B2_c_126_n N_B2_M1008_g N_B2_c_127_n
+ N_B2_M1010_g N_B2_c_128_n N_B2_M1019_g N_B2_c_129_n N_B2_M1017_g N_B2_c_134_n
+ N_B2_c_130_n B2 B2 PM_SKY130_FD_SC_HDLL__A221OI_2%B2
x_PM_SKY130_FD_SC_HDLL__A221OI_2%B1 N_B1_c_203_n N_B1_M1000_g N_B1_c_207_n
+ N_B1_M1001_g N_B1_c_208_n N_B1_M1005_g N_B1_c_204_n N_B1_M1011_g B1
+ N_B1_c_206_n B1 PM_SKY130_FD_SC_HDLL__A221OI_2%B1
x_PM_SKY130_FD_SC_HDLL__A221OI_2%A2 N_A2_c_247_n N_A2_M1002_g N_A2_c_248_n
+ N_A2_M1003_g N_A2_c_249_n N_A2_M1009_g N_A2_c_250_n N_A2_M1012_g N_A2_c_251_n
+ N_A2_c_258_n N_A2_c_259_n N_A2_c_252_n N_A2_c_253_n A2 A2
+ PM_SKY130_FD_SC_HDLL__A221OI_2%A2
x_PM_SKY130_FD_SC_HDLL__A221OI_2%A1 N_A1_c_324_n N_A1_M1006_g N_A1_c_328_n
+ N_A1_M1013_g N_A1_c_329_n N_A1_M1015_g N_A1_c_325_n N_A1_M1014_g A1
+ N_A1_c_327_n A1 PM_SKY130_FD_SC_HDLL__A221OI_2%A1
x_PM_SKY130_FD_SC_HDLL__A221OI_2%A_27_297# N_A_27_297#_M1004_s
+ N_A_27_297#_M1018_s N_A_27_297#_M1008_d N_A_27_297#_M1005_d
+ N_A_27_297#_c_369_n N_A_27_297#_c_370_n N_A_27_297#_c_371_n
+ N_A_27_297#_c_372_n N_A_27_297#_c_373_n N_A_27_297#_c_374_n
+ N_A_27_297#_c_395_n N_A_27_297#_c_375_n N_A_27_297#_c_396_n
+ N_A_27_297#_c_398_n PM_SKY130_FD_SC_HDLL__A221OI_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A221OI_2%Y N_Y_M1007_s N_Y_M1000_d N_Y_M1006_d
+ N_Y_M1004_d N_Y_c_431_n N_Y_c_432_n N_Y_c_433_n N_Y_c_434_n N_Y_c_435_n
+ N_Y_c_436_n Y Y Y Y Y N_Y_c_446_n PM_SKY130_FD_SC_HDLL__A221OI_2%Y
x_PM_SKY130_FD_SC_HDLL__A221OI_2%A_321_297# N_A_321_297#_M1008_s
+ N_A_321_297#_M1001_s N_A_321_297#_M1019_s N_A_321_297#_M1013_s
+ N_A_321_297#_M1009_s N_A_321_297#_c_509_n N_A_321_297#_c_510_n
+ N_A_321_297#_c_511_n N_A_321_297#_c_517_n N_A_321_297#_c_550_p
+ N_A_321_297#_c_520_n N_A_321_297#_c_505_n N_A_321_297#_c_551_p
+ N_A_321_297#_c_538_n N_A_321_297#_c_541_n N_A_321_297#_c_526_n
+ PM_SKY130_FD_SC_HDLL__A221OI_2%A_321_297#
x_PM_SKY130_FD_SC_HDLL__A221OI_2%VPWR N_VPWR_M1002_d N_VPWR_M1015_d
+ N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n
+ N_VPWR_c_571_n VPWR N_VPWR_c_572_n N_VPWR_c_565_n
+ PM_SKY130_FD_SC_HDLL__A221OI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A221OI_2%VGND N_VGND_M1007_d N_VGND_M1016_d
+ N_VGND_M1017_d N_VGND_M1012_s N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n
+ N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n N_VGND_c_640_n N_VGND_c_641_n
+ VGND N_VGND_c_642_n N_VGND_c_643_n N_VGND_c_644_n N_VGND_c_645_n
+ PM_SKY130_FD_SC_HDLL__A221OI_2%VGND
x_PM_SKY130_FD_SC_HDLL__A221OI_2%A_413_47# N_A_413_47#_M1010_s
+ N_A_413_47#_M1011_s N_A_413_47#_c_706_n
+ PM_SKY130_FD_SC_HDLL__A221OI_2%A_413_47#
x_PM_SKY130_FD_SC_HDLL__A221OI_2%A_805_47# N_A_805_47#_M1003_d
+ N_A_805_47#_M1014_s N_A_805_47#_c_721_n N_A_805_47#_c_738_n
+ N_A_805_47#_c_720_n PM_SKY130_FD_SC_HDLL__A221OI_2%A_805_47#
cc_1 VNB N_C1_c_86_n 0.0220726f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.995
cc_2 VNB N_C1_c_87_n 0.0219182f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.995
cc_3 VNB C1 0.00916578f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_C1_c_89_n 0.0706227f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.202
cc_5 VNB N_B2_c_126_n 0.0288833f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.41
cc_6 VNB N_B2_c_127_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.995
cc_7 VNB N_B2_c_128_n 0.0221931f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_8 VNB N_B2_c_129_n 0.0177944f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.995
cc_9 VNB N_B2_c_130_n 0.00349767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB B2 0.00662148f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.202
cc_11 VNB N_B1_c_203_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.41
cc_12 VNB N_B1_c_204_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.995
cc_13 VNB B1 0.00141641f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_14 VNB N_B1_c_206_n 0.0356367f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.202
cc_15 VNB N_A2_c_247_n 0.023686f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.41
cc_16 VNB N_A2_c_248_n 0.017338f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.995
cc_17 VNB N_A2_c_249_n 0.0316217f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_18 VNB N_A2_c_250_n 0.0221358f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.995
cc_19 VNB N_A2_c_251_n 0.0016889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_252_n 2.72331e-19 $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.202
cc_21 VNB N_A2_c_253_n 0.00192755f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.202
cc_22 VNB A2 0.0277194f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.202
cc_23 VNB N_A1_c_324_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.41
cc_24 VNB N_A1_c_325_n 0.0176137f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.995
cc_25 VNB A1 0.00231079f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_26 VNB N_A1_c_327_n 0.0356362f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.202
cc_27 VNB N_Y_c_431_n 8.41399e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_432_n 7.40341e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_433_n 0.023424f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.202
cc_30 VNB N_Y_c_434_n 0.00100041f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.202
cc_31 VNB N_Y_c_435_n 0.00278017f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_32 VNB N_Y_c_436_n 0.0144439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB Y 0.00172183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_565_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_634_n 0.010359f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_36 VNB N_VGND_c_635_n 0.0311542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_636_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.202
cc_38 VNB N_VGND_c_637_n 0.00712566f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_638_n 0.0413805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_639_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_640_n 0.0419047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_641_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_642_n 0.0124854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_643_n 0.302528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_644_n 0.0203884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_645_n 0.0208826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_805_47#_c_720_n 0.00285684f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_48 VPB N_C1_c_90_n 0.0196012f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.41
cc_49 VPB N_C1_c_91_n 0.0195801f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_50 VPB C1 0.0121511f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_51 VPB N_C1_c_89_n 0.0324367f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.202
cc_52 VPB N_B2_c_126_n 0.0301044f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.41
cc_53 VPB N_B2_c_128_n 0.0256643f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_54 VPB N_B2_c_134_n 0.00683421f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_55 VPB N_B2_c_130_n 0.00272899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB B2 0.0045697f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.202
cc_57 VPB N_B1_c_207_n 0.0159948f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.995
cc_58 VPB N_B1_c_208_n 0.0159958f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_59 VPB N_B1_c_206_n 0.0192932f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.202
cc_60 VPB N_A2_c_247_n 0.025619f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.41
cc_61 VPB N_A2_c_249_n 0.0331355f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_62 VPB N_A2_c_251_n 0.0021804f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A2_c_258_n 0.00783392f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_64 VPB N_A2_c_259_n 2.51985e-19 $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_65 VPB N_A2_c_252_n 0.00130718f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.202
cc_66 VPB N_A1_c_328_n 0.0159602f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.995
cc_67 VPB N_A1_c_329_n 0.0159756f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_68 VPB N_A1_c_327_n 0.0192976f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.202
cc_69 VPB N_A_27_297#_c_369_n 0.0198753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_297#_c_370_n 0.00190269f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.202
cc_71 VPB N_A_27_297#_c_371_n 0.00752692f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_72 VPB N_A_27_297#_c_372_n 0.00444976f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.202
cc_73 VPB N_A_27_297#_c_373_n 0.00410721f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_74 VPB N_A_27_297#_c_374_n 0.0129913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_297#_c_375_n 2.51509e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB Y 9.48779e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_321_297#_c_505_n 0.00341263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_566_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_79 VPB N_VPWR_c_567_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_80 VPB N_VPWR_c_568_n 0.0971875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_569_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.202
cc_82 VPB N_VPWR_c_570_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_83 VPB N_VPWR_c_571_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.202
cc_84 VPB N_VPWR_c_572_n 0.0242591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_565_n 0.0546019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 N_C1_c_91_n B2 0.00216536f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_87 N_C1_c_89_n B2 0.00901847f $X=0.975 $Y=1.202 $X2=0 $Y2=0
cc_88 C1 N_A_27_297#_M1004_s 0.00307229f $X=0.15 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_89 N_C1_c_90_n N_A_27_297#_c_369_n 0.00864808f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_90 N_C1_c_91_n N_A_27_297#_c_369_n 7.21945e-19 $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_91 C1 N_A_27_297#_c_369_n 0.0230777f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_92 N_C1_c_89_n N_A_27_297#_c_369_n 0.00115707f $X=0.975 $Y=1.202 $X2=0 $Y2=0
cc_93 N_C1_c_90_n N_A_27_297#_c_370_n 0.0129846f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_94 N_C1_c_91_n N_A_27_297#_c_370_n 0.0137768f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_95 N_C1_c_90_n N_A_27_297#_c_371_n 4.32652e-19 $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_96 N_C1_c_91_n N_A_27_297#_c_373_n 0.00723112f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_97 N_C1_c_91_n N_A_27_297#_c_375_n 0.00280942f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_98 N_C1_c_87_n N_Y_c_433_n 0.0174521f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_99 N_C1_c_90_n Y 6.46595e-19 $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_100 N_C1_c_86_n Y 0.00899777f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_101 N_C1_c_91_n Y 0.0123856f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_102 N_C1_c_87_n Y 0.00252485f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_103 C1 Y 0.0336807f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_104 N_C1_c_89_n Y 0.0456611f $X=0.975 $Y=1.202 $X2=0 $Y2=0
cc_105 N_C1_c_86_n N_Y_c_446_n 0.00684661f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_106 N_C1_c_90_n N_VPWR_c_568_n 0.00429425f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_107 N_C1_c_91_n N_VPWR_c_568_n 0.00429453f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_108 N_C1_c_90_n N_VPWR_c_565_n 0.0069856f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_109 N_C1_c_91_n N_VPWR_c_565_n 0.00734734f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_110 N_C1_c_86_n N_VGND_c_635_n 0.00733912f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_111 C1 N_VGND_c_635_n 0.0208398f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_112 N_C1_c_89_n N_VGND_c_635_n 0.00623008f $X=0.975 $Y=1.202 $X2=0 $Y2=0
cc_113 N_C1_c_86_n N_VGND_c_643_n 0.00891986f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_114 N_C1_c_87_n N_VGND_c_643_n 0.00733728f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_115 N_C1_c_86_n N_VGND_c_644_n 0.00470854f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_116 N_C1_c_87_n N_VGND_c_644_n 0.00437852f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C1_c_87_n N_VGND_c_645_n 0.00481673f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B2_c_127_n N_B1_c_203_n 0.0268983f $X=1.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_119 N_B2_c_126_n N_B1_c_207_n 0.036701f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B2_c_134_n N_B1_c_207_n 0.0112877f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_121 B2 N_B1_c_207_n 0.00111092f $X=1.955 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B2_c_128_n N_B1_c_208_n 0.0367644f $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B2_c_134_n N_B1_c_208_n 0.011241f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_124 N_B2_c_130_n N_B1_c_208_n 0.00101445f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_125 N_B2_c_129_n N_B1_c_204_n 0.0223996f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B2_c_126_n B1 2.06946e-19 $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_127 N_B2_c_128_n B1 6.86695e-19 $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B2_c_134_n B1 0.0461557f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_129 N_B2_c_130_n B1 0.0176354f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_130 B2 B1 0.0169932f $X=1.955 $Y=1.105 $X2=0 $Y2=0
cc_131 N_B2_c_126_n N_B1_c_206_n 0.0263618f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B2_c_128_n N_B1_c_206_n 0.0263033f $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_133 N_B2_c_134_n N_B1_c_206_n 0.00803891f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_134 N_B2_c_130_n N_B1_c_206_n 0.00392336f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_135 B2 N_B1_c_206_n 0.00489839f $X=1.955 $Y=1.105 $X2=0 $Y2=0
cc_136 N_B2_c_128_n N_A2_c_247_n 0.0396157f $X=3.375 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_137 N_B2_c_130_n N_A2_c_247_n 0.00168246f $X=3.35 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_138 N_B2_c_129_n N_A2_c_248_n 0.0217201f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B2_c_128_n N_A2_c_251_n 0.00113531f $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B2_c_130_n N_A2_c_251_n 0.0310908f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B2_c_128_n N_A2_c_259_n 5.73459e-19 $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B2_c_130_n N_A2_c_259_n 0.0147563f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_143 N_B2_c_134_n N_A_27_297#_M1008_d 0.00135043f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_144 B2 N_A_27_297#_M1008_d 0.00115658f $X=1.955 $Y=1.105 $X2=0 $Y2=0
cc_145 N_B2_c_134_n N_A_27_297#_M1005_d 0.00171997f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_146 N_B2_c_130_n N_A_27_297#_M1005_d 7.75307e-19 $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B2_c_126_n N_A_27_297#_c_372_n 0.00496988f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_148 B2 N_A_27_297#_c_372_n 0.00582192f $X=1.955 $Y=1.105 $X2=0 $Y2=0
cc_149 N_B2_c_126_n N_A_27_297#_c_373_n 0.00442724f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B2_c_126_n N_A_27_297#_c_374_n 0.0130414f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_151 B2 N_A_27_297#_c_374_n 0.0203631f $X=1.955 $Y=1.105 $X2=0 $Y2=0
cc_152 N_B2_c_134_n N_A_27_297#_c_395_n 0.0371166f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_153 N_B2_c_134_n N_A_27_297#_c_396_n 0.00754343f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_154 B2 N_A_27_297#_c_396_n 0.00648665f $X=1.955 $Y=1.105 $X2=0 $Y2=0
cc_155 N_B2_c_134_n N_A_27_297#_c_398_n 0.0102375f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_156 N_B2_c_130_n N_A_27_297#_c_398_n 0.00353817f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_157 N_B2_c_127_n N_Y_c_432_n 4.05448e-19 $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_158 N_B2_c_126_n N_Y_c_433_n 0.00437722f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_159 N_B2_c_127_n N_Y_c_433_n 0.0139778f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B2_c_134_n N_Y_c_433_n 0.01139f $X=3.185 $Y=1.53 $X2=0 $Y2=0
cc_161 B2 N_Y_c_433_n 0.036129f $X=1.955 $Y=1.105 $X2=0 $Y2=0
cc_162 N_B2_c_128_n N_Y_c_436_n 0.00437722f $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_163 N_B2_c_129_n N_Y_c_436_n 0.0134071f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B2_c_130_n N_Y_c_436_n 0.0294729f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_165 B2 N_A_321_297#_M1008_s 0.00285498f $X=1.955 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_166 N_B2_c_134_n N_A_321_297#_M1001_s 0.00187547f $X=3.185 $Y=1.53 $X2=0
+ $Y2=0
cc_167 N_B2_c_130_n N_A_321_297#_M1019_s 0.00158406f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B2_c_126_n N_A_321_297#_c_509_n 0.0099733f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B2_c_128_n N_A_321_297#_c_510_n 0.0143148f $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B2_c_130_n N_A_321_297#_c_511_n 0.00345721f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_171 N_B2_c_126_n N_VPWR_c_568_n 0.00429453f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B2_c_128_n N_VPWR_c_568_n 0.00429453f $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_173 N_B2_c_126_n N_VPWR_c_565_n 0.00737353f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B2_c_128_n N_VPWR_c_565_n 0.00629441f $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B2_c_129_n N_VGND_c_636_n 0.00533053f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B2_c_127_n N_VGND_c_638_n 0.00395199f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B2_c_129_n N_VGND_c_638_n 0.00437852f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B2_c_127_n N_VGND_c_643_n 0.00692334f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B2_c_129_n N_VGND_c_643_n 0.00645862f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B2_c_127_n N_VGND_c_645_n 0.00770185f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B2_c_127_n N_A_413_47#_c_706_n 0.005151f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_182 N_B1_c_207_n N_A_27_297#_c_395_n 0.0108425f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B1_c_208_n N_A_27_297#_c_395_n 0.0108425f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_184 N_B1_c_206_n N_Y_c_431_n 0.00473056f $X=2.905 $Y=1.202 $X2=0 $Y2=0
cc_185 N_B1_c_203_n N_Y_c_432_n 0.00408314f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_203_n N_Y_c_433_n 0.00696451f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_187 B1 N_Y_c_433_n 0.0473377f $X=2.67 $Y=1.105 $X2=0 $Y2=0
cc_188 N_B1_c_204_n N_Y_c_436_n 0.009629f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_207_n N_A_321_297#_c_509_n 0.0099733f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_190 N_B1_c_208_n N_A_321_297#_c_510_n 0.0099733f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B1_c_207_n N_VPWR_c_568_n 0.00429453f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B1_c_208_n N_VPWR_c_568_n 0.00429453f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B1_c_207_n N_VPWR_c_565_n 0.00609118f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B1_c_208_n N_VPWR_c_565_n 0.00609118f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_195 N_B1_c_203_n N_VGND_c_638_n 0.00357877f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B1_c_204_n N_VGND_c_638_n 0.00357877f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_197 N_B1_c_203_n N_VGND_c_643_n 0.005504f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B1_c_204_n N_VGND_c_643_n 0.00562222f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B1_c_203_n N_A_413_47#_c_706_n 0.00996116f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_200 N_B1_c_204_n N_A_413_47#_c_706_n 0.0101195f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A2_c_248_n N_A1_c_324_n 0.0269138f $X=3.95 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_202 N_A2_c_247_n N_A1_c_328_n 0.0372206f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A2_c_251_n N_A1_c_328_n 7.438e-19 $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A2_c_258_n N_A1_c_328_n 0.011867f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_205 N_A2_c_249_n N_A1_c_329_n 0.0364739f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A2_c_258_n N_A1_c_329_n 0.0130886f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_207 N_A2_c_252_n N_A1_c_329_n 7.34002e-19 $X=5.185 $Y=1.445 $X2=0 $Y2=0
cc_208 N_A2_c_250_n N_A1_c_325_n 0.0102225f $X=5.36 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A2_c_247_n A1 0.00125115f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A2_c_251_n A1 0.0166975f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A2_c_258_n A1 0.0482519f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_212 N_A2_c_253_n A1 0.0165531f $X=5.27 $Y=1.175 $X2=0 $Y2=0
cc_213 N_A2_c_247_n N_A1_c_327_n 0.0260737f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A2_c_249_n N_A1_c_327_n 0.026336f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A2_c_251_n N_A1_c_327_n 0.00245121f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A2_c_258_n N_A1_c_327_n 0.00816189f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_217 N_A2_c_252_n N_A1_c_327_n 0.0029218f $X=5.185 $Y=1.445 $X2=0 $Y2=0
cc_218 N_A2_c_253_n N_A1_c_327_n 0.00152454f $X=5.27 $Y=1.175 $X2=0 $Y2=0
cc_219 N_A2_c_248_n N_Y_c_435_n 3.90453e-19 $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A2_c_247_n N_Y_c_436_n 0.00448367f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A2_c_248_n N_Y_c_436_n 0.0124133f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_c_251_n N_Y_c_436_n 0.0254056f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A2_c_258_n N_Y_c_436_n 0.00574727f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_224 N_A2_c_259_n N_A_321_297#_M1019_s 0.00159543f $X=4.065 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A2_c_258_n N_A_321_297#_M1013_s 0.00187091f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_226 N_A2_c_259_n N_A_321_297#_c_511_n 0.00354737f $X=4.065 $Y=1.53 $X2=0
+ $Y2=0
cc_227 N_A2_c_247_n N_A_321_297#_c_517_n 0.0112531f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A2_c_258_n N_A_321_297#_c_517_n 0.02495f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_229 N_A2_c_259_n N_A_321_297#_c_517_n 0.0135462f $X=4.065 $Y=1.53 $X2=0 $Y2=0
cc_230 N_A2_c_249_n N_A_321_297#_c_520_n 0.0139685f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A2_c_258_n N_A_321_297#_c_520_n 0.0273762f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_232 A2 N_A_321_297#_c_520_n 0.00534422f $X=5.64 $Y=1.105 $X2=0 $Y2=0
cc_233 N_A2_c_249_n N_A_321_297#_c_505_n 0.004595f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A2_c_258_n N_A_321_297#_c_505_n 0.0104762f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_235 A2 N_A_321_297#_c_505_n 0.0166332f $X=5.64 $Y=1.105 $X2=0 $Y2=0
cc_236 N_A2_c_258_n N_A_321_297#_c_526_n 0.0143191f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_237 N_A2_c_258_n N_VPWR_M1002_d 0.00187547f $X=5.1 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_238 N_A2_c_258_n N_VPWR_M1015_d 0.00189646f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_239 N_A2_c_247_n N_VPWR_c_566_n 0.00300743f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A2_c_249_n N_VPWR_c_567_n 0.00300743f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A2_c_247_n N_VPWR_c_568_n 0.00702461f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A2_c_249_n N_VPWR_c_572_n 0.00702461f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A2_c_247_n N_VPWR_c_565_n 0.00716301f $X=3.925 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A2_c_249_n N_VPWR_c_565_n 0.00798376f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A2_c_248_n N_VGND_c_636_n 0.00638651f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A2_c_249_n N_VGND_c_637_n 2.31083e-19 $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A2_c_250_n N_VGND_c_637_n 0.0048389f $X=5.36 $Y=0.995 $X2=0 $Y2=0
cc_248 A2 N_VGND_c_637_n 0.0143134f $X=5.64 $Y=1.105 $X2=0 $Y2=0
cc_249 N_A2_c_248_n N_VGND_c_640_n 0.00395199f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A2_c_250_n N_VGND_c_640_n 0.00585385f $X=5.36 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A2_c_248_n N_VGND_c_643_n 0.00596736f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A2_c_250_n N_VGND_c_643_n 0.0117528f $X=5.36 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A2_c_248_n N_A_805_47#_c_721_n 0.00525851f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A2_c_249_n N_A_805_47#_c_720_n 0.00236971f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A2_c_258_n N_A_805_47#_c_720_n 0.00314708f $X=5.1 $Y=1.53 $X2=0 $Y2=0
cc_256 N_A2_c_253_n N_A_805_47#_c_720_n 0.0146598f $X=5.27 $Y=1.175 $X2=0 $Y2=0
cc_257 N_A1_c_324_n N_Y_c_435_n 0.00303345f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A1_c_325_n N_Y_c_435_n 2.04167e-19 $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A1_c_327_n N_Y_c_435_n 0.0047334f $X=4.865 $Y=1.202 $X2=0 $Y2=0
cc_260 N_A1_c_324_n N_Y_c_436_n 0.00762805f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_261 A1 N_Y_c_436_n 0.0411731f $X=4.725 $Y=1.105 $X2=0 $Y2=0
cc_262 N_A1_c_328_n N_A_321_297#_c_517_n 0.011229f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A1_c_329_n N_A_321_297#_c_520_n 0.011229f $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A1_c_328_n N_VPWR_c_566_n 0.00300743f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A1_c_329_n N_VPWR_c_567_n 0.00300743f $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A1_c_328_n N_VPWR_c_570_n 0.00702461f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A1_c_329_n N_VPWR_c_570_n 0.00702461f $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A1_c_328_n N_VPWR_c_565_n 0.00695979f $X=4.395 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A1_c_329_n N_VPWR_c_565_n 0.00695979f $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A1_c_324_n N_VGND_c_640_n 0.00357877f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A1_c_325_n N_VGND_c_640_n 0.00357877f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A1_c_324_n N_VGND_c_643_n 0.005504f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A1_c_325_n N_VGND_c_643_n 0.00562222f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A1_c_324_n N_A_805_47#_c_721_n 0.0100245f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A1_c_325_n N_A_805_47#_c_721_n 0.0125801f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_276 A1 N_A_805_47#_c_721_n 0.00271194f $X=4.725 $Y=1.105 $X2=0 $Y2=0
cc_277 N_A_27_297#_c_370_n N_Y_M1004_d 0.00352392f $X=1.125 $Y=2.38 $X2=0 $Y2=0
cc_278 N_A_27_297#_c_372_n N_Y_c_433_n 0.00842946f $X=1.21 $Y=1.66 $X2=0 $Y2=0
cc_279 N_A_27_297#_c_370_n Y 0.0147284f $X=1.125 $Y=2.38 $X2=0 $Y2=0
cc_280 N_A_27_297#_c_372_n Y 0.0179146f $X=1.21 $Y=1.66 $X2=0 $Y2=0
cc_281 N_A_27_297#_c_373_n Y 0.0104885f $X=1.25 $Y=2.295 $X2=0 $Y2=0
cc_282 N_A_27_297#_c_375_n Y 0.0114322f $X=1.25 $Y=1.87 $X2=0 $Y2=0
cc_283 N_A_27_297#_c_374_n N_A_321_297#_M1008_s 0.00876152f $X=2.075 $Y=1.87
+ $X2=-0.19 $Y2=1.305
cc_284 N_A_27_297#_c_395_n N_A_321_297#_M1001_s 0.00347905f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_285 N_A_27_297#_M1008_d N_A_321_297#_c_509_n 0.0035039f $X=2.055 $Y=1.485
+ $X2=0 $Y2=0
cc_286 N_A_27_297#_c_374_n N_A_321_297#_c_509_n 0.00608347f $X=2.075 $Y=1.87
+ $X2=0 $Y2=0
cc_287 N_A_27_297#_c_395_n N_A_321_297#_c_509_n 0.00608347f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_288 N_A_27_297#_c_396_n N_A_321_297#_c_509_n 0.0126551f $X=2.2 $Y=1.87 $X2=0
+ $Y2=0
cc_289 N_A_27_297#_M1005_d N_A_321_297#_c_510_n 0.0035039f $X=2.995 $Y=1.485
+ $X2=0 $Y2=0
cc_290 N_A_27_297#_c_395_n N_A_321_297#_c_510_n 0.00608347f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_291 N_A_27_297#_c_398_n N_A_321_297#_c_510_n 0.0126551f $X=3.14 $Y=1.87 $X2=0
+ $Y2=0
cc_292 N_A_27_297#_c_370_n N_A_321_297#_c_538_n 0.011663f $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_293 N_A_27_297#_c_373_n N_A_321_297#_c_538_n 0.0106948f $X=1.25 $Y=2.295
+ $X2=0 $Y2=0
cc_294 N_A_27_297#_c_374_n N_A_321_297#_c_538_n 0.0158267f $X=2.075 $Y=1.87
+ $X2=0 $Y2=0
cc_295 N_A_27_297#_c_395_n N_A_321_297#_c_541_n 0.0131392f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_296 N_A_27_297#_c_370_n N_VPWR_c_568_n 0.0557918f $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_297 N_A_27_297#_c_371_n N_VPWR_c_568_n 0.022203f $X=0.435 $Y=2.38 $X2=0 $Y2=0
cc_298 N_A_27_297#_M1004_s N_VPWR_c_565_n 0.00225715f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_299 N_A_27_297#_M1018_s N_VPWR_c_565_n 0.00217523f $X=1.065 $Y=1.485 $X2=0
+ $Y2=0
cc_300 N_A_27_297#_M1008_d N_VPWR_c_565_n 0.00231289f $X=2.055 $Y=1.485 $X2=0
+ $Y2=0
cc_301 N_A_27_297#_M1005_d N_VPWR_c_565_n 0.00232092f $X=2.995 $Y=1.485 $X2=0
+ $Y2=0
cc_302 N_A_27_297#_c_370_n N_VPWR_c_565_n 0.0336958f $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_303 N_A_27_297#_c_371_n N_VPWR_c_565_n 0.0131123f $X=0.435 $Y=2.38 $X2=0
+ $Y2=0
cc_304 N_A_27_297#_c_374_n N_VPWR_c_565_n 0.00942151f $X=2.075 $Y=1.87 $X2=0
+ $Y2=0
cc_305 N_A_27_297#_c_395_n N_VPWR_c_565_n 0.00153883f $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_306 N_Y_M1004_d N_VPWR_c_565_n 0.00232895f $X=0.595 $Y=1.485 $X2=0 $Y2=0
cc_307 N_Y_c_433_n N_VGND_M1016_d 0.0121649f $X=2.435 $Y=0.775 $X2=0 $Y2=0
cc_308 N_Y_c_436_n N_VGND_M1017_d 0.00432921f $X=4.415 $Y=0.775 $X2=0 $Y2=0
cc_309 Y N_VGND_c_635_n 0.0132149f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_310 N_Y_c_446_n N_VGND_c_635_n 0.0322239f $X=0.74 $Y=0.39 $X2=0 $Y2=0
cc_311 N_Y_c_436_n N_VGND_c_636_n 0.0131987f $X=4.415 $Y=0.775 $X2=0 $Y2=0
cc_312 N_Y_c_433_n N_VGND_c_638_n 0.00200011f $X=2.435 $Y=0.775 $X2=0 $Y2=0
cc_313 N_Y_c_436_n N_VGND_c_638_n 0.00315761f $X=4.415 $Y=0.775 $X2=0 $Y2=0
cc_314 N_Y_c_436_n N_VGND_c_640_n 0.00250893f $X=4.415 $Y=0.775 $X2=0 $Y2=0
cc_315 N_Y_M1007_s N_VGND_c_643_n 0.00267672f $X=0.605 $Y=0.235 $X2=0 $Y2=0
cc_316 N_Y_M1000_d N_VGND_c_643_n 0.00297142f $X=2.485 $Y=0.235 $X2=0 $Y2=0
cc_317 N_Y_M1006_d N_VGND_c_643_n 0.00297142f $X=4.445 $Y=0.235 $X2=0 $Y2=0
cc_318 N_Y_c_433_n N_VGND_c_643_n 0.0127285f $X=2.435 $Y=0.775 $X2=0 $Y2=0
cc_319 N_Y_c_436_n N_VGND_c_643_n 0.0140963f $X=4.415 $Y=0.775 $X2=0 $Y2=0
cc_320 N_Y_c_446_n N_VGND_c_643_n 0.0137337f $X=0.74 $Y=0.39 $X2=0 $Y2=0
cc_321 N_Y_c_433_n N_VGND_c_644_n 0.00254521f $X=2.435 $Y=0.775 $X2=0 $Y2=0
cc_322 N_Y_c_446_n N_VGND_c_644_n 0.0174746f $X=0.74 $Y=0.39 $X2=0 $Y2=0
cc_323 N_Y_c_433_n N_VGND_c_645_n 0.0533815f $X=2.435 $Y=0.775 $X2=0 $Y2=0
cc_324 N_Y_c_433_n N_A_413_47#_M1010_s 0.00191752f $X=2.435 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_325 N_Y_c_436_n N_A_413_47#_M1011_s 0.00253211f $X=4.415 $Y=0.775 $X2=0 $Y2=0
cc_326 N_Y_M1000_d N_A_413_47#_c_706_n 0.00507817f $X=2.485 $Y=0.235 $X2=0 $Y2=0
cc_327 N_Y_c_432_n N_A_413_47#_c_706_n 0.0218848f $X=2.565 $Y=0.775 $X2=0 $Y2=0
cc_328 N_Y_c_433_n N_A_413_47#_c_706_n 0.0163438f $X=2.435 $Y=0.775 $X2=0 $Y2=0
cc_329 N_Y_c_436_n N_A_413_47#_c_706_n 0.017531f $X=4.415 $Y=0.775 $X2=0 $Y2=0
cc_330 N_Y_c_436_n N_A_805_47#_M1003_d 0.00191752f $X=4.415 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_331 N_Y_M1006_d N_A_805_47#_c_721_n 0.00507817f $X=4.445 $Y=0.235 $X2=0 $Y2=0
cc_332 N_Y_c_435_n N_A_805_47#_c_721_n 0.0205972f $X=4.63 $Y=0.73 $X2=0 $Y2=0
cc_333 N_Y_c_436_n N_A_805_47#_c_721_n 0.0172789f $X=4.415 $Y=0.775 $X2=0 $Y2=0
cc_334 N_Y_c_435_n N_A_805_47#_c_720_n 0.00130066f $X=4.63 $Y=0.73 $X2=0 $Y2=0
cc_335 N_A_321_297#_c_517_n N_VPWR_M1002_d 0.00369247f $X=4.505 $Y=1.87
+ $X2=-0.19 $Y2=1.305
cc_336 N_A_321_297#_c_520_n N_VPWR_M1015_d 0.00369025f $X=5.49 $Y=1.87 $X2=0
+ $Y2=0
cc_337 N_A_321_297#_c_517_n N_VPWR_c_566_n 0.0139109f $X=4.505 $Y=1.87 $X2=0
+ $Y2=0
cc_338 N_A_321_297#_c_520_n N_VPWR_c_567_n 0.0139109f $X=5.49 $Y=1.87 $X2=0
+ $Y2=0
cc_339 N_A_321_297#_c_509_n N_VPWR_c_568_n 0.0386534f $X=2.545 $Y=2.38 $X2=0
+ $Y2=0
cc_340 N_A_321_297#_c_510_n N_VPWR_c_568_n 0.0576444f $X=3.525 $Y=2.38 $X2=0
+ $Y2=0
cc_341 N_A_321_297#_c_538_n N_VPWR_c_568_n 0.0154637f $X=1.73 $Y=2.3 $X2=0 $Y2=0
cc_342 N_A_321_297#_c_541_n N_VPWR_c_568_n 0.014332f $X=2.67 $Y=2.3 $X2=0 $Y2=0
cc_343 N_A_321_297#_c_550_p N_VPWR_c_570_n 0.0149311f $X=4.63 $Y=1.96 $X2=0
+ $Y2=0
cc_344 N_A_321_297#_c_551_p N_VPWR_c_572_n 0.0142751f $X=5.575 $Y=1.96 $X2=0
+ $Y2=0
cc_345 N_A_321_297#_M1008_s N_VPWR_c_565_n 0.00215913f $X=1.605 $Y=1.485 $X2=0
+ $Y2=0
cc_346 N_A_321_297#_M1001_s N_VPWR_c_565_n 0.00229658f $X=2.525 $Y=1.485 $X2=0
+ $Y2=0
cc_347 N_A_321_297#_M1019_s N_VPWR_c_565_n 0.00328363f $X=3.465 $Y=1.485 $X2=0
+ $Y2=0
cc_348 N_A_321_297#_M1013_s N_VPWR_c_565_n 0.00250817f $X=4.485 $Y=1.485 $X2=0
+ $Y2=0
cc_349 N_A_321_297#_M1009_s N_VPWR_c_565_n 0.00363111f $X=5.425 $Y=1.485 $X2=0
+ $Y2=0
cc_350 N_A_321_297#_c_509_n N_VPWR_c_565_n 0.0239144f $X=2.545 $Y=2.38 $X2=0
+ $Y2=0
cc_351 N_A_321_297#_c_510_n N_VPWR_c_565_n 0.0350242f $X=3.525 $Y=2.38 $X2=0
+ $Y2=0
cc_352 N_A_321_297#_c_517_n N_VPWR_c_565_n 0.0155943f $X=4.505 $Y=1.87 $X2=0
+ $Y2=0
cc_353 N_A_321_297#_c_550_p N_VPWR_c_565_n 0.00955092f $X=4.63 $Y=1.96 $X2=0
+ $Y2=0
cc_354 N_A_321_297#_c_520_n N_VPWR_c_565_n 0.0158107f $X=5.49 $Y=1.87 $X2=0
+ $Y2=0
cc_355 N_A_321_297#_c_551_p N_VPWR_c_565_n 0.00781789f $X=5.575 $Y=1.96 $X2=0
+ $Y2=0
cc_356 N_A_321_297#_c_538_n N_VPWR_c_565_n 0.00938745f $X=1.73 $Y=2.3 $X2=0
+ $Y2=0
cc_357 N_A_321_297#_c_541_n N_VPWR_c_565_n 0.00938745f $X=2.67 $Y=2.3 $X2=0
+ $Y2=0
cc_358 N_VGND_c_643_n N_A_413_47#_M1010_s 0.00215227f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_359 N_VGND_c_643_n N_A_413_47#_M1011_s 0.00264825f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_638_n N_A_413_47#_c_706_n 0.0749156f $X=3.57 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_643_n N_A_413_47#_c_706_n 0.0474961f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_362 N_VGND_c_645_n N_A_413_47#_c_706_n 0.0190752f $X=1.815 $Y=0.235 $X2=0
+ $Y2=0
cc_363 N_VGND_c_643_n N_A_805_47#_M1003_d 0.00215227f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_364 N_VGND_c_643_n N_A_805_47#_M1014_s 0.00321315f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_636_n N_A_805_47#_c_721_n 0.0148152f $X=3.655 $Y=0.39 $X2=0
+ $Y2=0
cc_366 N_VGND_c_640_n N_A_805_47#_c_721_n 0.0600765f $X=5.485 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_643_n N_A_805_47#_c_721_n 0.0381287f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_640_n N_A_805_47#_c_738_n 0.0159994f $X=5.485 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_643_n N_A_805_47#_c_738_n 0.00961661f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_637_n N_A_805_47#_c_720_n 0.00122902f $X=5.57 $Y=0.39 $X2=0
+ $Y2=0
