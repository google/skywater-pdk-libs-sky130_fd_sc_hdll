# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hdll__muxb
  CLASS BLOCK ;
  FOREIGN sky130_fd_sc_hdll__muxb ;
  ORIGIN  0.190000  0.240000 ;
  SIZE  225.7800 BY  5.920000 ;
  OBS
    LAYER li1 ;
      RECT   0.000000 -0.085000 225.400000 0.085000 ;
      RECT   0.000000  2.635000 107.835000 2.805000 ;
      RECT   0.090000  0.255000   0.345000 1.495000 ;
      RECT   0.090000  1.495000   0.425000 2.465000 ;
      RECT   0.515000  0.085000   0.895000 0.485000 ;
      RECT   0.515000  0.655000   1.610000 0.825000 ;
      RECT   0.515000  0.825000   0.685000 1.325000 ;
      RECT   0.645000  1.495000   0.815000 2.635000 ;
      RECT   0.995000  0.995000   1.270000 1.325000 ;
      RECT   1.070000  1.325000   1.270000 2.295000 ;
      RECT   1.070000  2.295000   3.415000 2.465000 ;
      RECT   1.435000  0.255000   1.955000 0.620000 ;
      RECT   1.435000  0.620000   1.610000 0.655000 ;
      RECT   1.440000  0.825000   1.610000 1.955000 ;
      RECT   1.440000  1.955000   2.885000 2.125000 ;
      RECT   1.780000  0.810000   1.950000 1.615000 ;
      RECT   1.780000  1.615000   3.075000 1.785000 ;
      RECT   2.290000  0.255000   2.615000 1.415000 ;
      RECT   2.785000  0.255000   3.075000 1.615000 ;
      RECT   3.245000  1.440000   3.995000 1.630000 ;
      RECT   3.245000  1.630000   3.415000 2.295000 ;
      RECT   3.250000  0.085000   3.765000 0.525000 ;
      RECT   3.325000  0.695000   4.385000 0.865000 ;
      RECT   3.325000  0.865000   3.495000 1.185000 ;
      RECT   3.585000  1.835000   3.815000 2.635000 ;
      RECT   3.805000  1.055000   3.995000 1.440000 ;
      RECT   3.985000  1.835000   4.385000 2.465000 ;
      RECT   4.035000  0.255000   4.280000 0.695000 ;
      RECT   4.215000  0.865000   4.385000 1.835000 ;
      RECT   4.735000  0.085000   4.985000 0.655000 ;
      RECT   4.735000  1.495000   4.980000 2.635000 ;
      RECT   5.155000  0.255000   5.405000 1.495000 ;
      RECT   5.155000  1.495000   5.495000 2.465000 ;
      RECT   5.575000  0.085000   5.955000 0.485000 ;
      RECT   5.575000  0.655000   6.670000 0.825000 ;
      RECT   5.575000  0.825000   5.745000 1.325000 ;
      RECT   5.675000  1.495000   5.925000 2.635000 ;
      RECT   6.055000  0.995000   6.330000 1.325000 ;
      RECT   6.130000  1.325000   6.330000 2.295000 ;
      RECT   6.130000  2.295000   8.475000 2.465000 ;
      RECT   6.495000  0.255000   7.180000 0.620000 ;
      RECT   6.495000  0.620000   6.670000 0.655000 ;
      RECT   6.500000  0.825000   6.670000 1.955000 ;
      RECT   6.500000  1.955000   7.945000 2.125000 ;
      RECT   6.840000  0.810000   7.010000 1.615000 ;
      RECT   6.840000  1.615000   8.135000 1.785000 ;
      RECT   7.350000  0.255000   7.675000 1.415000 ;
      RECT   7.845000  0.255000   8.135000 1.615000 ;
      RECT   8.305000  1.440000   9.055000 1.630000 ;
      RECT   8.305000  1.630000   8.475000 2.295000 ;
      RECT   8.310000  0.085000   8.825000 0.525000 ;
      RECT   8.385000  0.695000   9.445000 0.865000 ;
      RECT   8.385000  0.865000   8.555000 1.185000 ;
      RECT   8.645000  1.835000   8.875000 2.635000 ;
      RECT   8.865000  1.055000   9.055000 1.440000 ;
      RECT   9.045000  1.835000   9.445000 2.465000 ;
      RECT   9.095000  0.255000   9.340000 0.695000 ;
      RECT   9.275000  0.865000   9.445000 1.835000 ;
      RECT   9.795000  1.495000  10.055000 2.635000 ;
      RECT   9.835000  0.085000  10.080000 0.655000 ;
      RECT  10.225000  1.495000  10.555000 2.465000 ;
      RECT  10.250000  0.255000  10.510000 1.065000 ;
      RECT  10.250000  1.065000  11.405000 1.325000 ;
      RECT  10.250000  1.325000  10.510000 1.495000 ;
      RECT  10.715000  0.085000  10.965000 0.655000 ;
      RECT  10.725000  1.495000  10.965000 2.635000 ;
      RECT  11.135000  0.255000  11.405000 1.065000 ;
      RECT  11.135000  1.325000  11.405000 1.495000 ;
      RECT  11.135000  1.495000  11.495000 2.465000 ;
      RECT  11.575000  0.085000  11.935000 0.485000 ;
      RECT  11.575000  0.655000  12.650000 0.825000 ;
      RECT  11.575000  0.825000  11.745000 1.325000 ;
      RECT  11.665000  1.495000  11.940000 2.635000 ;
      RECT  12.035000  0.995000  12.310000 1.325000 ;
      RECT  12.110000  1.325000  12.310000 2.295000 ;
      RECT  12.110000  2.295000  14.455000 2.465000 ;
      RECT  12.475000  0.255000  13.160000 0.620000 ;
      RECT  12.475000  0.620000  12.650000 0.655000 ;
      RECT  12.480000  0.825000  12.650000 1.955000 ;
      RECT  12.480000  1.955000  13.925000 2.125000 ;
      RECT  12.820000  0.810000  12.990000 1.615000 ;
      RECT  12.820000  1.615000  14.115000 1.785000 ;
      RECT  13.330000  0.255000  13.655000 1.415000 ;
      RECT  13.825000  0.255000  14.115000 1.615000 ;
      RECT  14.285000  1.440000  15.035000 1.630000 ;
      RECT  14.285000  1.630000  14.455000 2.295000 ;
      RECT  14.290000  0.085000  14.805000 0.525000 ;
      RECT  14.365000  0.695000  15.425000 0.865000 ;
      RECT  14.365000  0.865000  14.535000 1.185000 ;
      RECT  14.625000  1.835000  14.855000 2.635000 ;
      RECT  14.845000  1.055000  15.035000 1.440000 ;
      RECT  15.025000  1.835000  15.425000 2.465000 ;
      RECT  15.075000  0.255000  15.320000 0.695000 ;
      RECT  15.255000  0.865000  15.425000 1.835000 ;
      RECT  15.735000  1.495000  16.065000 2.635000 ;
      RECT  15.770000  0.085000  16.030000 0.885000 ;
      RECT  15.975000  1.055000  16.370000 1.325000 ;
      RECT  16.200000  0.395000  16.475000 0.625000 ;
      RECT  16.200000  0.625000  16.370000 1.055000 ;
      RECT  16.540000  0.835000  16.930000 1.005000 ;
      RECT  16.540000  1.005000  16.710000 1.755000 ;
      RECT  16.540000  1.755000  16.935000 1.805000 ;
      RECT  16.540000  1.805000  17.060000 1.985000 ;
      RECT  16.685000  0.330000  16.930000 0.835000 ;
      RECT  16.730000  1.985000  17.060000 2.465000 ;
      RECT  16.880000  1.175000  17.270000 1.465000 ;
      RECT  16.880000  1.465000  17.580000 1.505000 ;
      RECT  17.100000  0.585000  17.540000 0.755000 ;
      RECT  17.100000  0.755000  17.270000 1.175000 ;
      RECT  17.100000  1.505000  17.580000 1.635000 ;
      RECT  17.250000  1.635000  17.580000 2.465000 ;
      RECT  17.290000  0.330000  17.540000 0.585000 ;
      RECT  17.445000  0.945000  17.795000 1.295000 ;
      RECT  17.775000  0.085000  18.105000 0.660000 ;
      RECT  17.805000  1.465000  18.105000 2.635000 ;
      RECT  18.085000  0.945000  18.435000 1.295000 ;
      RECT  18.300000  1.465000  19.000000 1.505000 ;
      RECT  18.300000  1.505000  18.780000 1.635000 ;
      RECT  18.300000  1.635000  18.630000 2.465000 ;
      RECT  18.340000  0.330000  18.590000 0.585000 ;
      RECT  18.340000  0.585000  18.780000 0.755000 ;
      RECT  18.610000  0.755000  18.780000 1.175000 ;
      RECT  18.610000  1.175000  19.000000 1.465000 ;
      RECT  18.820000  1.805000  19.340000 1.985000 ;
      RECT  18.820000  1.985000  19.150000 2.465000 ;
      RECT  18.945000  1.755000  19.340000 1.805000 ;
      RECT  18.950000  0.330000  19.195000 0.835000 ;
      RECT  18.950000  0.835000  19.340000 1.005000 ;
      RECT  19.170000  1.005000  19.340000 1.755000 ;
      RECT  19.405000  0.395000  19.680000 0.625000 ;
      RECT  19.510000  0.625000  19.680000 1.055000 ;
      RECT  19.510000  1.055000  19.905000 1.325000 ;
      RECT  19.815000  1.495000  20.205000 2.635000 ;
      RECT  19.850000  0.085000  20.170000 0.885000 ;
      RECT  20.115000  1.055000  20.510000 1.325000 ;
      RECT  20.340000  0.395000  20.615000 0.625000 ;
      RECT  20.340000  0.625000  20.510000 1.055000 ;
      RECT  20.680000  0.835000  21.070000 1.005000 ;
      RECT  20.680000  1.005000  20.850000 1.755000 ;
      RECT  20.680000  1.755000  21.075000 1.805000 ;
      RECT  20.680000  1.805000  21.200000 1.985000 ;
      RECT  20.825000  0.330000  21.070000 0.835000 ;
      RECT  20.870000  1.985000  21.200000 2.465000 ;
      RECT  21.020000  1.175000  21.410000 1.465000 ;
      RECT  21.020000  1.465000  21.720000 1.505000 ;
      RECT  21.240000  0.585000  21.680000 0.755000 ;
      RECT  21.240000  0.755000  21.410000 1.175000 ;
      RECT  21.240000  1.505000  21.720000 1.635000 ;
      RECT  21.390000  1.635000  21.720000 2.465000 ;
      RECT  21.430000  0.330000  21.680000 0.585000 ;
      RECT  21.585000  0.945000  21.935000 1.295000 ;
      RECT  21.915000  0.085000  22.245000 0.660000 ;
      RECT  21.915000  1.465000  22.215000 2.635000 ;
      RECT  22.225000  0.945000  22.575000 1.295000 ;
      RECT  22.440000  1.465000  23.140000 1.505000 ;
      RECT  22.440000  1.505000  22.920000 1.635000 ;
      RECT  22.440000  1.635000  22.770000 2.465000 ;
      RECT  22.480000  0.330000  22.730000 0.585000 ;
      RECT  22.480000  0.585000  22.920000 0.755000 ;
      RECT  22.750000  0.755000  22.920000 1.175000 ;
      RECT  22.750000  1.175000  23.140000 1.465000 ;
      RECT  22.960000  1.805000  23.480000 1.985000 ;
      RECT  22.960000  1.985000  23.290000 2.465000 ;
      RECT  23.085000  1.755000  23.480000 1.805000 ;
      RECT  23.090000  0.330000  23.335000 0.835000 ;
      RECT  23.090000  0.835000  23.480000 1.005000 ;
      RECT  23.310000  1.005000  23.480000 1.755000 ;
      RECT  23.545000  0.395000  23.820000 0.625000 ;
      RECT  23.650000  0.625000  23.820000 1.055000 ;
      RECT  23.650000  1.055000  24.045000 1.325000 ;
      RECT  23.955000  1.495000  24.285000 2.635000 ;
      RECT  23.990000  0.085000  24.250000 0.885000 ;
      RECT  24.475000  1.055000  25.295000 1.325000 ;
      RECT  24.475000  1.495000  25.665000 1.665000 ;
      RECT  24.475000  1.665000  24.775000 2.210000 ;
      RECT  24.475000  2.210000  24.805000 2.465000 ;
      RECT  24.525000  0.255000  24.855000 0.715000 ;
      RECT  24.525000  0.715000  25.715000 0.885000 ;
      RECT  24.945000  1.835000  25.275000 2.105000 ;
      RECT  24.975000  2.105000  25.275000 2.635000 ;
      RECT  25.025000  0.085000  25.240000 0.545000 ;
      RECT  25.410000  0.255000  26.555000 0.425000 ;
      RECT  25.410000  0.425000  25.715000 0.715000 ;
      RECT  25.410000  0.885000  25.715000 0.925000 ;
      RECT  25.495000  1.665000  25.665000 2.295000 ;
      RECT  25.495000  2.295000  26.660000 2.465000 ;
      RECT  25.845000  1.755000  26.275000 2.125000 ;
      RECT  25.885000  0.595000  26.215000 0.885000 ;
      RECT  25.965000  0.885000  26.135000 1.755000 ;
      RECT  26.385000  0.425000  26.555000 0.770000 ;
      RECT  26.480000  1.205000  26.895000 1.305000 ;
      RECT  26.480000  1.305000  27.000000 1.465000 ;
      RECT  26.480000  1.465000  27.260000 1.475000 ;
      RECT  26.490000  1.645000  26.660000 2.295000 ;
      RECT  26.725000  0.585000  27.305000 0.755000 ;
      RECT  26.725000  0.755000  26.895000 1.205000 ;
      RECT  26.830000  1.475000  27.260000 1.635000 ;
      RECT  26.930000  1.635000  27.260000 2.465000 ;
      RECT  27.055000  0.330000  27.305000 0.585000 ;
      RECT  27.170000  1.025000  27.505000 1.295000 ;
      RECT  27.435000  1.465000  27.765000 2.635000 ;
      RECT  27.475000  0.085000  27.725000 0.660000 ;
      RECT  27.695000  1.025000  28.030000 1.295000 ;
      RECT  27.895000  0.330000  28.145000 0.585000 ;
      RECT  27.895000  0.585000  28.475000 0.755000 ;
      RECT  27.940000  1.465000  28.720000 1.475000 ;
      RECT  27.940000  1.475000  28.370000 1.635000 ;
      RECT  27.940000  1.635000  28.270000 2.465000 ;
      RECT  28.200000  1.305000  28.720000 1.465000 ;
      RECT  28.305000  0.755000  28.475000 1.205000 ;
      RECT  28.305000  1.205000  28.720000 1.305000 ;
      RECT  28.540000  1.645000  28.710000 2.295000 ;
      RECT  28.540000  2.295000  29.705000 2.465000 ;
      RECT  28.645000  0.255000  29.790000 0.425000 ;
      RECT  28.645000  0.425000  28.815000 0.770000 ;
      RECT  28.925000  1.755000  29.355000 2.125000 ;
      RECT  28.985000  0.595000  29.315000 0.885000 ;
      RECT  29.065000  0.885000  29.235000 1.755000 ;
      RECT  29.485000  0.425000  29.790000 0.715000 ;
      RECT  29.485000  0.715000  30.675000 0.885000 ;
      RECT  29.485000  0.885000  29.790000 0.925000 ;
      RECT  29.535000  1.495000  30.725000 1.665000 ;
      RECT  29.535000  1.665000  29.705000 2.295000 ;
      RECT  29.905000  1.055000  30.725000 1.325000 ;
      RECT  29.925000  1.835000  30.255000 2.105000 ;
      RECT  29.925000  2.105000  30.225000 2.635000 ;
      RECT  29.960000  0.085000  30.175000 0.545000 ;
      RECT  30.345000  0.255000  30.675000 0.715000 ;
      RECT  30.395000  2.210000  30.725000 2.465000 ;
      RECT  30.425000  1.665000  30.725000 2.210000 ;
      RECT  30.915000  1.055000  31.735000 1.325000 ;
      RECT  30.915000  1.495000  32.105000 1.665000 ;
      RECT  30.915000  1.665000  31.215000 2.210000 ;
      RECT  30.915000  2.210000  31.245000 2.465000 ;
      RECT  30.965000  0.255000  31.295000 0.715000 ;
      RECT  30.965000  0.715000  32.155000 0.885000 ;
      RECT  31.385000  1.835000  31.715000 2.105000 ;
      RECT  31.415000  2.105000  31.715000 2.635000 ;
      RECT  31.465000  0.085000  31.680000 0.545000 ;
      RECT  31.850000  0.255000  32.995000 0.425000 ;
      RECT  31.850000  0.425000  32.155000 0.715000 ;
      RECT  31.850000  0.885000  32.155000 0.925000 ;
      RECT  31.935000  1.665000  32.105000 2.295000 ;
      RECT  31.935000  2.295000  33.100000 2.465000 ;
      RECT  32.285000  1.755000  32.715000 2.125000 ;
      RECT  32.325000  0.595000  32.655000 0.885000 ;
      RECT  32.405000  0.885000  32.575000 1.755000 ;
      RECT  32.825000  0.425000  32.995000 0.770000 ;
      RECT  32.920000  1.205000  33.335000 1.305000 ;
      RECT  32.920000  1.305000  33.440000 1.465000 ;
      RECT  32.920000  1.465000  33.700000 1.475000 ;
      RECT  32.930000  1.645000  33.100000 2.295000 ;
      RECT  33.165000  0.585000  33.745000 0.755000 ;
      RECT  33.165000  0.755000  33.335000 1.205000 ;
      RECT  33.270000  1.475000  33.700000 1.635000 ;
      RECT  33.370000  1.635000  33.700000 2.465000 ;
      RECT  33.495000  0.330000  33.745000 0.585000 ;
      RECT  33.610000  1.025000  33.945000 1.295000 ;
      RECT  33.875000  1.465000  34.205000 2.635000 ;
      RECT  33.915000  0.085000  34.165000 0.660000 ;
      RECT  34.135000  1.025000  34.470000 1.295000 ;
      RECT  34.335000  0.330000  34.585000 0.585000 ;
      RECT  34.335000  0.585000  34.915000 0.755000 ;
      RECT  34.380000  1.465000  35.160000 1.475000 ;
      RECT  34.380000  1.475000  34.810000 1.635000 ;
      RECT  34.380000  1.635000  34.710000 2.465000 ;
      RECT  34.640000  1.305000  35.160000 1.465000 ;
      RECT  34.745000  0.755000  34.915000 1.205000 ;
      RECT  34.745000  1.205000  35.160000 1.305000 ;
      RECT  34.980000  1.645000  35.150000 2.295000 ;
      RECT  34.980000  2.295000  36.145000 2.465000 ;
      RECT  35.085000  0.255000  36.230000 0.425000 ;
      RECT  35.085000  0.425000  35.255000 0.770000 ;
      RECT  35.365000  1.755000  35.795000 2.125000 ;
      RECT  35.425000  0.595000  35.755000 0.885000 ;
      RECT  35.505000  0.885000  35.675000 1.755000 ;
      RECT  35.925000  0.425000  36.230000 0.715000 ;
      RECT  35.925000  0.715000  37.115000 0.885000 ;
      RECT  35.925000  0.885000  36.230000 0.925000 ;
      RECT  35.975000  1.495000  37.165000 1.665000 ;
      RECT  35.975000  1.665000  36.145000 2.295000 ;
      RECT  36.345000  1.055000  37.165000 1.325000 ;
      RECT  36.365000  1.835000  36.695000 2.105000 ;
      RECT  36.365000  2.105000  36.665000 2.635000 ;
      RECT  36.400000  0.085000  36.615000 0.545000 ;
      RECT  36.785000  0.255000  37.115000 0.715000 ;
      RECT  36.835000  2.210000  37.165000 2.465000 ;
      RECT  36.865000  1.665000  37.165000 2.210000 ;
      RECT  37.385000  1.495000  37.655000 2.635000 ;
      RECT  37.405000  0.085000  37.655000 0.885000 ;
      RECT  37.655000  1.055000  39.045000 1.325000 ;
      RECT  37.825000  0.255000  38.155000 0.715000 ;
      RECT  37.825000  0.715000  39.955000 0.885000 ;
      RECT  37.825000  1.495000  40.055000 1.665000 ;
      RECT  37.825000  1.665000  38.155000 2.465000 ;
      RECT  38.325000  0.085000  38.595000 0.545000 ;
      RECT  38.325000  1.835000  38.595000 2.635000 ;
      RECT  38.765000  0.255000  39.095000 0.715000 ;
      RECT  38.765000  1.665000  39.095000 2.465000 ;
      RECT  39.265000  0.085000  39.515000 0.545000 ;
      RECT  39.265000  1.835000  39.535000 2.635000 ;
      RECT  39.685000  0.255000  41.715000 0.425000 ;
      RECT  39.685000  0.425000  39.955000 0.715000 ;
      RECT  39.755000  1.665000  40.055000 2.295000 ;
      RECT  39.755000  2.295000  41.965000 2.465000 ;
      RECT  40.125000  0.595000  40.455000 0.885000 ;
      RECT  40.225000  0.885000  40.455000 1.065000 ;
      RECT  40.225000  1.065000  41.495000 1.365000 ;
      RECT  40.225000  1.365000  40.555000 2.125000 ;
      RECT  40.625000  0.425000  40.795000 0.770000 ;
      RECT  40.725000  1.535000  40.995000 2.295000 ;
      RECT  40.965000  0.595000  41.295000 1.065000 ;
      RECT  41.165000  1.365000  41.495000 2.125000 ;
      RECT  41.465000  0.425000  41.715000 0.770000 ;
      RECT  41.665000  1.065000  42.850000 1.395000 ;
      RECT  41.665000  1.565000  41.965000 2.295000 ;
      RECT  42.210000  1.605000  42.485000 2.635000 ;
      RECT  42.220000  0.085000  42.510000 0.610000 ;
      RECT  42.680000  0.280000  42.930000 0.825000 ;
      RECT  42.680000  0.825000  42.850000 1.065000 ;
      RECT  42.680000  1.395000  42.850000 1.605000 ;
      RECT  42.680000  1.605000  43.010000 2.465000 ;
      RECT  43.020000  0.995000  43.615000 1.325000 ;
      RECT  43.140000  0.085000  43.430000 0.610000 ;
      RECT  43.180000  1.605000  43.480000 2.635000 ;
      RECT  43.785000  0.995000  44.380000 1.325000 ;
      RECT  43.920000  1.605000  44.220000 2.635000 ;
      RECT  43.970000  0.085000  44.260000 0.610000 ;
      RECT  44.390000  1.605000  44.720000 2.465000 ;
      RECT  44.470000  0.280000  44.720000 0.825000 ;
      RECT  44.550000  0.825000  44.720000 1.065000 ;
      RECT  44.550000  1.065000  45.735000 1.395000 ;
      RECT  44.550000  1.395000  44.720000 1.605000 ;
      RECT  44.890000  0.085000  45.180000 0.610000 ;
      RECT  44.915000  1.605000  45.190000 2.635000 ;
      RECT  45.435000  1.565000  45.735000 2.295000 ;
      RECT  45.435000  2.295000  47.645000 2.465000 ;
      RECT  45.685000  0.255000  47.715000 0.425000 ;
      RECT  45.685000  0.425000  45.935000 0.770000 ;
      RECT  45.905000  1.065000  47.175000 1.365000 ;
      RECT  45.905000  1.365000  46.235000 2.125000 ;
      RECT  46.105000  0.595000  46.435000 1.065000 ;
      RECT  46.405000  1.535000  46.675000 2.295000 ;
      RECT  46.605000  0.425000  46.775000 0.770000 ;
      RECT  46.845000  1.365000  47.175000 2.125000 ;
      RECT  46.945000  0.595000  47.275000 0.885000 ;
      RECT  46.945000  0.885000  47.175000 1.065000 ;
      RECT  47.345000  1.495000  49.575000 1.665000 ;
      RECT  47.345000  1.665000  47.645000 2.295000 ;
      RECT  47.445000  0.425000  47.715000 0.715000 ;
      RECT  47.445000  0.715000  49.575000 0.885000 ;
      RECT  47.865000  1.835000  48.135000 2.635000 ;
      RECT  47.885000  0.085000  48.135000 0.545000 ;
      RECT  48.305000  0.255000  48.635000 0.715000 ;
      RECT  48.305000  1.665000  48.635000 2.465000 ;
      RECT  48.355000  1.055000  49.745000 1.325000 ;
      RECT  48.805000  0.085000  49.075000 0.545000 ;
      RECT  48.805000  1.835000  49.075000 2.635000 ;
      RECT  49.245000  0.255000  49.575000 0.715000 ;
      RECT  49.245000  1.665000  49.575000 2.465000 ;
      RECT  49.745000  0.085000  49.995000 0.885000 ;
      RECT  49.745000  1.495000  50.015000 2.635000 ;
      RECT  50.265000  1.495000  50.535000 2.635000 ;
      RECT  50.285000  0.085000  50.535000 0.885000 ;
      RECT  50.535000  1.055000  51.925000 1.325000 ;
      RECT  50.705000  0.255000  51.035000 0.715000 ;
      RECT  50.705000  0.715000  52.835000 0.885000 ;
      RECT  50.705000  1.495000  52.935000 1.665000 ;
      RECT  50.705000  1.665000  51.035000 2.465000 ;
      RECT  51.205000  0.085000  51.475000 0.545000 ;
      RECT  51.205000  1.835000  51.475000 2.635000 ;
      RECT  51.645000  0.255000  51.975000 0.715000 ;
      RECT  51.645000  1.665000  51.975000 2.465000 ;
      RECT  52.145000  0.085000  52.395000 0.545000 ;
      RECT  52.145000  1.835000  52.415000 2.635000 ;
      RECT  52.565000  0.255000  54.595000 0.425000 ;
      RECT  52.565000  0.425000  52.835000 0.715000 ;
      RECT  52.635000  1.665000  52.935000 2.295000 ;
      RECT  52.635000  2.295000  54.845000 2.465000 ;
      RECT  53.005000  0.595000  53.335000 0.885000 ;
      RECT  53.105000  0.885000  53.335000 1.065000 ;
      RECT  53.105000  1.065000  54.375000 1.365000 ;
      RECT  53.105000  1.365000  53.435000 2.125000 ;
      RECT  53.505000  0.425000  53.675000 0.770000 ;
      RECT  53.605000  1.535000  53.875000 2.295000 ;
      RECT  53.845000  0.595000  54.175000 1.065000 ;
      RECT  54.045000  1.365000  54.375000 2.125000 ;
      RECT  54.345000  0.425000  54.595000 0.770000 ;
      RECT  54.545000  1.065000  55.730000 1.395000 ;
      RECT  54.545000  1.565000  54.845000 2.295000 ;
      RECT  55.090000  1.605000  55.365000 2.635000 ;
      RECT  55.100000  0.085000  55.390000 0.610000 ;
      RECT  55.560000  0.280000  55.810000 0.825000 ;
      RECT  55.560000  0.825000  55.730000 1.065000 ;
      RECT  55.560000  1.395000  55.730000 1.605000 ;
      RECT  55.560000  1.605000  55.890000 2.465000 ;
      RECT  55.900000  0.995000  56.495000 1.325000 ;
      RECT  56.020000  0.085000  56.310000 0.610000 ;
      RECT  56.060000  1.605000  56.360000 2.635000 ;
      RECT  56.665000  0.995000  57.260000 1.325000 ;
      RECT  56.800000  1.605000  57.100000 2.635000 ;
      RECT  56.850000  0.085000  57.140000 0.610000 ;
      RECT  57.270000  1.605000  57.600000 2.465000 ;
      RECT  57.350000  0.280000  57.600000 0.825000 ;
      RECT  57.430000  0.825000  57.600000 1.065000 ;
      RECT  57.430000  1.065000  58.615000 1.395000 ;
      RECT  57.430000  1.395000  57.600000 1.605000 ;
      RECT  57.770000  0.085000  58.060000 0.610000 ;
      RECT  57.795000  1.605000  58.070000 2.635000 ;
      RECT  58.315000  1.565000  58.615000 2.295000 ;
      RECT  58.315000  2.295000  60.525000 2.465000 ;
      RECT  58.565000  0.255000  60.595000 0.425000 ;
      RECT  58.565000  0.425000  58.815000 0.770000 ;
      RECT  58.785000  1.065000  60.055000 1.365000 ;
      RECT  58.785000  1.365000  59.115000 2.125000 ;
      RECT  58.985000  0.595000  59.315000 1.065000 ;
      RECT  59.285000  1.535000  59.555000 2.295000 ;
      RECT  59.485000  0.425000  59.655000 0.770000 ;
      RECT  59.725000  1.365000  60.055000 2.125000 ;
      RECT  59.825000  0.595000  60.155000 0.885000 ;
      RECT  59.825000  0.885000  60.055000 1.065000 ;
      RECT  60.225000  1.495000  62.455000 1.665000 ;
      RECT  60.225000  1.665000  60.525000 2.295000 ;
      RECT  60.325000  0.425000  60.595000 0.715000 ;
      RECT  60.325000  0.715000  62.455000 0.885000 ;
      RECT  60.745000  1.835000  61.015000 2.635000 ;
      RECT  60.765000  0.085000  61.015000 0.545000 ;
      RECT  61.185000  0.255000  61.515000 0.715000 ;
      RECT  61.185000  1.665000  61.515000 2.465000 ;
      RECT  61.235000  1.055000  62.625000 1.325000 ;
      RECT  61.685000  0.085000  61.955000 0.545000 ;
      RECT  61.685000  1.835000  61.955000 2.635000 ;
      RECT  62.125000  0.255000  62.455000 0.715000 ;
      RECT  62.125000  1.665000  62.455000 2.465000 ;
      RECT  62.625000  0.085000  62.875000 0.885000 ;
      RECT  62.625000  1.495000  62.895000 2.635000 ;
      RECT  63.115000  1.495000  63.445000 2.635000 ;
      RECT  63.150000  0.085000  63.410000 0.885000 ;
      RECT  63.355000  1.055000  63.750000 1.325000 ;
      RECT  63.580000  0.395000  63.855000 0.625000 ;
      RECT  63.580000  0.625000  63.750000 1.055000 ;
      RECT  63.920000  0.835000  64.310000 1.005000 ;
      RECT  63.920000  1.005000  64.090000 1.755000 ;
      RECT  63.920000  1.755000  64.315000 1.805000 ;
      RECT  63.920000  1.805000  64.440000 1.985000 ;
      RECT  64.065000  0.330000  64.310000 0.835000 ;
      RECT  64.110000  1.985000  64.440000 2.465000 ;
      RECT  64.260000  1.175000  64.650000 1.465000 ;
      RECT  64.260000  1.465000  64.960000 1.505000 ;
      RECT  64.480000  0.585000  64.920000 0.755000 ;
      RECT  64.480000  0.755000  64.650000 1.175000 ;
      RECT  64.480000  1.505000  64.960000 1.635000 ;
      RECT  64.630000  1.635000  64.960000 2.465000 ;
      RECT  64.670000  0.330000  64.920000 0.585000 ;
      RECT  64.825000  0.945000  65.225000 1.295000 ;
      RECT  65.155000  0.085000  65.485000 0.660000 ;
      RECT  65.155000  1.465000  65.485000 2.635000 ;
      RECT  65.415000  0.945000  65.815000 1.295000 ;
      RECT  65.680000  1.465000  66.380000 1.505000 ;
      RECT  65.680000  1.505000  66.160000 1.635000 ;
      RECT  65.680000  1.635000  66.010000 2.465000 ;
      RECT  65.720000  0.330000  65.970000 0.585000 ;
      RECT  65.720000  0.585000  66.160000 0.755000 ;
      RECT  65.990000  0.755000  66.160000 1.175000 ;
      RECT  65.990000  1.175000  66.380000 1.465000 ;
      RECT  66.200000  1.805000  66.720000 1.985000 ;
      RECT  66.200000  1.985000  66.530000 2.465000 ;
      RECT  66.325000  1.755000  66.720000 1.805000 ;
      RECT  66.330000  0.330000  66.575000 0.835000 ;
      RECT  66.330000  0.835000  66.720000 1.005000 ;
      RECT  66.550000  1.005000  66.720000 1.755000 ;
      RECT  66.785000  0.395000  67.060000 0.625000 ;
      RECT  66.890000  0.625000  67.060000 1.055000 ;
      RECT  66.890000  1.055000  67.285000 1.325000 ;
      RECT  67.195000  1.495000  67.585000 2.635000 ;
      RECT  67.230000  0.085000  67.550000 0.885000 ;
      RECT  67.495000  1.055000  67.890000 1.325000 ;
      RECT  67.720000  0.395000  67.995000 0.625000 ;
      RECT  67.720000  0.625000  67.890000 1.055000 ;
      RECT  68.060000  0.835000  68.450000 1.005000 ;
      RECT  68.060000  1.005000  68.230000 1.755000 ;
      RECT  68.060000  1.755000  68.455000 1.805000 ;
      RECT  68.060000  1.805000  68.580000 1.985000 ;
      RECT  68.205000  0.330000  68.450000 0.835000 ;
      RECT  68.250000  1.985000  68.580000 2.465000 ;
      RECT  68.400000  1.175000  68.790000 1.465000 ;
      RECT  68.400000  1.465000  69.100000 1.505000 ;
      RECT  68.620000  0.585000  69.060000 0.755000 ;
      RECT  68.620000  0.755000  68.790000 1.175000 ;
      RECT  68.620000  1.505000  69.100000 1.635000 ;
      RECT  68.770000  1.635000  69.100000 2.465000 ;
      RECT  68.810000  0.330000  69.060000 0.585000 ;
      RECT  68.965000  0.945000  69.365000 1.295000 ;
      RECT  69.295000  0.085000  69.625000 0.660000 ;
      RECT  69.295000  1.465000  69.625000 2.635000 ;
      RECT  69.555000  0.945000  69.955000 1.295000 ;
      RECT  69.820000  1.465000  70.520000 1.505000 ;
      RECT  69.820000  1.505000  70.300000 1.635000 ;
      RECT  69.820000  1.635000  70.150000 2.465000 ;
      RECT  69.860000  0.330000  70.110000 0.585000 ;
      RECT  69.860000  0.585000  70.300000 0.755000 ;
      RECT  70.130000  0.755000  70.300000 1.175000 ;
      RECT  70.130000  1.175000  70.520000 1.465000 ;
      RECT  70.340000  1.805000  70.860000 1.985000 ;
      RECT  70.340000  1.985000  70.670000 2.465000 ;
      RECT  70.465000  1.755000  70.860000 1.805000 ;
      RECT  70.470000  0.330000  70.715000 0.835000 ;
      RECT  70.470000  0.835000  70.860000 1.005000 ;
      RECT  70.690000  1.005000  70.860000 1.755000 ;
      RECT  70.925000  0.395000  71.200000 0.625000 ;
      RECT  71.030000  0.625000  71.200000 1.055000 ;
      RECT  71.030000  1.055000  71.425000 1.325000 ;
      RECT  71.335000  1.495000  71.725000 2.635000 ;
      RECT  71.370000  0.085000  71.690000 0.885000 ;
      RECT  71.635000  1.055000  72.030000 1.325000 ;
      RECT  71.860000  0.395000  72.135000 0.625000 ;
      RECT  71.860000  0.625000  72.030000 1.055000 ;
      RECT  72.200000  0.835000  72.590000 1.005000 ;
      RECT  72.200000  1.005000  72.370000 1.755000 ;
      RECT  72.200000  1.755000  72.595000 1.805000 ;
      RECT  72.200000  1.805000  72.720000 1.985000 ;
      RECT  72.345000  0.330000  72.590000 0.835000 ;
      RECT  72.390000  1.985000  72.720000 2.465000 ;
      RECT  72.540000  1.175000  72.930000 1.465000 ;
      RECT  72.540000  1.465000  73.240000 1.505000 ;
      RECT  72.760000  0.585000  73.200000 0.755000 ;
      RECT  72.760000  0.755000  72.930000 1.175000 ;
      RECT  72.760000  1.505000  73.240000 1.635000 ;
      RECT  72.910000  1.635000  73.240000 2.465000 ;
      RECT  72.950000  0.330000  73.200000 0.585000 ;
      RECT  73.105000  0.945000  73.505000 1.295000 ;
      RECT  73.435000  0.085000  73.765000 0.660000 ;
      RECT  73.435000  1.465000  73.765000 2.635000 ;
      RECT  73.695000  0.945000  74.095000 1.295000 ;
      RECT  73.960000  1.465000  74.660000 1.505000 ;
      RECT  73.960000  1.505000  74.440000 1.635000 ;
      RECT  73.960000  1.635000  74.290000 2.465000 ;
      RECT  74.000000  0.330000  74.250000 0.585000 ;
      RECT  74.000000  0.585000  74.440000 0.755000 ;
      RECT  74.270000  0.755000  74.440000 1.175000 ;
      RECT  74.270000  1.175000  74.660000 1.465000 ;
      RECT  74.480000  1.805000  75.000000 1.985000 ;
      RECT  74.480000  1.985000  74.810000 2.465000 ;
      RECT  74.605000  1.755000  75.000000 1.805000 ;
      RECT  74.610000  0.330000  74.855000 0.835000 ;
      RECT  74.610000  0.835000  75.000000 1.005000 ;
      RECT  74.830000  1.005000  75.000000 1.755000 ;
      RECT  75.065000  0.395000  75.340000 0.625000 ;
      RECT  75.170000  0.625000  75.340000 1.055000 ;
      RECT  75.170000  1.055000  75.565000 1.325000 ;
      RECT  75.475000  1.495000  75.865000 2.635000 ;
      RECT  75.510000  0.085000  75.830000 0.885000 ;
      RECT  75.775000  1.055000  76.170000 1.325000 ;
      RECT  76.000000  0.395000  76.275000 0.625000 ;
      RECT  76.000000  0.625000  76.170000 1.055000 ;
      RECT  76.340000  0.835000  76.730000 1.005000 ;
      RECT  76.340000  1.005000  76.510000 1.755000 ;
      RECT  76.340000  1.755000  76.735000 1.805000 ;
      RECT  76.340000  1.805000  76.860000 1.985000 ;
      RECT  76.485000  0.330000  76.730000 0.835000 ;
      RECT  76.530000  1.985000  76.860000 2.465000 ;
      RECT  76.680000  1.175000  77.070000 1.465000 ;
      RECT  76.680000  1.465000  77.380000 1.505000 ;
      RECT  76.900000  0.585000  77.340000 0.755000 ;
      RECT  76.900000  0.755000  77.070000 1.175000 ;
      RECT  76.900000  1.505000  77.380000 1.635000 ;
      RECT  77.050000  1.635000  77.380000 2.465000 ;
      RECT  77.090000  0.330000  77.340000 0.585000 ;
      RECT  77.245000  0.945000  77.645000 1.295000 ;
      RECT  77.575000  0.085000  77.905000 0.660000 ;
      RECT  77.575000  1.465000  77.905000 2.635000 ;
      RECT  77.835000  0.945000  78.235000 1.295000 ;
      RECT  78.100000  1.465000  78.800000 1.505000 ;
      RECT  78.100000  1.505000  78.580000 1.635000 ;
      RECT  78.100000  1.635000  78.430000 2.465000 ;
      RECT  78.140000  0.330000  78.390000 0.585000 ;
      RECT  78.140000  0.585000  78.580000 0.755000 ;
      RECT  78.410000  0.755000  78.580000 1.175000 ;
      RECT  78.410000  1.175000  78.800000 1.465000 ;
      RECT  78.620000  1.805000  79.140000 1.985000 ;
      RECT  78.620000  1.985000  78.950000 2.465000 ;
      RECT  78.745000  1.755000  79.140000 1.805000 ;
      RECT  78.750000  0.330000  78.995000 0.835000 ;
      RECT  78.750000  0.835000  79.140000 1.005000 ;
      RECT  78.970000  1.005000  79.140000 1.755000 ;
      RECT  79.205000  0.395000  79.480000 0.625000 ;
      RECT  79.310000  0.625000  79.480000 1.055000 ;
      RECT  79.310000  1.055000  79.705000 1.325000 ;
      RECT  79.615000  1.495000  79.945000 2.635000 ;
      RECT  79.650000  0.085000  79.910000 0.885000 ;
      RECT  80.135000  1.055000  80.955000 1.325000 ;
      RECT  80.135000  1.495000  81.325000 1.665000 ;
      RECT  80.135000  1.665000  80.435000 2.210000 ;
      RECT  80.135000  2.210000  80.465000 2.465000 ;
      RECT  80.185000  0.255000  80.515000 0.715000 ;
      RECT  80.185000  0.715000  81.375000 0.885000 ;
      RECT  80.605000  1.835000  80.935000 2.105000 ;
      RECT  80.635000  2.105000  80.935000 2.635000 ;
      RECT  80.685000  0.085000  80.900000 0.545000 ;
      RECT  81.070000  0.255000  82.215000 0.425000 ;
      RECT  81.070000  0.425000  81.375000 0.715000 ;
      RECT  81.070000  0.885000  81.375000 0.925000 ;
      RECT  81.155000  1.665000  81.325000 2.295000 ;
      RECT  81.155000  2.295000  82.320000 2.465000 ;
      RECT  81.505000  1.755000  81.935000 2.125000 ;
      RECT  81.545000  0.595000  81.875000 0.885000 ;
      RECT  81.625000  0.885000  81.795000 1.755000 ;
      RECT  82.045000  0.425000  82.215000 0.770000 ;
      RECT  82.140000  1.205000  82.555000 1.305000 ;
      RECT  82.140000  1.305000  82.660000 1.465000 ;
      RECT  82.140000  1.465000  82.920000 1.475000 ;
      RECT  82.150000  1.645000  82.320000 2.295000 ;
      RECT  82.385000  0.585000  82.965000 0.755000 ;
      RECT  82.385000  0.755000  82.555000 1.205000 ;
      RECT  82.490000  1.475000  82.920000 1.635000 ;
      RECT  82.590000  1.635000  82.920000 2.465000 ;
      RECT  82.715000  0.330000  82.965000 0.585000 ;
      RECT  82.830000  1.025000  83.165000 1.295000 ;
      RECT  83.095000  1.465000  83.425000 2.635000 ;
      RECT  83.135000  0.085000  83.385000 0.660000 ;
      RECT  83.355000  1.025000  83.690000 1.295000 ;
      RECT  83.555000  0.330000  83.805000 0.585000 ;
      RECT  83.555000  0.585000  84.135000 0.755000 ;
      RECT  83.600000  1.465000  84.380000 1.475000 ;
      RECT  83.600000  1.475000  84.030000 1.635000 ;
      RECT  83.600000  1.635000  83.930000 2.465000 ;
      RECT  83.860000  1.305000  84.380000 1.465000 ;
      RECT  83.965000  0.755000  84.135000 1.205000 ;
      RECT  83.965000  1.205000  84.380000 1.305000 ;
      RECT  84.200000  1.645000  84.370000 2.295000 ;
      RECT  84.200000  2.295000  85.365000 2.465000 ;
      RECT  84.305000  0.255000  85.450000 0.425000 ;
      RECT  84.305000  0.425000  84.475000 0.770000 ;
      RECT  84.585000  1.755000  85.015000 2.125000 ;
      RECT  84.645000  0.595000  84.975000 0.885000 ;
      RECT  84.725000  0.885000  84.895000 1.755000 ;
      RECT  85.145000  0.425000  85.450000 0.715000 ;
      RECT  85.145000  0.715000  86.335000 0.885000 ;
      RECT  85.145000  0.885000  85.450000 0.925000 ;
      RECT  85.195000  1.495000  86.385000 1.665000 ;
      RECT  85.195000  1.665000  85.365000 2.295000 ;
      RECT  85.565000  1.055000  86.385000 1.325000 ;
      RECT  85.585000  1.835000  85.915000 2.105000 ;
      RECT  85.585000  2.105000  85.885000 2.635000 ;
      RECT  85.620000  0.085000  85.835000 0.545000 ;
      RECT  86.005000  0.255000  86.335000 0.715000 ;
      RECT  86.055000  2.210000  86.385000 2.465000 ;
      RECT  86.085000  1.665000  86.385000 2.210000 ;
      RECT  86.575000  1.055000  87.395000 1.325000 ;
      RECT  86.575000  1.495000  87.765000 1.665000 ;
      RECT  86.575000  1.665000  86.875000 2.210000 ;
      RECT  86.575000  2.210000  86.905000 2.465000 ;
      RECT  86.625000  0.255000  86.955000 0.715000 ;
      RECT  86.625000  0.715000  87.815000 0.885000 ;
      RECT  87.045000  1.835000  87.375000 2.105000 ;
      RECT  87.075000  2.105000  87.375000 2.635000 ;
      RECT  87.125000  0.085000  87.340000 0.545000 ;
      RECT  87.510000  0.255000  88.655000 0.425000 ;
      RECT  87.510000  0.425000  87.815000 0.715000 ;
      RECT  87.510000  0.885000  87.815000 0.925000 ;
      RECT  87.595000  1.665000  87.765000 2.295000 ;
      RECT  87.595000  2.295000  88.760000 2.465000 ;
      RECT  87.945000  1.755000  88.375000 2.125000 ;
      RECT  87.985000  0.595000  88.315000 0.885000 ;
      RECT  88.065000  0.885000  88.235000 1.755000 ;
      RECT  88.485000  0.425000  88.655000 0.770000 ;
      RECT  88.580000  1.205000  88.995000 1.305000 ;
      RECT  88.580000  1.305000  89.100000 1.465000 ;
      RECT  88.580000  1.465000  89.360000 1.475000 ;
      RECT  88.590000  1.645000  88.760000 2.295000 ;
      RECT  88.825000  0.585000  89.405000 0.755000 ;
      RECT  88.825000  0.755000  88.995000 1.205000 ;
      RECT  88.930000  1.475000  89.360000 1.635000 ;
      RECT  89.030000  1.635000  89.360000 2.465000 ;
      RECT  89.155000  0.330000  89.405000 0.585000 ;
      RECT  89.270000  1.025000  89.605000 1.295000 ;
      RECT  89.535000  1.465000  89.865000 2.635000 ;
      RECT  89.575000  0.085000  89.825000 0.660000 ;
      RECT  89.795000  1.025000  90.130000 1.295000 ;
      RECT  89.995000  0.330000  90.245000 0.585000 ;
      RECT  89.995000  0.585000  90.575000 0.755000 ;
      RECT  90.040000  1.465000  90.820000 1.475000 ;
      RECT  90.040000  1.475000  90.470000 1.635000 ;
      RECT  90.040000  1.635000  90.370000 2.465000 ;
      RECT  90.300000  1.305000  90.820000 1.465000 ;
      RECT  90.405000  0.755000  90.575000 1.205000 ;
      RECT  90.405000  1.205000  90.820000 1.305000 ;
      RECT  90.640000  1.645000  90.810000 2.295000 ;
      RECT  90.640000  2.295000  91.805000 2.465000 ;
      RECT  90.745000  0.255000  91.890000 0.425000 ;
      RECT  90.745000  0.425000  90.915000 0.770000 ;
      RECT  91.025000  1.755000  91.455000 2.125000 ;
      RECT  91.085000  0.595000  91.415000 0.885000 ;
      RECT  91.165000  0.885000  91.335000 1.755000 ;
      RECT  91.585000  0.425000  91.890000 0.715000 ;
      RECT  91.585000  0.715000  92.775000 0.885000 ;
      RECT  91.585000  0.885000  91.890000 0.925000 ;
      RECT  91.635000  1.495000  92.825000 1.665000 ;
      RECT  91.635000  1.665000  91.805000 2.295000 ;
      RECT  92.005000  1.055000  92.825000 1.325000 ;
      RECT  92.025000  1.835000  92.355000 2.105000 ;
      RECT  92.025000  2.105000  92.325000 2.635000 ;
      RECT  92.060000  0.085000  92.275000 0.545000 ;
      RECT  92.445000  0.255000  92.775000 0.715000 ;
      RECT  92.495000  2.210000  92.825000 2.465000 ;
      RECT  92.525000  1.665000  92.825000 2.210000 ;
      RECT  93.015000  1.055000  93.835000 1.325000 ;
      RECT  93.015000  1.495000  94.205000 1.665000 ;
      RECT  93.015000  1.665000  93.315000 2.210000 ;
      RECT  93.015000  2.210000  93.345000 2.465000 ;
      RECT  93.065000  0.255000  93.395000 0.715000 ;
      RECT  93.065000  0.715000  94.255000 0.885000 ;
      RECT  93.485000  1.835000  93.815000 2.105000 ;
      RECT  93.515000  2.105000  93.815000 2.635000 ;
      RECT  93.565000  0.085000  93.780000 0.545000 ;
      RECT  93.950000  0.255000  95.095000 0.425000 ;
      RECT  93.950000  0.425000  94.255000 0.715000 ;
      RECT  93.950000  0.885000  94.255000 0.925000 ;
      RECT  94.035000  1.665000  94.205000 2.295000 ;
      RECT  94.035000  2.295000  95.200000 2.465000 ;
      RECT  94.385000  1.755000  94.815000 2.125000 ;
      RECT  94.425000  0.595000  94.755000 0.885000 ;
      RECT  94.505000  0.885000  94.675000 1.755000 ;
      RECT  94.925000  0.425000  95.095000 0.770000 ;
      RECT  95.020000  1.205000  95.435000 1.305000 ;
      RECT  95.020000  1.305000  95.540000 1.465000 ;
      RECT  95.020000  1.465000  95.800000 1.475000 ;
      RECT  95.030000  1.645000  95.200000 2.295000 ;
      RECT  95.265000  0.585000  95.845000 0.755000 ;
      RECT  95.265000  0.755000  95.435000 1.205000 ;
      RECT  95.370000  1.475000  95.800000 1.635000 ;
      RECT  95.470000  1.635000  95.800000 2.465000 ;
      RECT  95.595000  0.330000  95.845000 0.585000 ;
      RECT  95.710000  1.025000  96.045000 1.295000 ;
      RECT  95.975000  1.465000  96.305000 2.635000 ;
      RECT  96.015000  0.085000  96.265000 0.660000 ;
      RECT  96.235000  1.025000  96.570000 1.295000 ;
      RECT  96.435000  0.330000  96.685000 0.585000 ;
      RECT  96.435000  0.585000  97.015000 0.755000 ;
      RECT  96.480000  1.465000  97.260000 1.475000 ;
      RECT  96.480000  1.475000  96.910000 1.635000 ;
      RECT  96.480000  1.635000  96.810000 2.465000 ;
      RECT  96.740000  1.305000  97.260000 1.465000 ;
      RECT  96.845000  0.755000  97.015000 1.205000 ;
      RECT  96.845000  1.205000  97.260000 1.305000 ;
      RECT  97.080000  1.645000  97.250000 2.295000 ;
      RECT  97.080000  2.295000  98.245000 2.465000 ;
      RECT  97.185000  0.255000  98.330000 0.425000 ;
      RECT  97.185000  0.425000  97.355000 0.770000 ;
      RECT  97.465000  1.755000  97.895000 2.125000 ;
      RECT  97.525000  0.595000  97.855000 0.885000 ;
      RECT  97.605000  0.885000  97.775000 1.755000 ;
      RECT  98.025000  0.425000  98.330000 0.715000 ;
      RECT  98.025000  0.715000  99.215000 0.885000 ;
      RECT  98.025000  0.885000  98.330000 0.925000 ;
      RECT  98.075000  1.495000  99.265000 1.665000 ;
      RECT  98.075000  1.665000  98.245000 2.295000 ;
      RECT  98.445000  1.055000  99.265000 1.325000 ;
      RECT  98.465000  1.835000  98.795000 2.105000 ;
      RECT  98.465000  2.105000  98.765000 2.635000 ;
      RECT  98.500000  0.085000  98.715000 0.545000 ;
      RECT  98.885000  0.255000  99.215000 0.715000 ;
      RECT  98.935000  2.210000  99.265000 2.465000 ;
      RECT  98.965000  1.665000  99.265000 2.210000 ;
      RECT  99.455000  1.055000 100.275000 1.325000 ;
      RECT  99.455000  1.495000 100.645000 1.665000 ;
      RECT  99.455000  1.665000  99.755000 2.210000 ;
      RECT  99.455000  2.210000  99.785000 2.465000 ;
      RECT  99.505000  0.255000  99.835000 0.715000 ;
      RECT  99.505000  0.715000 100.695000 0.885000 ;
      RECT  99.925000  1.835000 100.255000 2.105000 ;
      RECT  99.955000  2.105000 100.255000 2.635000 ;
      RECT 100.005000  0.085000 100.220000 0.545000 ;
      RECT 100.390000  0.255000 101.535000 0.425000 ;
      RECT 100.390000  0.425000 100.695000 0.715000 ;
      RECT 100.390000  0.885000 100.695000 0.925000 ;
      RECT 100.475000  1.665000 100.645000 2.295000 ;
      RECT 100.475000  2.295000 101.640000 2.465000 ;
      RECT 100.825000  1.755000 101.255000 2.125000 ;
      RECT 100.865000  0.595000 101.195000 0.885000 ;
      RECT 100.945000  0.885000 101.115000 1.755000 ;
      RECT 101.365000  0.425000 101.535000 0.770000 ;
      RECT 101.460000  1.205000 101.875000 1.305000 ;
      RECT 101.460000  1.305000 101.980000 1.465000 ;
      RECT 101.460000  1.465000 102.240000 1.475000 ;
      RECT 101.470000  1.645000 101.640000 2.295000 ;
      RECT 101.705000  0.585000 102.285000 0.755000 ;
      RECT 101.705000  0.755000 101.875000 1.205000 ;
      RECT 101.810000  1.475000 102.240000 1.635000 ;
      RECT 101.910000  1.635000 102.240000 2.465000 ;
      RECT 102.035000  0.330000 102.285000 0.585000 ;
      RECT 102.150000  1.025000 102.485000 1.295000 ;
      RECT 102.415000  1.465000 102.745000 2.635000 ;
      RECT 102.455000  0.085000 102.705000 0.660000 ;
      RECT 102.675000  1.025000 103.010000 1.295000 ;
      RECT 102.875000  0.330000 103.125000 0.585000 ;
      RECT 102.875000  0.585000 103.455000 0.755000 ;
      RECT 102.920000  1.465000 103.700000 1.475000 ;
      RECT 102.920000  1.475000 103.350000 1.635000 ;
      RECT 102.920000  1.635000 103.250000 2.465000 ;
      RECT 103.180000  1.305000 103.700000 1.465000 ;
      RECT 103.285000  0.755000 103.455000 1.205000 ;
      RECT 103.285000  1.205000 103.700000 1.305000 ;
      RECT 103.520000  1.645000 103.690000 2.295000 ;
      RECT 103.520000  2.295000 104.685000 2.465000 ;
      RECT 103.625000  0.255000 104.770000 0.425000 ;
      RECT 103.625000  0.425000 103.795000 0.770000 ;
      RECT 103.905000  1.755000 104.335000 2.125000 ;
      RECT 103.965000  0.595000 104.295000 0.885000 ;
      RECT 104.045000  0.885000 104.215000 1.755000 ;
      RECT 104.465000  0.425000 104.770000 0.715000 ;
      RECT 104.465000  0.715000 105.655000 0.885000 ;
      RECT 104.465000  0.885000 104.770000 0.925000 ;
      RECT 104.515000  1.495000 105.705000 1.665000 ;
      RECT 104.515000  1.665000 104.685000 2.295000 ;
      RECT 104.885000  1.055000 105.705000 1.325000 ;
      RECT 104.905000  1.835000 105.235000 2.105000 ;
      RECT 104.905000  2.105000 105.205000 2.635000 ;
      RECT 104.940000  0.085000 105.155000 0.545000 ;
      RECT 105.325000  0.255000 105.655000 0.715000 ;
      RECT 105.375000  2.210000 105.705000 2.465000 ;
      RECT 105.405000  1.665000 105.705000 2.210000 ;
      RECT 105.800000  5.355000 225.400000 5.525000 ;
      RECT 105.885000  0.995000 106.480000 1.325000 ;
      RECT 105.885000  4.115000 106.480000 4.445000 ;
      RECT 106.020000  1.605000 106.320000 2.635000 ;
      RECT 106.020000  2.805000 106.320000 3.835000 ;
      RECT 106.070000  0.085000 106.360000 0.610000 ;
      RECT 106.070000  4.830000 106.360000 5.355000 ;
      RECT 106.490000  1.605000 106.820000 2.465000 ;
      RECT 106.490000  2.975000 106.820000 3.835000 ;
      RECT 106.570000  0.280000 106.820000 0.825000 ;
      RECT 106.570000  4.615000 106.820000 5.160000 ;
      RECT 106.650000  0.825000 106.820000 1.065000 ;
      RECT 106.650000  1.065000 107.835000 1.395000 ;
      RECT 106.650000  1.395000 106.820000 1.605000 ;
      RECT 106.650000  3.835000 106.820000 4.045000 ;
      RECT 106.650000  4.045000 107.835000 4.375000 ;
      RECT 106.650000  4.375000 106.820000 4.615000 ;
      RECT 106.990000  0.085000 107.280000 0.610000 ;
      RECT 106.990000  4.830000 107.280000 5.355000 ;
      RECT 107.015000  1.605000 107.290000 2.635000 ;
      RECT 107.015000  2.805000 107.290000 3.835000 ;
      RECT 107.535000  1.565000 107.835000 2.465000 ;
      RECT 107.535000  2.975000 107.835000 3.875000 ;
      RECT 107.785000  0.255000 109.815000 0.425000 ;
      RECT 107.785000  0.425000 108.035000 0.770000 ;
      RECT 107.785000  4.670000 108.035000 5.015000 ;
      RECT 107.785000  5.015000 109.815000 5.185000 ;
      RECT 108.005000  1.065000 109.275000 1.365000 ;
      RECT 108.005000  1.365000 108.335000 4.075000 ;
      RECT 108.005000  4.075000 109.275000 4.375000 ;
      RECT 108.205000  0.595000 108.535000 1.065000 ;
      RECT 108.205000  4.375000 108.535000 4.845000 ;
      RECT 108.505000  1.535000 108.775000 2.465000 ;
      RECT 108.505000  2.975000 108.775000 3.905000 ;
      RECT 108.705000  0.425000 108.875000 0.770000 ;
      RECT 108.705000  4.670000 108.875000 5.015000 ;
      RECT 108.945000  1.365000 109.275000 4.075000 ;
      RECT 109.045000  0.595000 109.375000 0.885000 ;
      RECT 109.045000  0.885000 109.275000 1.065000 ;
      RECT 109.045000  4.375000 109.275000 4.555000 ;
      RECT 109.045000  4.555000 109.375000 4.845000 ;
      RECT 109.445000  1.495000 111.675000 1.665000 ;
      RECT 109.445000  1.665000 109.745000 2.465000 ;
      RECT 109.445000  2.635000 114.575000 2.805000 ;
      RECT 109.445000  2.975000 109.745000 3.775000 ;
      RECT 109.445000  3.775000 111.675000 3.945000 ;
      RECT 109.545000  0.425000 109.815000 0.715000 ;
      RECT 109.545000  0.715000 111.675000 0.885000 ;
      RECT 109.545000  4.555000 111.675000 4.725000 ;
      RECT 109.545000  4.725000 109.815000 5.015000 ;
      RECT 109.965000  1.835000 110.235000 2.635000 ;
      RECT 109.965000  2.805000 110.235000 3.605000 ;
      RECT 109.985000  0.085000 110.235000 0.545000 ;
      RECT 109.985000  4.895000 110.235000 5.355000 ;
      RECT 110.405000  0.255000 110.735000 0.715000 ;
      RECT 110.405000  1.665000 110.735000 2.465000 ;
      RECT 110.405000  2.975000 110.735000 3.775000 ;
      RECT 110.405000  4.725000 110.735000 5.185000 ;
      RECT 110.455000  1.055000 111.845000 1.325000 ;
      RECT 110.455000  4.115000 111.845000 4.385000 ;
      RECT 110.905000  0.085000 111.175000 0.545000 ;
      RECT 110.905000  1.835000 111.175000 2.635000 ;
      RECT 110.905000  2.805000 111.175000 3.605000 ;
      RECT 110.905000  4.895000 111.175000 5.355000 ;
      RECT 111.345000  0.255000 111.675000 0.715000 ;
      RECT 111.345000  1.665000 111.675000 2.465000 ;
      RECT 111.345000  2.975000 111.675000 3.775000 ;
      RECT 111.345000  4.725000 111.675000 5.185000 ;
      RECT 111.845000  0.085000 112.175000 0.885000 ;
      RECT 111.845000  1.495000 112.175000 2.635000 ;
      RECT 111.845000  2.805000 112.175000 3.945000 ;
      RECT 111.845000  4.555000 112.175000 5.355000 ;
      RECT 112.175000  1.055000 113.565000 1.325000 ;
      RECT 112.175000  4.115000 113.565000 4.385000 ;
      RECT 112.345000  0.255000 112.675000 0.715000 ;
      RECT 112.345000  0.715000 114.475000 0.885000 ;
      RECT 112.345000  1.495000 114.575000 1.665000 ;
      RECT 112.345000  1.665000 112.675000 2.465000 ;
      RECT 112.345000  2.975000 112.675000 3.775000 ;
      RECT 112.345000  3.775000 114.575000 3.945000 ;
      RECT 112.345000  4.555000 114.475000 4.725000 ;
      RECT 112.345000  4.725000 112.675000 5.185000 ;
      RECT 112.845000  0.085000 113.115000 0.545000 ;
      RECT 112.845000  1.835000 113.115000 2.635000 ;
      RECT 112.845000  2.805000 113.115000 3.605000 ;
      RECT 112.845000  4.895000 113.115000 5.355000 ;
      RECT 113.285000  0.255000 113.615000 0.715000 ;
      RECT 113.285000  1.665000 113.615000 2.465000 ;
      RECT 113.285000  2.975000 113.615000 3.775000 ;
      RECT 113.285000  4.725000 113.615000 5.185000 ;
      RECT 113.785000  0.085000 114.035000 0.545000 ;
      RECT 113.785000  1.835000 114.055000 2.635000 ;
      RECT 113.785000  2.805000 114.055000 3.605000 ;
      RECT 113.785000  4.895000 114.035000 5.355000 ;
      RECT 114.205000  0.255000 116.235000 0.425000 ;
      RECT 114.205000  0.425000 114.475000 0.715000 ;
      RECT 114.205000  4.725000 114.475000 5.015000 ;
      RECT 114.205000  5.015000 116.235000 5.185000 ;
      RECT 114.275000  1.665000 114.575000 2.465000 ;
      RECT 114.275000  2.975000 114.575000 3.775000 ;
      RECT 114.645000  0.595000 114.975000 0.885000 ;
      RECT 114.645000  4.555000 114.975000 4.845000 ;
      RECT 114.745000  0.885000 114.975000 1.065000 ;
      RECT 114.745000  1.065000 116.015000 1.365000 ;
      RECT 114.745000  1.365000 115.075000 4.075000 ;
      RECT 114.745000  4.075000 116.015000 4.375000 ;
      RECT 114.745000  4.375000 114.975000 4.555000 ;
      RECT 115.145000  0.425000 115.315000 0.770000 ;
      RECT 115.145000  4.670000 115.315000 5.015000 ;
      RECT 115.245000  1.535000 115.515000 2.465000 ;
      RECT 115.245000  2.975000 115.515000 3.905000 ;
      RECT 115.485000  0.595000 115.815000 1.065000 ;
      RECT 115.485000  4.375000 115.815000 4.845000 ;
      RECT 115.685000  1.365000 116.015000 4.075000 ;
      RECT 115.985000  0.425000 116.235000 0.770000 ;
      RECT 115.985000  4.670000 116.235000 5.015000 ;
      RECT 116.185000  1.065000 117.370000 1.395000 ;
      RECT 116.185000  1.565000 116.485000 2.465000 ;
      RECT 116.185000  2.635000 120.255000 2.805000 ;
      RECT 116.185000  2.975000 116.485000 3.875000 ;
      RECT 116.185000  4.045000 117.370000 4.375000 ;
      RECT 116.730000  1.605000 117.005000 2.635000 ;
      RECT 116.730000  2.805000 117.005000 3.835000 ;
      RECT 116.740000  0.085000 117.030000 0.610000 ;
      RECT 116.740000  4.830000 117.030000 5.355000 ;
      RECT 117.200000  0.280000 117.450000 0.825000 ;
      RECT 117.200000  0.825000 117.370000 1.065000 ;
      RECT 117.200000  1.395000 117.370000 1.605000 ;
      RECT 117.200000  1.605000 117.530000 2.465000 ;
      RECT 117.200000  2.975000 117.530000 3.835000 ;
      RECT 117.200000  3.835000 117.370000 4.045000 ;
      RECT 117.200000  4.375000 117.370000 4.615000 ;
      RECT 117.200000  4.615000 117.450000 5.160000 ;
      RECT 117.540000  0.995000 118.135000 1.325000 ;
      RECT 117.540000  4.115000 118.135000 4.445000 ;
      RECT 117.660000  0.085000 117.950000 0.610000 ;
      RECT 117.660000  4.830000 117.950000 5.355000 ;
      RECT 117.700000  1.605000 118.000000 2.635000 ;
      RECT 117.700000  2.805000 118.000000 3.835000 ;
      RECT 118.305000  0.995000 118.900000 1.325000 ;
      RECT 118.305000  4.115000 118.900000 4.445000 ;
      RECT 118.440000  1.605000 118.740000 2.635000 ;
      RECT 118.440000  2.805000 118.740000 3.835000 ;
      RECT 118.490000  0.085000 118.780000 0.610000 ;
      RECT 118.490000  4.830000 118.780000 5.355000 ;
      RECT 118.910000  1.605000 119.240000 2.465000 ;
      RECT 118.910000  2.975000 119.240000 3.835000 ;
      RECT 118.990000  0.280000 119.240000 0.825000 ;
      RECT 118.990000  4.615000 119.240000 5.160000 ;
      RECT 119.070000  0.825000 119.240000 1.065000 ;
      RECT 119.070000  1.065000 120.255000 1.395000 ;
      RECT 119.070000  1.395000 119.240000 1.605000 ;
      RECT 119.070000  3.835000 119.240000 4.045000 ;
      RECT 119.070000  4.045000 120.255000 4.375000 ;
      RECT 119.070000  4.375000 119.240000 4.615000 ;
      RECT 119.410000  0.085000 119.700000 0.610000 ;
      RECT 119.410000  4.830000 119.700000 5.355000 ;
      RECT 119.435000  1.605000 119.710000 2.635000 ;
      RECT 119.435000  2.805000 119.710000 3.835000 ;
      RECT 119.955000  1.565000 120.255000 2.465000 ;
      RECT 119.955000  2.975000 120.255000 3.875000 ;
      RECT 120.205000  0.255000 122.235000 0.425000 ;
      RECT 120.205000  0.425000 120.455000 0.770000 ;
      RECT 120.205000  4.670000 120.455000 5.015000 ;
      RECT 120.205000  5.015000 122.235000 5.185000 ;
      RECT 120.425000  1.065000 121.695000 1.365000 ;
      RECT 120.425000  1.365000 120.755000 4.075000 ;
      RECT 120.425000  4.075000 121.695000 4.375000 ;
      RECT 120.625000  0.595000 120.955000 1.065000 ;
      RECT 120.625000  4.375000 120.955000 4.845000 ;
      RECT 120.925000  1.535000 121.195000 2.465000 ;
      RECT 120.925000  2.975000 121.195000 3.905000 ;
      RECT 121.125000  0.425000 121.295000 0.770000 ;
      RECT 121.125000  4.670000 121.295000 5.015000 ;
      RECT 121.365000  1.365000 121.695000 4.075000 ;
      RECT 121.465000  0.595000 121.795000 0.885000 ;
      RECT 121.465000  0.885000 121.695000 1.065000 ;
      RECT 121.465000  4.375000 121.695000 4.555000 ;
      RECT 121.465000  4.555000 121.795000 4.845000 ;
      RECT 121.865000  1.495000 124.095000 1.665000 ;
      RECT 121.865000  1.665000 122.165000 2.465000 ;
      RECT 121.865000  2.635000 126.995000 2.805000 ;
      RECT 121.865000  2.975000 122.165000 3.775000 ;
      RECT 121.865000  3.775000 124.095000 3.945000 ;
      RECT 121.965000  0.425000 122.235000 0.715000 ;
      RECT 121.965000  0.715000 124.095000 0.885000 ;
      RECT 121.965000  4.555000 124.095000 4.725000 ;
      RECT 121.965000  4.725000 122.235000 5.015000 ;
      RECT 122.385000  1.835000 122.655000 2.635000 ;
      RECT 122.385000  2.805000 122.655000 3.605000 ;
      RECT 122.405000  0.085000 122.655000 0.545000 ;
      RECT 122.405000  4.895000 122.655000 5.355000 ;
      RECT 122.825000  0.255000 123.155000 0.715000 ;
      RECT 122.825000  1.665000 123.155000 2.465000 ;
      RECT 122.825000  2.975000 123.155000 3.775000 ;
      RECT 122.825000  4.725000 123.155000 5.185000 ;
      RECT 122.875000  1.055000 124.265000 1.325000 ;
      RECT 122.875000  4.115000 124.265000 4.385000 ;
      RECT 123.325000  0.085000 123.595000 0.545000 ;
      RECT 123.325000  1.835000 123.595000 2.635000 ;
      RECT 123.325000  2.805000 123.595000 3.605000 ;
      RECT 123.325000  4.895000 123.595000 5.355000 ;
      RECT 123.765000  0.255000 124.095000 0.715000 ;
      RECT 123.765000  1.665000 124.095000 2.465000 ;
      RECT 123.765000  2.975000 124.095000 3.775000 ;
      RECT 123.765000  4.725000 124.095000 5.185000 ;
      RECT 124.265000  0.085000 124.595000 0.885000 ;
      RECT 124.265000  1.495000 124.595000 2.635000 ;
      RECT 124.265000  2.805000 124.595000 3.945000 ;
      RECT 124.265000  4.555000 124.595000 5.355000 ;
      RECT 124.595000  1.055000 125.985000 1.325000 ;
      RECT 124.595000  4.115000 125.985000 4.385000 ;
      RECT 124.765000  0.255000 125.095000 0.715000 ;
      RECT 124.765000  0.715000 126.895000 0.885000 ;
      RECT 124.765000  1.495000 126.995000 1.665000 ;
      RECT 124.765000  1.665000 125.095000 2.465000 ;
      RECT 124.765000  2.975000 125.095000 3.775000 ;
      RECT 124.765000  3.775000 126.995000 3.945000 ;
      RECT 124.765000  4.555000 126.895000 4.725000 ;
      RECT 124.765000  4.725000 125.095000 5.185000 ;
      RECT 125.265000  0.085000 125.535000 0.545000 ;
      RECT 125.265000  1.835000 125.535000 2.635000 ;
      RECT 125.265000  2.805000 125.535000 3.605000 ;
      RECT 125.265000  4.895000 125.535000 5.355000 ;
      RECT 125.705000  0.255000 126.035000 0.715000 ;
      RECT 125.705000  1.665000 126.035000 2.465000 ;
      RECT 125.705000  2.975000 126.035000 3.775000 ;
      RECT 125.705000  4.725000 126.035000 5.185000 ;
      RECT 126.205000  0.085000 126.455000 0.545000 ;
      RECT 126.205000  1.835000 126.475000 2.635000 ;
      RECT 126.205000  2.805000 126.475000 3.605000 ;
      RECT 126.205000  4.895000 126.455000 5.355000 ;
      RECT 126.625000  0.255000 128.655000 0.425000 ;
      RECT 126.625000  0.425000 126.895000 0.715000 ;
      RECT 126.625000  4.725000 126.895000 5.015000 ;
      RECT 126.625000  5.015000 128.655000 5.185000 ;
      RECT 126.695000  1.665000 126.995000 2.465000 ;
      RECT 126.695000  2.975000 126.995000 3.775000 ;
      RECT 127.065000  0.595000 127.395000 0.885000 ;
      RECT 127.065000  4.555000 127.395000 4.845000 ;
      RECT 127.165000  0.885000 127.395000 1.065000 ;
      RECT 127.165000  1.065000 128.435000 1.365000 ;
      RECT 127.165000  1.365000 127.495000 4.075000 ;
      RECT 127.165000  4.075000 128.435000 4.375000 ;
      RECT 127.165000  4.375000 127.395000 4.555000 ;
      RECT 127.565000  0.425000 127.735000 0.770000 ;
      RECT 127.565000  4.670000 127.735000 5.015000 ;
      RECT 127.665000  1.535000 127.935000 2.465000 ;
      RECT 127.665000  2.975000 127.935000 3.905000 ;
      RECT 127.905000  0.595000 128.235000 1.065000 ;
      RECT 127.905000  4.375000 128.235000 4.845000 ;
      RECT 128.105000  1.365000 128.435000 4.075000 ;
      RECT 128.405000  0.425000 128.655000 0.770000 ;
      RECT 128.405000  4.670000 128.655000 5.015000 ;
      RECT 128.605000  1.065000 129.790000 1.395000 ;
      RECT 128.605000  1.565000 128.905000 2.465000 ;
      RECT 128.605000  2.635000 131.560000 2.805000 ;
      RECT 128.605000  2.975000 128.905000 3.875000 ;
      RECT 128.605000  4.045000 129.790000 4.375000 ;
      RECT 129.150000  1.605000 129.425000 2.635000 ;
      RECT 129.150000  2.805000 129.425000 3.835000 ;
      RECT 129.160000  0.085000 129.450000 0.610000 ;
      RECT 129.160000  4.830000 129.450000 5.355000 ;
      RECT 129.620000  0.280000 129.870000 0.825000 ;
      RECT 129.620000  0.825000 129.790000 1.065000 ;
      RECT 129.620000  1.395000 129.790000 1.605000 ;
      RECT 129.620000  1.605000 129.950000 2.465000 ;
      RECT 129.620000  2.975000 129.950000 3.835000 ;
      RECT 129.620000  3.835000 129.790000 4.045000 ;
      RECT 129.620000  4.375000 129.790000 4.615000 ;
      RECT 129.620000  4.615000 129.870000 5.160000 ;
      RECT 129.960000  0.995000 130.555000 1.325000 ;
      RECT 129.960000  4.115000 130.555000 4.445000 ;
      RECT 130.080000  0.085000 130.370000 0.610000 ;
      RECT 130.080000  4.830000 130.370000 5.355000 ;
      RECT 130.120000  1.605000 130.420000 2.635000 ;
      RECT 130.120000  2.805000 130.420000 3.835000 ;
      RECT 130.735000  1.495000 131.065000 2.635000 ;
      RECT 130.735000  2.805000 131.065000 3.945000 ;
      RECT 130.770000  0.085000 131.030000 0.885000 ;
      RECT 130.770000  4.555000 131.030000 5.355000 ;
      RECT 130.975000  1.055000 131.370000 1.325000 ;
      RECT 130.975000  4.115000 131.370000 4.385000 ;
      RECT 131.200000  0.395000 131.475000 0.625000 ;
      RECT 131.200000  0.625000 131.370000 1.055000 ;
      RECT 131.200000  4.385000 131.370000 4.815000 ;
      RECT 131.200000  4.815000 131.475000 5.045000 ;
      RECT 131.540000  0.835000 131.930000 1.005000 ;
      RECT 131.540000  1.005000 131.710000 1.755000 ;
      RECT 131.540000  1.755000 131.935000 1.805000 ;
      RECT 131.540000  1.805000 132.060000 1.985000 ;
      RECT 131.540000  3.455000 132.060000 3.635000 ;
      RECT 131.540000  3.635000 131.935000 3.685000 ;
      RECT 131.540000  3.685000 131.710000 4.435000 ;
      RECT 131.540000  4.435000 131.930000 4.605000 ;
      RECT 131.685000  0.330000 131.930000 0.835000 ;
      RECT 131.685000  4.605000 131.930000 5.110000 ;
      RECT 131.730000  1.985000 132.060000 2.465000 ;
      RECT 131.730000  2.465000 131.935000 2.975000 ;
      RECT 131.730000  2.975000 132.060000 3.455000 ;
      RECT 131.880000  1.175000 132.270000 1.465000 ;
      RECT 131.880000  1.465000 132.580000 1.505000 ;
      RECT 131.880000  3.935000 132.580000 3.975000 ;
      RECT 131.880000  3.975000 132.270000 4.265000 ;
      RECT 132.100000  0.585000 132.540000 0.755000 ;
      RECT 132.100000  0.755000 132.270000 1.175000 ;
      RECT 132.100000  1.505000 132.580000 1.635000 ;
      RECT 132.100000  3.805000 132.580000 3.935000 ;
      RECT 132.100000  4.265000 132.270000 4.685000 ;
      RECT 132.100000  4.685000 132.540000 4.855000 ;
      RECT 132.105000  2.635000 133.775000 2.805000 ;
      RECT 132.250000  1.635000 132.580000 2.465000 ;
      RECT 132.250000  2.975000 132.580000 3.805000 ;
      RECT 132.290000  0.330000 132.540000 0.585000 ;
      RECT 132.290000  4.855000 132.540000 5.110000 ;
      RECT 132.445000  0.945000 132.845000 1.295000 ;
      RECT 132.445000  4.145000 132.845000 4.495000 ;
      RECT 132.775000  0.085000 133.105000 0.660000 ;
      RECT 132.775000  1.465000 133.105000 2.635000 ;
      RECT 132.775000  2.805000 133.105000 3.975000 ;
      RECT 132.775000  4.780000 133.105000 5.355000 ;
      RECT 133.035000  0.945000 133.435000 1.295000 ;
      RECT 133.035000  4.145000 133.435000 4.495000 ;
      RECT 133.300000  1.465000 134.000000 1.505000 ;
      RECT 133.300000  1.505000 133.780000 1.635000 ;
      RECT 133.300000  1.635000 133.630000 2.465000 ;
      RECT 133.300000  2.975000 133.630000 3.805000 ;
      RECT 133.300000  3.805000 133.780000 3.935000 ;
      RECT 133.300000  3.935000 134.000000 3.975000 ;
      RECT 133.340000  0.330000 133.590000 0.585000 ;
      RECT 133.340000  0.585000 133.780000 0.755000 ;
      RECT 133.340000  4.685000 133.780000 4.855000 ;
      RECT 133.340000  4.855000 133.590000 5.110000 ;
      RECT 133.610000  0.755000 133.780000 1.175000 ;
      RECT 133.610000  1.175000 134.000000 1.465000 ;
      RECT 133.610000  3.975000 134.000000 4.265000 ;
      RECT 133.610000  4.265000 133.780000 4.685000 ;
      RECT 133.820000  1.805000 134.340000 1.985000 ;
      RECT 133.820000  1.985000 134.150000 2.465000 ;
      RECT 133.820000  2.975000 134.150000 3.455000 ;
      RECT 133.820000  3.455000 134.340000 3.635000 ;
      RECT 133.945000  1.755000 134.340000 1.805000 ;
      RECT 133.945000  2.465000 134.150000 2.975000 ;
      RECT 133.945000  3.635000 134.340000 3.685000 ;
      RECT 133.950000  0.330000 134.195000 0.835000 ;
      RECT 133.950000  0.835000 134.340000 1.005000 ;
      RECT 133.950000  4.435000 134.340000 4.605000 ;
      RECT 133.950000  4.605000 134.195000 5.110000 ;
      RECT 134.170000  1.005000 134.340000 1.755000 ;
      RECT 134.170000  3.685000 134.340000 4.435000 ;
      RECT 134.320000  2.635000 135.700000 2.805000 ;
      RECT 134.405000  0.395000 134.680000 0.625000 ;
      RECT 134.405000  4.815000 134.680000 5.045000 ;
      RECT 134.510000  0.625000 134.680000 1.055000 ;
      RECT 134.510000  1.055000 134.905000 1.325000 ;
      RECT 134.510000  4.115000 134.905000 4.385000 ;
      RECT 134.510000  4.385000 134.680000 4.815000 ;
      RECT 134.815000  1.495000 135.205000 2.635000 ;
      RECT 134.815000  2.805000 135.205000 3.945000 ;
      RECT 134.850000  0.085000 135.170000 0.885000 ;
      RECT 134.850000  4.555000 135.170000 5.355000 ;
      RECT 135.115000  1.055000 135.510000 1.325000 ;
      RECT 135.115000  4.115000 135.510000 4.385000 ;
      RECT 135.340000  0.395000 135.615000 0.625000 ;
      RECT 135.340000  0.625000 135.510000 1.055000 ;
      RECT 135.340000  4.385000 135.510000 4.815000 ;
      RECT 135.340000  4.815000 135.615000 5.045000 ;
      RECT 135.680000  0.835000 136.070000 1.005000 ;
      RECT 135.680000  1.005000 135.850000 1.755000 ;
      RECT 135.680000  1.755000 136.075000 1.805000 ;
      RECT 135.680000  1.805000 136.200000 1.985000 ;
      RECT 135.680000  3.455000 136.200000 3.635000 ;
      RECT 135.680000  3.635000 136.075000 3.685000 ;
      RECT 135.680000  3.685000 135.850000 4.435000 ;
      RECT 135.680000  4.435000 136.070000 4.605000 ;
      RECT 135.825000  0.330000 136.070000 0.835000 ;
      RECT 135.825000  4.605000 136.070000 5.110000 ;
      RECT 135.870000  1.985000 136.200000 2.465000 ;
      RECT 135.870000  2.465000 136.075000 2.975000 ;
      RECT 135.870000  2.975000 136.200000 3.455000 ;
      RECT 136.020000  1.175000 136.410000 1.465000 ;
      RECT 136.020000  1.465000 136.720000 1.505000 ;
      RECT 136.020000  3.935000 136.720000 3.975000 ;
      RECT 136.020000  3.975000 136.410000 4.265000 ;
      RECT 136.240000  0.585000 136.680000 0.755000 ;
      RECT 136.240000  0.755000 136.410000 1.175000 ;
      RECT 136.240000  1.505000 136.720000 1.635000 ;
      RECT 136.240000  3.805000 136.720000 3.935000 ;
      RECT 136.240000  4.265000 136.410000 4.685000 ;
      RECT 136.240000  4.685000 136.680000 4.855000 ;
      RECT 136.245000  2.635000 137.915000 2.805000 ;
      RECT 136.390000  1.635000 136.720000 2.465000 ;
      RECT 136.390000  2.975000 136.720000 3.805000 ;
      RECT 136.430000  0.330000 136.680000 0.585000 ;
      RECT 136.430000  4.855000 136.680000 5.110000 ;
      RECT 136.585000  0.945000 136.985000 1.295000 ;
      RECT 136.585000  4.145000 136.985000 4.495000 ;
      RECT 136.915000  0.085000 137.245000 0.660000 ;
      RECT 136.915000  1.465000 137.245000 2.635000 ;
      RECT 136.915000  2.805000 137.245000 3.975000 ;
      RECT 136.915000  4.780000 137.245000 5.355000 ;
      RECT 137.175000  0.945000 137.575000 1.295000 ;
      RECT 137.175000  4.145000 137.575000 4.495000 ;
      RECT 137.440000  1.465000 138.140000 1.505000 ;
      RECT 137.440000  1.505000 137.920000 1.635000 ;
      RECT 137.440000  1.635000 137.770000 2.465000 ;
      RECT 137.440000  2.975000 137.770000 3.805000 ;
      RECT 137.440000  3.805000 137.920000 3.935000 ;
      RECT 137.440000  3.935000 138.140000 3.975000 ;
      RECT 137.480000  0.330000 137.730000 0.585000 ;
      RECT 137.480000  0.585000 137.920000 0.755000 ;
      RECT 137.480000  4.685000 137.920000 4.855000 ;
      RECT 137.480000  4.855000 137.730000 5.110000 ;
      RECT 137.750000  0.755000 137.920000 1.175000 ;
      RECT 137.750000  1.175000 138.140000 1.465000 ;
      RECT 137.750000  3.975000 138.140000 4.265000 ;
      RECT 137.750000  4.265000 137.920000 4.685000 ;
      RECT 137.960000  1.805000 138.480000 1.985000 ;
      RECT 137.960000  1.985000 138.290000 2.465000 ;
      RECT 137.960000  2.975000 138.290000 3.455000 ;
      RECT 137.960000  3.455000 138.480000 3.635000 ;
      RECT 138.085000  1.755000 138.480000 1.805000 ;
      RECT 138.085000  2.465000 138.290000 2.975000 ;
      RECT 138.085000  3.635000 138.480000 3.685000 ;
      RECT 138.090000  0.330000 138.335000 0.835000 ;
      RECT 138.090000  0.835000 138.480000 1.005000 ;
      RECT 138.090000  4.435000 138.480000 4.605000 ;
      RECT 138.090000  4.605000 138.335000 5.110000 ;
      RECT 138.310000  1.005000 138.480000 1.755000 ;
      RECT 138.310000  3.685000 138.480000 4.435000 ;
      RECT 138.460000  2.635000 139.840000 2.805000 ;
      RECT 138.545000  0.395000 138.820000 0.625000 ;
      RECT 138.545000  4.815000 138.820000 5.045000 ;
      RECT 138.650000  0.625000 138.820000 1.055000 ;
      RECT 138.650000  1.055000 139.045000 1.325000 ;
      RECT 138.650000  4.115000 139.045000 4.385000 ;
      RECT 138.650000  4.385000 138.820000 4.815000 ;
      RECT 138.955000  1.495000 139.345000 2.635000 ;
      RECT 138.955000  2.805000 139.345000 3.945000 ;
      RECT 138.990000  0.085000 139.310000 0.885000 ;
      RECT 138.990000  4.555000 139.310000 5.355000 ;
      RECT 139.255000  1.055000 139.650000 1.325000 ;
      RECT 139.255000  4.115000 139.650000 4.385000 ;
      RECT 139.480000  0.395000 139.755000 0.625000 ;
      RECT 139.480000  0.625000 139.650000 1.055000 ;
      RECT 139.480000  4.385000 139.650000 4.815000 ;
      RECT 139.480000  4.815000 139.755000 5.045000 ;
      RECT 139.820000  0.835000 140.210000 1.005000 ;
      RECT 139.820000  1.005000 139.990000 1.755000 ;
      RECT 139.820000  1.755000 140.215000 1.805000 ;
      RECT 139.820000  1.805000 140.340000 1.985000 ;
      RECT 139.820000  3.455000 140.340000 3.635000 ;
      RECT 139.820000  3.635000 140.215000 3.685000 ;
      RECT 139.820000  3.685000 139.990000 4.435000 ;
      RECT 139.820000  4.435000 140.210000 4.605000 ;
      RECT 139.965000  0.330000 140.210000 0.835000 ;
      RECT 139.965000  4.605000 140.210000 5.110000 ;
      RECT 140.010000  1.985000 140.340000 2.465000 ;
      RECT 140.010000  2.465000 140.215000 2.975000 ;
      RECT 140.010000  2.975000 140.340000 3.455000 ;
      RECT 140.160000  1.175000 140.550000 1.465000 ;
      RECT 140.160000  1.465000 140.860000 1.505000 ;
      RECT 140.160000  3.935000 140.860000 3.975000 ;
      RECT 140.160000  3.975000 140.550000 4.265000 ;
      RECT 140.380000  0.585000 140.820000 0.755000 ;
      RECT 140.380000  0.755000 140.550000 1.175000 ;
      RECT 140.380000  1.505000 140.860000 1.635000 ;
      RECT 140.380000  3.805000 140.860000 3.935000 ;
      RECT 140.380000  4.265000 140.550000 4.685000 ;
      RECT 140.380000  4.685000 140.820000 4.855000 ;
      RECT 140.385000  2.635000 142.055000 2.805000 ;
      RECT 140.530000  1.635000 140.860000 2.465000 ;
      RECT 140.530000  2.975000 140.860000 3.805000 ;
      RECT 140.570000  0.330000 140.820000 0.585000 ;
      RECT 140.570000  4.855000 140.820000 5.110000 ;
      RECT 140.725000  0.945000 141.125000 1.295000 ;
      RECT 140.725000  4.145000 141.125000 4.495000 ;
      RECT 141.055000  0.085000 141.385000 0.660000 ;
      RECT 141.055000  1.465000 141.385000 2.635000 ;
      RECT 141.055000  2.805000 141.385000 3.975000 ;
      RECT 141.055000  4.780000 141.385000 5.355000 ;
      RECT 141.315000  0.945000 141.715000 1.295000 ;
      RECT 141.315000  4.145000 141.715000 4.495000 ;
      RECT 141.580000  1.465000 142.280000 1.505000 ;
      RECT 141.580000  1.505000 142.060000 1.635000 ;
      RECT 141.580000  1.635000 141.910000 2.465000 ;
      RECT 141.580000  2.975000 141.910000 3.805000 ;
      RECT 141.580000  3.805000 142.060000 3.935000 ;
      RECT 141.580000  3.935000 142.280000 3.975000 ;
      RECT 141.620000  0.330000 141.870000 0.585000 ;
      RECT 141.620000  0.585000 142.060000 0.755000 ;
      RECT 141.620000  4.685000 142.060000 4.855000 ;
      RECT 141.620000  4.855000 141.870000 5.110000 ;
      RECT 141.890000  0.755000 142.060000 1.175000 ;
      RECT 141.890000  1.175000 142.280000 1.465000 ;
      RECT 141.890000  3.975000 142.280000 4.265000 ;
      RECT 141.890000  4.265000 142.060000 4.685000 ;
      RECT 142.100000  1.805000 142.620000 1.985000 ;
      RECT 142.100000  1.985000 142.430000 2.465000 ;
      RECT 142.100000  2.975000 142.430000 3.455000 ;
      RECT 142.100000  3.455000 142.620000 3.635000 ;
      RECT 142.225000  1.755000 142.620000 1.805000 ;
      RECT 142.225000  2.465000 142.430000 2.975000 ;
      RECT 142.225000  3.635000 142.620000 3.685000 ;
      RECT 142.230000  0.330000 142.475000 0.835000 ;
      RECT 142.230000  0.835000 142.620000 1.005000 ;
      RECT 142.230000  4.435000 142.620000 4.605000 ;
      RECT 142.230000  4.605000 142.475000 5.110000 ;
      RECT 142.450000  1.005000 142.620000 1.755000 ;
      RECT 142.450000  3.685000 142.620000 4.435000 ;
      RECT 142.600000  2.635000 143.980000 2.805000 ;
      RECT 142.685000  0.395000 142.960000 0.625000 ;
      RECT 142.685000  4.815000 142.960000 5.045000 ;
      RECT 142.790000  0.625000 142.960000 1.055000 ;
      RECT 142.790000  1.055000 143.185000 1.325000 ;
      RECT 142.790000  4.115000 143.185000 4.385000 ;
      RECT 142.790000  4.385000 142.960000 4.815000 ;
      RECT 143.095000  1.495000 143.485000 2.635000 ;
      RECT 143.095000  2.805000 143.485000 3.945000 ;
      RECT 143.130000  0.085000 143.450000 0.885000 ;
      RECT 143.130000  4.555000 143.450000 5.355000 ;
      RECT 143.395000  1.055000 143.790000 1.325000 ;
      RECT 143.395000  4.115000 143.790000 4.385000 ;
      RECT 143.620000  0.395000 143.895000 0.625000 ;
      RECT 143.620000  0.625000 143.790000 1.055000 ;
      RECT 143.620000  4.385000 143.790000 4.815000 ;
      RECT 143.620000  4.815000 143.895000 5.045000 ;
      RECT 143.960000  0.835000 144.350000 1.005000 ;
      RECT 143.960000  1.005000 144.130000 1.755000 ;
      RECT 143.960000  1.755000 144.355000 1.805000 ;
      RECT 143.960000  1.805000 144.480000 1.985000 ;
      RECT 143.960000  3.455000 144.480000 3.635000 ;
      RECT 143.960000  3.635000 144.355000 3.685000 ;
      RECT 143.960000  3.685000 144.130000 4.435000 ;
      RECT 143.960000  4.435000 144.350000 4.605000 ;
      RECT 144.105000  0.330000 144.350000 0.835000 ;
      RECT 144.105000  4.605000 144.350000 5.110000 ;
      RECT 144.150000  1.985000 144.480000 2.465000 ;
      RECT 144.150000  2.465000 144.355000 2.975000 ;
      RECT 144.150000  2.975000 144.480000 3.455000 ;
      RECT 144.300000  1.175000 144.690000 1.465000 ;
      RECT 144.300000  1.465000 145.000000 1.505000 ;
      RECT 144.300000  3.935000 145.000000 3.975000 ;
      RECT 144.300000  3.975000 144.690000 4.265000 ;
      RECT 144.520000  0.585000 144.960000 0.755000 ;
      RECT 144.520000  0.755000 144.690000 1.175000 ;
      RECT 144.520000  1.505000 145.000000 1.635000 ;
      RECT 144.520000  3.805000 145.000000 3.935000 ;
      RECT 144.520000  4.265000 144.690000 4.685000 ;
      RECT 144.520000  4.685000 144.960000 4.855000 ;
      RECT 144.525000  2.635000 146.195000 2.805000 ;
      RECT 144.670000  1.635000 145.000000 2.465000 ;
      RECT 144.670000  2.975000 145.000000 3.805000 ;
      RECT 144.710000  0.330000 144.960000 0.585000 ;
      RECT 144.710000  4.855000 144.960000 5.110000 ;
      RECT 144.865000  0.945000 145.265000 1.295000 ;
      RECT 144.865000  4.145000 145.265000 4.495000 ;
      RECT 145.195000  0.085000 145.525000 0.660000 ;
      RECT 145.195000  1.465000 145.525000 2.635000 ;
      RECT 145.195000  2.805000 145.525000 3.975000 ;
      RECT 145.195000  4.780000 145.525000 5.355000 ;
      RECT 145.455000  0.945000 145.855000 1.295000 ;
      RECT 145.455000  4.145000 145.855000 4.495000 ;
      RECT 145.720000  1.465000 146.420000 1.505000 ;
      RECT 145.720000  1.505000 146.200000 1.635000 ;
      RECT 145.720000  1.635000 146.050000 2.465000 ;
      RECT 145.720000  2.975000 146.050000 3.805000 ;
      RECT 145.720000  3.805000 146.200000 3.935000 ;
      RECT 145.720000  3.935000 146.420000 3.975000 ;
      RECT 145.760000  0.330000 146.010000 0.585000 ;
      RECT 145.760000  0.585000 146.200000 0.755000 ;
      RECT 145.760000  4.685000 146.200000 4.855000 ;
      RECT 145.760000  4.855000 146.010000 5.110000 ;
      RECT 146.030000  0.755000 146.200000 1.175000 ;
      RECT 146.030000  1.175000 146.420000 1.465000 ;
      RECT 146.030000  3.975000 146.420000 4.265000 ;
      RECT 146.030000  4.265000 146.200000 4.685000 ;
      RECT 146.240000  1.805000 146.760000 1.985000 ;
      RECT 146.240000  1.985000 146.570000 2.465000 ;
      RECT 146.240000  2.975000 146.570000 3.455000 ;
      RECT 146.240000  3.455000 146.760000 3.635000 ;
      RECT 146.365000  1.755000 146.760000 1.805000 ;
      RECT 146.365000  2.465000 146.570000 2.975000 ;
      RECT 146.365000  3.635000 146.760000 3.685000 ;
      RECT 146.370000  0.330000 146.615000 0.835000 ;
      RECT 146.370000  0.835000 146.760000 1.005000 ;
      RECT 146.370000  4.435000 146.760000 4.605000 ;
      RECT 146.370000  4.605000 146.615000 5.110000 ;
      RECT 146.590000  1.005000 146.760000 1.755000 ;
      RECT 146.590000  3.685000 146.760000 4.435000 ;
      RECT 146.740000  2.635000 149.075000 2.805000 ;
      RECT 146.825000  0.395000 147.100000 0.625000 ;
      RECT 146.825000  4.815000 147.100000 5.045000 ;
      RECT 146.930000  0.625000 147.100000 1.055000 ;
      RECT 146.930000  1.055000 147.325000 1.325000 ;
      RECT 146.930000  4.115000 147.325000 4.385000 ;
      RECT 146.930000  4.385000 147.100000 4.815000 ;
      RECT 147.235000  1.495000 147.565000 2.635000 ;
      RECT 147.235000  2.805000 147.565000 3.945000 ;
      RECT 147.270000  0.085000 147.530000 0.885000 ;
      RECT 147.270000  4.555000 147.530000 5.355000 ;
      RECT 147.755000  1.055000 148.575000 1.325000 ;
      RECT 147.755000  1.495000 148.945000 1.665000 ;
      RECT 147.755000  1.665000 148.055000 2.210000 ;
      RECT 147.755000  2.210000 148.085000 2.465000 ;
      RECT 147.755000  2.975000 148.085000 3.230000 ;
      RECT 147.755000  3.230000 148.055000 3.775000 ;
      RECT 147.755000  3.775000 148.945000 3.945000 ;
      RECT 147.755000  4.115000 148.575000 4.385000 ;
      RECT 147.805000  0.255000 148.135000 0.715000 ;
      RECT 147.805000  0.715000 148.995000 0.885000 ;
      RECT 147.805000  4.555000 148.995000 4.725000 ;
      RECT 147.805000  4.725000 148.135000 5.185000 ;
      RECT 148.225000  1.835000 148.555000 2.105000 ;
      RECT 148.225000  3.335000 148.555000 3.605000 ;
      RECT 148.255000  2.105000 148.555000 2.635000 ;
      RECT 148.255000  2.805000 148.555000 3.335000 ;
      RECT 148.305000  0.085000 148.520000 0.545000 ;
      RECT 148.305000  4.895000 148.520000 5.355000 ;
      RECT 148.690000  0.255000 149.835000 0.425000 ;
      RECT 148.690000  0.425000 148.995000 0.715000 ;
      RECT 148.690000  0.885000 148.995000 0.925000 ;
      RECT 148.690000  4.515000 148.995000 4.555000 ;
      RECT 148.690000  4.725000 148.995000 5.015000 ;
      RECT 148.690000  5.015000 149.835000 5.185000 ;
      RECT 148.775000  1.665000 148.945000 2.295000 ;
      RECT 148.775000  2.295000 149.075000 2.465000 ;
      RECT 148.775000  2.975000 149.075000 3.145000 ;
      RECT 148.775000  3.145000 148.945000 3.775000 ;
      RECT 149.125000  1.755000 149.555000 2.125000 ;
      RECT 149.125000  3.315000 149.555000 3.685000 ;
      RECT 149.165000  0.595000 149.495000 0.885000 ;
      RECT 149.165000  4.555000 149.495000 4.845000 ;
      RECT 149.245000  0.885000 149.415000 1.755000 ;
      RECT 149.245000  2.125000 149.415000 3.315000 ;
      RECT 149.245000  3.685000 149.415000 4.555000 ;
      RECT 149.585000  2.295000 149.940000 2.465000 ;
      RECT 149.585000  2.635000 152.175000 2.805000 ;
      RECT 149.585000  2.975000 149.940000 3.145000 ;
      RECT 149.665000  0.425000 149.835000 0.770000 ;
      RECT 149.665000  4.670000 149.835000 5.015000 ;
      RECT 149.760000  1.205000 150.175000 1.305000 ;
      RECT 149.760000  1.305000 150.280000 1.465000 ;
      RECT 149.760000  1.465000 150.540000 1.475000 ;
      RECT 149.760000  3.965000 150.540000 3.975000 ;
      RECT 149.760000  3.975000 150.280000 4.135000 ;
      RECT 149.760000  4.135000 150.175000 4.235000 ;
      RECT 149.770000  1.645000 149.940000 2.295000 ;
      RECT 149.770000  3.145000 149.940000 3.795000 ;
      RECT 150.005000  0.585000 150.585000 0.755000 ;
      RECT 150.005000  0.755000 150.175000 1.205000 ;
      RECT 150.005000  4.235000 150.175000 4.685000 ;
      RECT 150.005000  4.685000 150.585000 4.855000 ;
      RECT 150.110000  1.475000 150.540000 1.635000 ;
      RECT 150.110000  3.805000 150.540000 3.965000 ;
      RECT 150.210000  1.635000 150.540000 2.465000 ;
      RECT 150.210000  2.975000 150.540000 3.805000 ;
      RECT 150.335000  0.330000 150.585000 0.585000 ;
      RECT 150.335000  4.855000 150.585000 5.110000 ;
      RECT 150.450000  1.025000 150.785000 1.295000 ;
      RECT 150.450000  4.145000 150.785000 4.415000 ;
      RECT 150.715000  1.465000 151.045000 2.635000 ;
      RECT 150.715000  2.805000 151.045000 3.975000 ;
      RECT 150.755000  0.085000 151.005000 0.660000 ;
      RECT 150.755000  4.780000 151.005000 5.355000 ;
      RECT 150.975000  1.025000 151.310000 1.295000 ;
      RECT 150.975000  4.145000 151.310000 4.415000 ;
      RECT 151.175000  0.330000 151.425000 0.585000 ;
      RECT 151.175000  0.585000 151.755000 0.755000 ;
      RECT 151.175000  4.685000 151.755000 4.855000 ;
      RECT 151.175000  4.855000 151.425000 5.110000 ;
      RECT 151.220000  1.465000 152.000000 1.475000 ;
      RECT 151.220000  1.475000 151.650000 1.635000 ;
      RECT 151.220000  1.635000 151.550000 2.465000 ;
      RECT 151.220000  2.975000 151.550000 3.805000 ;
      RECT 151.220000  3.805000 151.650000 3.965000 ;
      RECT 151.220000  3.965000 152.000000 3.975000 ;
      RECT 151.480000  1.305000 152.000000 1.465000 ;
      RECT 151.480000  3.975000 152.000000 4.135000 ;
      RECT 151.585000  0.755000 151.755000 1.205000 ;
      RECT 151.585000  1.205000 152.000000 1.305000 ;
      RECT 151.585000  4.135000 152.000000 4.235000 ;
      RECT 151.585000  4.235000 151.755000 4.685000 ;
      RECT 151.820000  1.645000 151.990000 2.295000 ;
      RECT 151.820000  2.295000 152.175000 2.465000 ;
      RECT 151.820000  2.975000 152.175000 3.145000 ;
      RECT 151.820000  3.145000 151.990000 3.795000 ;
      RECT 151.925000  0.255000 153.070000 0.425000 ;
      RECT 151.925000  0.425000 152.095000 0.770000 ;
      RECT 151.925000  4.670000 152.095000 5.015000 ;
      RECT 151.925000  5.015000 153.070000 5.185000 ;
      RECT 152.205000  1.755000 152.635000 2.125000 ;
      RECT 152.205000  3.315000 152.635000 3.685000 ;
      RECT 152.265000  0.595000 152.595000 0.885000 ;
      RECT 152.265000  4.555000 152.595000 4.845000 ;
      RECT 152.345000  0.885000 152.515000 1.755000 ;
      RECT 152.345000  2.125000 152.515000 3.315000 ;
      RECT 152.345000  3.685000 152.515000 4.555000 ;
      RECT 152.685000  2.295000 152.985000 2.465000 ;
      RECT 152.685000  2.635000 155.515000 2.805000 ;
      RECT 152.685000  2.975000 152.985000 3.145000 ;
      RECT 152.765000  0.425000 153.070000 0.715000 ;
      RECT 152.765000  0.715000 153.955000 0.885000 ;
      RECT 152.765000  0.885000 153.070000 0.925000 ;
      RECT 152.765000  4.515000 153.070000 4.555000 ;
      RECT 152.765000  4.555000 153.955000 4.725000 ;
      RECT 152.765000  4.725000 153.070000 5.015000 ;
      RECT 152.815000  1.495000 154.005000 1.665000 ;
      RECT 152.815000  1.665000 152.985000 2.295000 ;
      RECT 152.815000  3.145000 152.985000 3.775000 ;
      RECT 152.815000  3.775000 154.005000 3.945000 ;
      RECT 153.185000  1.055000 154.005000 1.325000 ;
      RECT 153.185000  4.115000 154.005000 4.385000 ;
      RECT 153.205000  1.835000 153.535000 2.105000 ;
      RECT 153.205000  2.105000 153.505000 2.635000 ;
      RECT 153.205000  2.805000 153.505000 3.335000 ;
      RECT 153.205000  3.335000 153.535000 3.605000 ;
      RECT 153.240000  0.085000 153.455000 0.545000 ;
      RECT 153.240000  4.895000 153.455000 5.355000 ;
      RECT 153.625000  0.255000 153.955000 0.715000 ;
      RECT 153.625000  4.725000 153.955000 5.185000 ;
      RECT 153.675000  2.210000 154.005000 2.465000 ;
      RECT 153.675000  2.975000 154.005000 3.230000 ;
      RECT 153.705000  1.665000 154.005000 2.210000 ;
      RECT 153.705000  3.230000 154.005000 3.775000 ;
      RECT 154.195000  1.055000 155.015000 1.325000 ;
      RECT 154.195000  1.495000 155.385000 1.665000 ;
      RECT 154.195000  1.665000 154.495000 2.210000 ;
      RECT 154.195000  2.210000 154.525000 2.465000 ;
      RECT 154.195000  2.975000 154.525000 3.230000 ;
      RECT 154.195000  3.230000 154.495000 3.775000 ;
      RECT 154.195000  3.775000 155.385000 3.945000 ;
      RECT 154.195000  4.115000 155.015000 4.385000 ;
      RECT 154.245000  0.255000 154.575000 0.715000 ;
      RECT 154.245000  0.715000 155.435000 0.885000 ;
      RECT 154.245000  4.555000 155.435000 4.725000 ;
      RECT 154.245000  4.725000 154.575000 5.185000 ;
      RECT 154.665000  1.835000 154.995000 2.105000 ;
      RECT 154.665000  3.335000 154.995000 3.605000 ;
      RECT 154.695000  2.105000 154.995000 2.635000 ;
      RECT 154.695000  2.805000 154.995000 3.335000 ;
      RECT 154.745000  0.085000 154.960000 0.545000 ;
      RECT 154.745000  4.895000 154.960000 5.355000 ;
      RECT 155.130000  0.255000 156.275000 0.425000 ;
      RECT 155.130000  0.425000 155.435000 0.715000 ;
      RECT 155.130000  0.885000 155.435000 0.925000 ;
      RECT 155.130000  4.515000 155.435000 4.555000 ;
      RECT 155.130000  4.725000 155.435000 5.015000 ;
      RECT 155.130000  5.015000 156.275000 5.185000 ;
      RECT 155.215000  1.665000 155.385000 2.295000 ;
      RECT 155.215000  2.295000 155.515000 2.465000 ;
      RECT 155.215000  2.975000 155.515000 3.145000 ;
      RECT 155.215000  3.145000 155.385000 3.775000 ;
      RECT 155.565000  1.755000 155.995000 2.125000 ;
      RECT 155.565000  3.315000 155.995000 3.685000 ;
      RECT 155.605000  0.595000 155.935000 0.885000 ;
      RECT 155.605000  4.555000 155.935000 4.845000 ;
      RECT 155.685000  0.885000 155.855000 1.755000 ;
      RECT 155.685000  2.125000 155.855000 3.315000 ;
      RECT 155.685000  3.685000 155.855000 4.555000 ;
      RECT 156.025000  2.295000 156.380000 2.465000 ;
      RECT 156.025000  2.635000 158.615000 2.805000 ;
      RECT 156.025000  2.975000 156.380000 3.145000 ;
      RECT 156.105000  0.425000 156.275000 0.770000 ;
      RECT 156.105000  4.670000 156.275000 5.015000 ;
      RECT 156.200000  1.205000 156.615000 1.305000 ;
      RECT 156.200000  1.305000 156.720000 1.465000 ;
      RECT 156.200000  1.465000 156.980000 1.475000 ;
      RECT 156.200000  3.965000 156.980000 3.975000 ;
      RECT 156.200000  3.975000 156.720000 4.135000 ;
      RECT 156.200000  4.135000 156.615000 4.235000 ;
      RECT 156.210000  1.645000 156.380000 2.295000 ;
      RECT 156.210000  3.145000 156.380000 3.795000 ;
      RECT 156.445000  0.585000 157.025000 0.755000 ;
      RECT 156.445000  0.755000 156.615000 1.205000 ;
      RECT 156.445000  4.235000 156.615000 4.685000 ;
      RECT 156.445000  4.685000 157.025000 4.855000 ;
      RECT 156.550000  1.475000 156.980000 1.635000 ;
      RECT 156.550000  3.805000 156.980000 3.965000 ;
      RECT 156.650000  1.635000 156.980000 2.465000 ;
      RECT 156.650000  2.975000 156.980000 3.805000 ;
      RECT 156.775000  0.330000 157.025000 0.585000 ;
      RECT 156.775000  4.855000 157.025000 5.110000 ;
      RECT 156.890000  1.025000 157.225000 1.295000 ;
      RECT 156.890000  4.145000 157.225000 4.415000 ;
      RECT 157.155000  1.465000 157.485000 2.635000 ;
      RECT 157.155000  2.805000 157.485000 3.975000 ;
      RECT 157.195000  0.085000 157.445000 0.660000 ;
      RECT 157.195000  4.780000 157.445000 5.355000 ;
      RECT 157.415000  1.025000 157.750000 1.295000 ;
      RECT 157.415000  4.145000 157.750000 4.415000 ;
      RECT 157.615000  0.330000 157.865000 0.585000 ;
      RECT 157.615000  0.585000 158.195000 0.755000 ;
      RECT 157.615000  4.685000 158.195000 4.855000 ;
      RECT 157.615000  4.855000 157.865000 5.110000 ;
      RECT 157.660000  1.465000 158.440000 1.475000 ;
      RECT 157.660000  1.475000 158.090000 1.635000 ;
      RECT 157.660000  1.635000 157.990000 2.465000 ;
      RECT 157.660000  2.975000 157.990000 3.805000 ;
      RECT 157.660000  3.805000 158.090000 3.965000 ;
      RECT 157.660000  3.965000 158.440000 3.975000 ;
      RECT 157.920000  1.305000 158.440000 1.465000 ;
      RECT 157.920000  3.975000 158.440000 4.135000 ;
      RECT 158.025000  0.755000 158.195000 1.205000 ;
      RECT 158.025000  1.205000 158.440000 1.305000 ;
      RECT 158.025000  4.135000 158.440000 4.235000 ;
      RECT 158.025000  4.235000 158.195000 4.685000 ;
      RECT 158.260000  1.645000 158.430000 2.295000 ;
      RECT 158.260000  2.295000 158.615000 2.465000 ;
      RECT 158.260000  2.975000 158.615000 3.145000 ;
      RECT 158.260000  3.145000 158.430000 3.795000 ;
      RECT 158.365000  0.255000 159.510000 0.425000 ;
      RECT 158.365000  0.425000 158.535000 0.770000 ;
      RECT 158.365000  4.670000 158.535000 5.015000 ;
      RECT 158.365000  5.015000 159.510000 5.185000 ;
      RECT 158.645000  1.755000 159.075000 2.125000 ;
      RECT 158.645000  3.315000 159.075000 3.685000 ;
      RECT 158.705000  0.595000 159.035000 0.885000 ;
      RECT 158.705000  4.555000 159.035000 4.845000 ;
      RECT 158.785000  0.885000 158.955000 1.755000 ;
      RECT 158.785000  2.125000 158.955000 3.315000 ;
      RECT 158.785000  3.685000 158.955000 4.555000 ;
      RECT 159.125000  2.295000 159.425000 2.465000 ;
      RECT 159.125000  2.635000 161.955000 2.805000 ;
      RECT 159.125000  2.975000 159.425000 3.145000 ;
      RECT 159.205000  0.425000 159.510000 0.715000 ;
      RECT 159.205000  0.715000 160.395000 0.885000 ;
      RECT 159.205000  0.885000 159.510000 0.925000 ;
      RECT 159.205000  4.515000 159.510000 4.555000 ;
      RECT 159.205000  4.555000 160.395000 4.725000 ;
      RECT 159.205000  4.725000 159.510000 5.015000 ;
      RECT 159.255000  1.495000 160.445000 1.665000 ;
      RECT 159.255000  1.665000 159.425000 2.295000 ;
      RECT 159.255000  3.145000 159.425000 3.775000 ;
      RECT 159.255000  3.775000 160.445000 3.945000 ;
      RECT 159.625000  1.055000 160.445000 1.325000 ;
      RECT 159.625000  4.115000 160.445000 4.385000 ;
      RECT 159.645000  1.835000 159.975000 2.105000 ;
      RECT 159.645000  2.105000 159.945000 2.635000 ;
      RECT 159.645000  2.805000 159.945000 3.335000 ;
      RECT 159.645000  3.335000 159.975000 3.605000 ;
      RECT 159.680000  0.085000 159.895000 0.545000 ;
      RECT 159.680000  4.895000 159.895000 5.355000 ;
      RECT 160.065000  0.255000 160.395000 0.715000 ;
      RECT 160.065000  4.725000 160.395000 5.185000 ;
      RECT 160.115000  2.210000 160.445000 2.465000 ;
      RECT 160.115000  2.975000 160.445000 3.230000 ;
      RECT 160.145000  1.665000 160.445000 2.210000 ;
      RECT 160.145000  3.230000 160.445000 3.775000 ;
      RECT 160.635000  1.055000 161.455000 1.325000 ;
      RECT 160.635000  1.495000 161.825000 1.665000 ;
      RECT 160.635000  1.665000 160.935000 2.210000 ;
      RECT 160.635000  2.210000 160.965000 2.465000 ;
      RECT 160.635000  2.975000 160.965000 3.230000 ;
      RECT 160.635000  3.230000 160.935000 3.775000 ;
      RECT 160.635000  3.775000 161.825000 3.945000 ;
      RECT 160.635000  4.115000 161.455000 4.385000 ;
      RECT 160.685000  0.255000 161.015000 0.715000 ;
      RECT 160.685000  0.715000 161.875000 0.885000 ;
      RECT 160.685000  4.555000 161.875000 4.725000 ;
      RECT 160.685000  4.725000 161.015000 5.185000 ;
      RECT 161.105000  1.835000 161.435000 2.105000 ;
      RECT 161.105000  3.335000 161.435000 3.605000 ;
      RECT 161.135000  2.105000 161.435000 2.635000 ;
      RECT 161.135000  2.805000 161.435000 3.335000 ;
      RECT 161.185000  0.085000 161.400000 0.545000 ;
      RECT 161.185000  4.895000 161.400000 5.355000 ;
      RECT 161.570000  0.255000 162.715000 0.425000 ;
      RECT 161.570000  0.425000 161.875000 0.715000 ;
      RECT 161.570000  0.885000 161.875000 0.925000 ;
      RECT 161.570000  4.515000 161.875000 4.555000 ;
      RECT 161.570000  4.725000 161.875000 5.015000 ;
      RECT 161.570000  5.015000 162.715000 5.185000 ;
      RECT 161.655000  1.665000 161.825000 2.295000 ;
      RECT 161.655000  2.295000 161.955000 2.465000 ;
      RECT 161.655000  2.975000 161.955000 3.145000 ;
      RECT 161.655000  3.145000 161.825000 3.775000 ;
      RECT 162.005000  1.755000 162.435000 2.125000 ;
      RECT 162.005000  3.315000 162.435000 3.685000 ;
      RECT 162.045000  0.595000 162.375000 0.885000 ;
      RECT 162.045000  4.555000 162.375000 4.845000 ;
      RECT 162.125000  0.885000 162.295000 1.755000 ;
      RECT 162.125000  2.125000 162.295000 3.315000 ;
      RECT 162.125000  3.685000 162.295000 4.555000 ;
      RECT 162.465000  2.295000 162.820000 2.465000 ;
      RECT 162.465000  2.635000 165.055000 2.805000 ;
      RECT 162.465000  2.975000 162.820000 3.145000 ;
      RECT 162.545000  0.425000 162.715000 0.770000 ;
      RECT 162.545000  4.670000 162.715000 5.015000 ;
      RECT 162.640000  1.205000 163.055000 1.305000 ;
      RECT 162.640000  1.305000 163.160000 1.465000 ;
      RECT 162.640000  1.465000 163.420000 1.475000 ;
      RECT 162.640000  3.965000 163.420000 3.975000 ;
      RECT 162.640000  3.975000 163.160000 4.135000 ;
      RECT 162.640000  4.135000 163.055000 4.235000 ;
      RECT 162.650000  1.645000 162.820000 2.295000 ;
      RECT 162.650000  3.145000 162.820000 3.795000 ;
      RECT 162.885000  0.585000 163.465000 0.755000 ;
      RECT 162.885000  0.755000 163.055000 1.205000 ;
      RECT 162.885000  4.235000 163.055000 4.685000 ;
      RECT 162.885000  4.685000 163.465000 4.855000 ;
      RECT 162.990000  1.475000 163.420000 1.635000 ;
      RECT 162.990000  3.805000 163.420000 3.965000 ;
      RECT 163.090000  1.635000 163.420000 2.465000 ;
      RECT 163.090000  2.975000 163.420000 3.805000 ;
      RECT 163.215000  0.330000 163.465000 0.585000 ;
      RECT 163.215000  4.855000 163.465000 5.110000 ;
      RECT 163.330000  1.025000 163.665000 1.295000 ;
      RECT 163.330000  4.145000 163.665000 4.415000 ;
      RECT 163.595000  1.465000 163.925000 2.635000 ;
      RECT 163.595000  2.805000 163.925000 3.975000 ;
      RECT 163.635000  0.085000 163.885000 0.660000 ;
      RECT 163.635000  4.780000 163.885000 5.355000 ;
      RECT 163.855000  1.025000 164.190000 1.295000 ;
      RECT 163.855000  4.145000 164.190000 4.415000 ;
      RECT 164.055000  0.330000 164.305000 0.585000 ;
      RECT 164.055000  0.585000 164.635000 0.755000 ;
      RECT 164.055000  4.685000 164.635000 4.855000 ;
      RECT 164.055000  4.855000 164.305000 5.110000 ;
      RECT 164.100000  1.465000 164.880000 1.475000 ;
      RECT 164.100000  1.475000 164.530000 1.635000 ;
      RECT 164.100000  1.635000 164.430000 2.465000 ;
      RECT 164.100000  2.975000 164.430000 3.805000 ;
      RECT 164.100000  3.805000 164.530000 3.965000 ;
      RECT 164.100000  3.965000 164.880000 3.975000 ;
      RECT 164.360000  1.305000 164.880000 1.465000 ;
      RECT 164.360000  3.975000 164.880000 4.135000 ;
      RECT 164.465000  0.755000 164.635000 1.205000 ;
      RECT 164.465000  1.205000 164.880000 1.305000 ;
      RECT 164.465000  4.135000 164.880000 4.235000 ;
      RECT 164.465000  4.235000 164.635000 4.685000 ;
      RECT 164.700000  1.645000 164.870000 2.295000 ;
      RECT 164.700000  2.295000 165.055000 2.465000 ;
      RECT 164.700000  2.975000 165.055000 3.145000 ;
      RECT 164.700000  3.145000 164.870000 3.795000 ;
      RECT 164.805000  0.255000 165.950000 0.425000 ;
      RECT 164.805000  0.425000 164.975000 0.770000 ;
      RECT 164.805000  4.670000 164.975000 5.015000 ;
      RECT 164.805000  5.015000 165.950000 5.185000 ;
      RECT 165.085000  1.755000 165.515000 2.125000 ;
      RECT 165.085000  3.315000 165.515000 3.685000 ;
      RECT 165.145000  0.595000 165.475000 0.885000 ;
      RECT 165.145000  4.555000 165.475000 4.845000 ;
      RECT 165.225000  0.885000 165.395000 1.755000 ;
      RECT 165.225000  2.125000 165.395000 3.315000 ;
      RECT 165.225000  3.685000 165.395000 4.555000 ;
      RECT 165.565000  2.295000 165.865000 2.465000 ;
      RECT 165.565000  2.635000 168.395000 2.805000 ;
      RECT 165.565000  2.975000 165.865000 3.145000 ;
      RECT 165.645000  0.425000 165.950000 0.715000 ;
      RECT 165.645000  0.715000 166.835000 0.885000 ;
      RECT 165.645000  0.885000 165.950000 0.925000 ;
      RECT 165.645000  4.515000 165.950000 4.555000 ;
      RECT 165.645000  4.555000 166.835000 4.725000 ;
      RECT 165.645000  4.725000 165.950000 5.015000 ;
      RECT 165.695000  1.495000 166.885000 1.665000 ;
      RECT 165.695000  1.665000 165.865000 2.295000 ;
      RECT 165.695000  3.145000 165.865000 3.775000 ;
      RECT 165.695000  3.775000 166.885000 3.945000 ;
      RECT 166.065000  1.055000 166.885000 1.325000 ;
      RECT 166.065000  4.115000 166.885000 4.385000 ;
      RECT 166.085000  1.835000 166.415000 2.105000 ;
      RECT 166.085000  2.105000 166.385000 2.635000 ;
      RECT 166.085000  2.805000 166.385000 3.335000 ;
      RECT 166.085000  3.335000 166.415000 3.605000 ;
      RECT 166.120000  0.085000 166.335000 0.545000 ;
      RECT 166.120000  4.895000 166.335000 5.355000 ;
      RECT 166.505000  0.255000 166.835000 0.715000 ;
      RECT 166.505000  4.725000 166.835000 5.185000 ;
      RECT 166.555000  2.210000 166.885000 2.465000 ;
      RECT 166.555000  2.975000 166.885000 3.230000 ;
      RECT 166.585000  1.665000 166.885000 2.210000 ;
      RECT 166.585000  3.230000 166.885000 3.775000 ;
      RECT 167.075000  1.055000 167.895000 1.325000 ;
      RECT 167.075000  1.495000 168.265000 1.665000 ;
      RECT 167.075000  1.665000 167.375000 2.210000 ;
      RECT 167.075000  2.210000 167.405000 2.465000 ;
      RECT 167.075000  2.975000 167.405000 3.230000 ;
      RECT 167.075000  3.230000 167.375000 3.775000 ;
      RECT 167.075000  3.775000 168.265000 3.945000 ;
      RECT 167.075000  4.115000 167.895000 4.385000 ;
      RECT 167.125000  0.255000 167.455000 0.715000 ;
      RECT 167.125000  0.715000 168.315000 0.885000 ;
      RECT 167.125000  4.555000 168.315000 4.725000 ;
      RECT 167.125000  4.725000 167.455000 5.185000 ;
      RECT 167.545000  1.835000 167.875000 2.105000 ;
      RECT 167.545000  3.335000 167.875000 3.605000 ;
      RECT 167.575000  2.105000 167.875000 2.635000 ;
      RECT 167.575000  2.805000 167.875000 3.335000 ;
      RECT 167.625000  0.085000 167.840000 0.545000 ;
      RECT 167.625000  4.895000 167.840000 5.355000 ;
      RECT 168.010000  0.255000 169.155000 0.425000 ;
      RECT 168.010000  0.425000 168.315000 0.715000 ;
      RECT 168.010000  0.885000 168.315000 0.925000 ;
      RECT 168.010000  4.515000 168.315000 4.555000 ;
      RECT 168.010000  4.725000 168.315000 5.015000 ;
      RECT 168.010000  5.015000 169.155000 5.185000 ;
      RECT 168.095000  1.665000 168.265000 2.295000 ;
      RECT 168.095000  2.295000 168.395000 2.465000 ;
      RECT 168.095000  2.975000 168.395000 3.145000 ;
      RECT 168.095000  3.145000 168.265000 3.775000 ;
      RECT 168.445000  1.755000 168.875000 2.125000 ;
      RECT 168.445000  3.315000 168.875000 3.685000 ;
      RECT 168.485000  0.595000 168.815000 0.885000 ;
      RECT 168.485000  4.555000 168.815000 4.845000 ;
      RECT 168.565000  0.885000 168.735000 1.755000 ;
      RECT 168.565000  2.125000 168.735000 3.315000 ;
      RECT 168.565000  3.685000 168.735000 4.555000 ;
      RECT 168.905000  2.295000 169.260000 2.465000 ;
      RECT 168.905000  2.635000 171.495000 2.805000 ;
      RECT 168.905000  2.975000 169.260000 3.145000 ;
      RECT 168.985000  0.425000 169.155000 0.770000 ;
      RECT 168.985000  4.670000 169.155000 5.015000 ;
      RECT 169.080000  1.205000 169.495000 1.305000 ;
      RECT 169.080000  1.305000 169.600000 1.465000 ;
      RECT 169.080000  1.465000 169.860000 1.475000 ;
      RECT 169.080000  3.965000 169.860000 3.975000 ;
      RECT 169.080000  3.975000 169.600000 4.135000 ;
      RECT 169.080000  4.135000 169.495000 4.235000 ;
      RECT 169.090000  1.645000 169.260000 2.295000 ;
      RECT 169.090000  3.145000 169.260000 3.795000 ;
      RECT 169.325000  0.585000 169.905000 0.755000 ;
      RECT 169.325000  0.755000 169.495000 1.205000 ;
      RECT 169.325000  4.235000 169.495000 4.685000 ;
      RECT 169.325000  4.685000 169.905000 4.855000 ;
      RECT 169.430000  1.475000 169.860000 1.635000 ;
      RECT 169.430000  3.805000 169.860000 3.965000 ;
      RECT 169.530000  1.635000 169.860000 2.465000 ;
      RECT 169.530000  2.975000 169.860000 3.805000 ;
      RECT 169.655000  0.330000 169.905000 0.585000 ;
      RECT 169.655000  4.855000 169.905000 5.110000 ;
      RECT 169.770000  1.025000 170.105000 1.295000 ;
      RECT 169.770000  4.145000 170.105000 4.415000 ;
      RECT 170.035000  1.465000 170.365000 2.635000 ;
      RECT 170.035000  2.805000 170.365000 3.975000 ;
      RECT 170.075000  0.085000 170.325000 0.660000 ;
      RECT 170.075000  4.780000 170.325000 5.355000 ;
      RECT 170.295000  1.025000 170.630000 1.295000 ;
      RECT 170.295000  4.145000 170.630000 4.415000 ;
      RECT 170.495000  0.330000 170.745000 0.585000 ;
      RECT 170.495000  0.585000 171.075000 0.755000 ;
      RECT 170.495000  4.685000 171.075000 4.855000 ;
      RECT 170.495000  4.855000 170.745000 5.110000 ;
      RECT 170.540000  1.465000 171.320000 1.475000 ;
      RECT 170.540000  1.475000 170.970000 1.635000 ;
      RECT 170.540000  1.635000 170.870000 2.465000 ;
      RECT 170.540000  2.975000 170.870000 3.805000 ;
      RECT 170.540000  3.805000 170.970000 3.965000 ;
      RECT 170.540000  3.965000 171.320000 3.975000 ;
      RECT 170.800000  1.305000 171.320000 1.465000 ;
      RECT 170.800000  3.975000 171.320000 4.135000 ;
      RECT 170.905000  0.755000 171.075000 1.205000 ;
      RECT 170.905000  1.205000 171.320000 1.305000 ;
      RECT 170.905000  4.135000 171.320000 4.235000 ;
      RECT 170.905000  4.235000 171.075000 4.685000 ;
      RECT 171.140000  1.645000 171.310000 2.295000 ;
      RECT 171.140000  2.295000 171.495000 2.465000 ;
      RECT 171.140000  2.975000 171.495000 3.145000 ;
      RECT 171.140000  3.145000 171.310000 3.795000 ;
      RECT 171.245000  0.255000 172.390000 0.425000 ;
      RECT 171.245000  0.425000 171.415000 0.770000 ;
      RECT 171.245000  4.670000 171.415000 5.015000 ;
      RECT 171.245000  5.015000 172.390000 5.185000 ;
      RECT 171.525000  1.755000 171.955000 2.125000 ;
      RECT 171.525000  3.315000 171.955000 3.685000 ;
      RECT 171.585000  0.595000 171.915000 0.885000 ;
      RECT 171.585000  4.555000 171.915000 4.845000 ;
      RECT 171.665000  0.885000 171.835000 1.755000 ;
      RECT 171.665000  2.125000 171.835000 3.315000 ;
      RECT 171.665000  3.685000 171.835000 4.555000 ;
      RECT 172.005000  2.295000 172.305000 2.465000 ;
      RECT 172.005000  2.635000 176.215000 2.805000 ;
      RECT 172.005000  2.975000 172.305000 3.145000 ;
      RECT 172.085000  0.425000 172.390000 0.715000 ;
      RECT 172.085000  0.715000 173.275000 0.885000 ;
      RECT 172.085000  0.885000 172.390000 0.925000 ;
      RECT 172.085000  4.515000 172.390000 4.555000 ;
      RECT 172.085000  4.555000 173.275000 4.725000 ;
      RECT 172.085000  4.725000 172.390000 5.015000 ;
      RECT 172.135000  1.495000 173.325000 1.665000 ;
      RECT 172.135000  1.665000 172.305000 2.295000 ;
      RECT 172.135000  3.145000 172.305000 3.775000 ;
      RECT 172.135000  3.775000 173.325000 3.945000 ;
      RECT 172.505000  1.055000 173.325000 1.325000 ;
      RECT 172.505000  4.115000 173.325000 4.385000 ;
      RECT 172.525000  1.835000 172.855000 2.105000 ;
      RECT 172.525000  2.105000 172.825000 2.635000 ;
      RECT 172.525000  2.805000 172.825000 3.335000 ;
      RECT 172.525000  3.335000 172.855000 3.605000 ;
      RECT 172.560000  0.085000 172.775000 0.545000 ;
      RECT 172.560000  4.895000 172.775000 5.355000 ;
      RECT 172.945000  0.255000 173.275000 0.715000 ;
      RECT 172.945000  4.725000 173.275000 5.185000 ;
      RECT 172.995000  2.210000 173.325000 2.465000 ;
      RECT 172.995000  2.975000 173.325000 3.230000 ;
      RECT 173.025000  1.665000 173.325000 2.210000 ;
      RECT 173.025000  3.230000 173.325000 3.775000 ;
      RECT 173.545000  1.495000 173.815000 2.635000 ;
      RECT 173.545000  2.805000 173.815000 3.945000 ;
      RECT 173.565000  0.085000 173.815000 0.885000 ;
      RECT 173.565000  4.555000 173.815000 5.355000 ;
      RECT 173.815000  1.055000 175.205000 1.325000 ;
      RECT 173.815000  4.115000 175.205000 4.385000 ;
      RECT 173.985000  0.255000 174.315000 0.715000 ;
      RECT 173.985000  0.715000 176.115000 0.885000 ;
      RECT 173.985000  1.495000 176.215000 1.665000 ;
      RECT 173.985000  1.665000 174.315000 2.465000 ;
      RECT 173.985000  2.975000 174.315000 3.775000 ;
      RECT 173.985000  3.775000 176.215000 3.945000 ;
      RECT 173.985000  4.555000 176.115000 4.725000 ;
      RECT 173.985000  4.725000 174.315000 5.185000 ;
      RECT 174.485000  0.085000 174.755000 0.545000 ;
      RECT 174.485000  1.835000 174.755000 2.635000 ;
      RECT 174.485000  2.805000 174.755000 3.605000 ;
      RECT 174.485000  4.895000 174.755000 5.355000 ;
      RECT 174.925000  0.255000 175.255000 0.715000 ;
      RECT 174.925000  1.665000 175.255000 2.465000 ;
      RECT 174.925000  2.975000 175.255000 3.775000 ;
      RECT 174.925000  4.725000 175.255000 5.185000 ;
      RECT 175.425000  0.085000 175.675000 0.545000 ;
      RECT 175.425000  1.835000 175.695000 2.635000 ;
      RECT 175.425000  2.805000 175.695000 3.605000 ;
      RECT 175.425000  4.895000 175.675000 5.355000 ;
      RECT 175.845000  0.255000 177.875000 0.425000 ;
      RECT 175.845000  0.425000 176.115000 0.715000 ;
      RECT 175.845000  4.725000 176.115000 5.015000 ;
      RECT 175.845000  5.015000 177.875000 5.185000 ;
      RECT 175.915000  1.665000 176.215000 2.465000 ;
      RECT 175.915000  2.975000 176.215000 3.775000 ;
      RECT 176.285000  0.595000 176.615000 0.885000 ;
      RECT 176.285000  4.555000 176.615000 4.845000 ;
      RECT 176.385000  0.885000 176.615000 1.065000 ;
      RECT 176.385000  1.065000 177.655000 1.365000 ;
      RECT 176.385000  1.365000 176.715000 4.075000 ;
      RECT 176.385000  4.075000 177.655000 4.375000 ;
      RECT 176.385000  4.375000 176.615000 4.555000 ;
      RECT 176.785000  0.425000 176.955000 0.770000 ;
      RECT 176.785000  4.670000 176.955000 5.015000 ;
      RECT 176.885000  1.535000 177.155000 2.465000 ;
      RECT 176.885000  2.975000 177.155000 3.905000 ;
      RECT 177.125000  0.595000 177.455000 1.065000 ;
      RECT 177.125000  4.375000 177.455000 4.845000 ;
      RECT 177.325000  1.365000 177.655000 4.075000 ;
      RECT 177.625000  0.425000 177.875000 0.770000 ;
      RECT 177.625000  4.670000 177.875000 5.015000 ;
      RECT 177.825000  1.065000 179.010000 1.395000 ;
      RECT 177.825000  1.565000 178.125000 2.465000 ;
      RECT 177.825000  2.635000 181.895000 2.805000 ;
      RECT 177.825000  2.975000 178.125000 3.875000 ;
      RECT 177.825000  4.045000 179.010000 4.375000 ;
      RECT 178.370000  1.605000 178.645000 2.635000 ;
      RECT 178.370000  2.805000 178.645000 3.835000 ;
      RECT 178.380000  0.085000 178.670000 0.610000 ;
      RECT 178.380000  4.830000 178.670000 5.355000 ;
      RECT 178.840000  0.280000 179.090000 0.825000 ;
      RECT 178.840000  0.825000 179.010000 1.065000 ;
      RECT 178.840000  1.395000 179.010000 1.605000 ;
      RECT 178.840000  1.605000 179.170000 2.465000 ;
      RECT 178.840000  2.975000 179.170000 3.835000 ;
      RECT 178.840000  3.835000 179.010000 4.045000 ;
      RECT 178.840000  4.375000 179.010000 4.615000 ;
      RECT 178.840000  4.615000 179.090000 5.160000 ;
      RECT 179.180000  0.995000 179.775000 1.325000 ;
      RECT 179.180000  4.115000 179.775000 4.445000 ;
      RECT 179.300000  0.085000 179.590000 0.610000 ;
      RECT 179.300000  4.830000 179.590000 5.355000 ;
      RECT 179.340000  1.605000 179.640000 2.635000 ;
      RECT 179.340000  2.805000 179.640000 3.835000 ;
      RECT 179.945000  0.995000 180.540000 1.325000 ;
      RECT 179.945000  4.115000 180.540000 4.445000 ;
      RECT 180.080000  1.605000 180.380000 2.635000 ;
      RECT 180.080000  2.805000 180.380000 3.835000 ;
      RECT 180.130000  0.085000 180.420000 0.610000 ;
      RECT 180.130000  4.830000 180.420000 5.355000 ;
      RECT 180.550000  1.605000 180.880000 2.465000 ;
      RECT 180.550000  2.975000 180.880000 3.835000 ;
      RECT 180.630000  0.280000 180.880000 0.825000 ;
      RECT 180.630000  4.615000 180.880000 5.160000 ;
      RECT 180.710000  0.825000 180.880000 1.065000 ;
      RECT 180.710000  1.065000 181.895000 1.395000 ;
      RECT 180.710000  1.395000 180.880000 1.605000 ;
      RECT 180.710000  3.835000 180.880000 4.045000 ;
      RECT 180.710000  4.045000 181.895000 4.375000 ;
      RECT 180.710000  4.375000 180.880000 4.615000 ;
      RECT 181.050000  0.085000 181.340000 0.610000 ;
      RECT 181.050000  4.830000 181.340000 5.355000 ;
      RECT 181.075000  1.605000 181.350000 2.635000 ;
      RECT 181.075000  2.805000 181.350000 3.835000 ;
      RECT 181.595000  1.565000 181.895000 2.465000 ;
      RECT 181.595000  2.975000 181.895000 3.875000 ;
      RECT 181.845000  0.255000 183.875000 0.425000 ;
      RECT 181.845000  0.425000 182.095000 0.770000 ;
      RECT 181.845000  4.670000 182.095000 5.015000 ;
      RECT 181.845000  5.015000 183.875000 5.185000 ;
      RECT 182.065000  1.065000 183.335000 1.365000 ;
      RECT 182.065000  1.365000 182.395000 4.075000 ;
      RECT 182.065000  4.075000 183.335000 4.375000 ;
      RECT 182.265000  0.595000 182.595000 1.065000 ;
      RECT 182.265000  4.375000 182.595000 4.845000 ;
      RECT 182.565000  1.535000 182.835000 2.465000 ;
      RECT 182.565000  2.975000 182.835000 3.905000 ;
      RECT 182.765000  0.425000 182.935000 0.770000 ;
      RECT 182.765000  4.670000 182.935000 5.015000 ;
      RECT 183.005000  1.365000 183.335000 4.075000 ;
      RECT 183.105000  0.595000 183.435000 0.885000 ;
      RECT 183.105000  0.885000 183.335000 1.065000 ;
      RECT 183.105000  4.375000 183.335000 4.555000 ;
      RECT 183.105000  4.555000 183.435000 4.845000 ;
      RECT 183.505000  1.495000 185.735000 1.665000 ;
      RECT 183.505000  1.665000 183.805000 2.465000 ;
      RECT 183.505000  2.635000 189.095000 2.805000 ;
      RECT 183.505000  2.975000 183.805000 3.775000 ;
      RECT 183.505000  3.775000 185.735000 3.945000 ;
      RECT 183.605000  0.425000 183.875000 0.715000 ;
      RECT 183.605000  0.715000 185.735000 0.885000 ;
      RECT 183.605000  4.555000 185.735000 4.725000 ;
      RECT 183.605000  4.725000 183.875000 5.015000 ;
      RECT 184.025000  1.835000 184.295000 2.635000 ;
      RECT 184.025000  2.805000 184.295000 3.605000 ;
      RECT 184.045000  0.085000 184.295000 0.545000 ;
      RECT 184.045000  4.895000 184.295000 5.355000 ;
      RECT 184.465000  0.255000 184.795000 0.715000 ;
      RECT 184.465000  1.665000 184.795000 2.465000 ;
      RECT 184.465000  2.975000 184.795000 3.775000 ;
      RECT 184.465000  4.725000 184.795000 5.185000 ;
      RECT 184.515000  1.055000 185.905000 1.325000 ;
      RECT 184.515000  4.115000 185.905000 4.385000 ;
      RECT 184.965000  0.085000 185.235000 0.545000 ;
      RECT 184.965000  1.835000 185.235000 2.635000 ;
      RECT 184.965000  2.805000 185.235000 3.605000 ;
      RECT 184.965000  4.895000 185.235000 5.355000 ;
      RECT 185.405000  0.255000 185.735000 0.715000 ;
      RECT 185.405000  1.665000 185.735000 2.465000 ;
      RECT 185.405000  2.975000 185.735000 3.775000 ;
      RECT 185.405000  4.725000 185.735000 5.185000 ;
      RECT 185.905000  0.085000 186.155000 0.885000 ;
      RECT 185.905000  1.495000 186.175000 2.635000 ;
      RECT 185.905000  2.805000 186.175000 3.945000 ;
      RECT 185.905000  4.555000 186.155000 5.355000 ;
      RECT 186.425000  1.495000 186.695000 2.635000 ;
      RECT 186.425000  2.805000 186.695000 3.945000 ;
      RECT 186.445000  0.085000 186.695000 0.885000 ;
      RECT 186.445000  4.555000 186.695000 5.355000 ;
      RECT 186.695000  1.055000 188.085000 1.325000 ;
      RECT 186.695000  4.115000 188.085000 4.385000 ;
      RECT 186.865000  0.255000 187.195000 0.715000 ;
      RECT 186.865000  0.715000 188.995000 0.885000 ;
      RECT 186.865000  1.495000 189.095000 1.665000 ;
      RECT 186.865000  1.665000 187.195000 2.465000 ;
      RECT 186.865000  2.975000 187.195000 3.775000 ;
      RECT 186.865000  3.775000 189.095000 3.945000 ;
      RECT 186.865000  4.555000 188.995000 4.725000 ;
      RECT 186.865000  4.725000 187.195000 5.185000 ;
      RECT 187.365000  0.085000 187.635000 0.545000 ;
      RECT 187.365000  1.835000 187.635000 2.635000 ;
      RECT 187.365000  2.805000 187.635000 3.605000 ;
      RECT 187.365000  4.895000 187.635000 5.355000 ;
      RECT 187.805000  0.255000 188.135000 0.715000 ;
      RECT 187.805000  1.665000 188.135000 2.465000 ;
      RECT 187.805000  2.975000 188.135000 3.775000 ;
      RECT 187.805000  4.725000 188.135000 5.185000 ;
      RECT 188.305000  0.085000 188.555000 0.545000 ;
      RECT 188.305000  1.835000 188.575000 2.635000 ;
      RECT 188.305000  2.805000 188.575000 3.605000 ;
      RECT 188.305000  4.895000 188.555000 5.355000 ;
      RECT 188.725000  0.255000 190.755000 0.425000 ;
      RECT 188.725000  0.425000 188.995000 0.715000 ;
      RECT 188.725000  4.725000 188.995000 5.015000 ;
      RECT 188.725000  5.015000 190.755000 5.185000 ;
      RECT 188.795000  1.665000 189.095000 2.465000 ;
      RECT 188.795000  2.975000 189.095000 3.775000 ;
      RECT 189.165000  0.595000 189.495000 0.885000 ;
      RECT 189.165000  4.555000 189.495000 4.845000 ;
      RECT 189.265000  0.885000 189.495000 1.065000 ;
      RECT 189.265000  1.065000 190.535000 1.365000 ;
      RECT 189.265000  1.365000 189.595000 4.075000 ;
      RECT 189.265000  4.075000 190.535000 4.375000 ;
      RECT 189.265000  4.375000 189.495000 4.555000 ;
      RECT 189.665000  0.425000 189.835000 0.770000 ;
      RECT 189.665000  4.670000 189.835000 5.015000 ;
      RECT 189.765000  1.535000 190.035000 2.465000 ;
      RECT 189.765000  2.975000 190.035000 3.905000 ;
      RECT 190.005000  0.595000 190.335000 1.065000 ;
      RECT 190.005000  4.375000 190.335000 4.845000 ;
      RECT 190.205000  1.365000 190.535000 4.075000 ;
      RECT 190.505000  0.425000 190.755000 0.770000 ;
      RECT 190.505000  4.670000 190.755000 5.015000 ;
      RECT 190.705000  1.065000 191.890000 1.395000 ;
      RECT 190.705000  1.565000 191.005000 2.465000 ;
      RECT 190.705000  2.635000 194.775000 2.805000 ;
      RECT 190.705000  2.975000 191.005000 3.875000 ;
      RECT 190.705000  4.045000 191.890000 4.375000 ;
      RECT 191.250000  1.605000 191.525000 2.635000 ;
      RECT 191.250000  2.805000 191.525000 3.835000 ;
      RECT 191.260000  0.085000 191.550000 0.610000 ;
      RECT 191.260000  4.830000 191.550000 5.355000 ;
      RECT 191.720000  0.280000 191.970000 0.825000 ;
      RECT 191.720000  0.825000 191.890000 1.065000 ;
      RECT 191.720000  1.395000 191.890000 1.605000 ;
      RECT 191.720000  1.605000 192.050000 2.465000 ;
      RECT 191.720000  2.975000 192.050000 3.835000 ;
      RECT 191.720000  3.835000 191.890000 4.045000 ;
      RECT 191.720000  4.375000 191.890000 4.615000 ;
      RECT 191.720000  4.615000 191.970000 5.160000 ;
      RECT 192.060000  0.995000 192.655000 1.325000 ;
      RECT 192.060000  4.115000 192.655000 4.445000 ;
      RECT 192.180000  0.085000 192.470000 0.610000 ;
      RECT 192.180000  4.830000 192.470000 5.355000 ;
      RECT 192.220000  1.605000 192.520000 2.635000 ;
      RECT 192.220000  2.805000 192.520000 3.835000 ;
      RECT 192.825000  0.995000 193.420000 1.325000 ;
      RECT 192.825000  4.115000 193.420000 4.445000 ;
      RECT 192.960000  1.605000 193.260000 2.635000 ;
      RECT 192.960000  2.805000 193.260000 3.835000 ;
      RECT 193.010000  0.085000 193.300000 0.610000 ;
      RECT 193.010000  4.830000 193.300000 5.355000 ;
      RECT 193.430000  1.605000 193.760000 2.465000 ;
      RECT 193.430000  2.975000 193.760000 3.835000 ;
      RECT 193.510000  0.280000 193.760000 0.825000 ;
      RECT 193.510000  4.615000 193.760000 5.160000 ;
      RECT 193.590000  0.825000 193.760000 1.065000 ;
      RECT 193.590000  1.065000 194.775000 1.395000 ;
      RECT 193.590000  1.395000 193.760000 1.605000 ;
      RECT 193.590000  3.835000 193.760000 4.045000 ;
      RECT 193.590000  4.045000 194.775000 4.375000 ;
      RECT 193.590000  4.375000 193.760000 4.615000 ;
      RECT 193.930000  0.085000 194.220000 0.610000 ;
      RECT 193.930000  4.830000 194.220000 5.355000 ;
      RECT 193.955000  1.605000 194.230000 2.635000 ;
      RECT 193.955000  2.805000 194.230000 3.835000 ;
      RECT 194.475000  1.565000 194.775000 2.465000 ;
      RECT 194.475000  2.975000 194.775000 3.875000 ;
      RECT 194.725000  0.255000 196.755000 0.425000 ;
      RECT 194.725000  0.425000 194.975000 0.770000 ;
      RECT 194.725000  4.670000 194.975000 5.015000 ;
      RECT 194.725000  5.015000 196.755000 5.185000 ;
      RECT 194.945000  1.065000 196.215000 1.365000 ;
      RECT 194.945000  1.365000 195.275000 4.075000 ;
      RECT 194.945000  4.075000 196.215000 4.375000 ;
      RECT 195.145000  0.595000 195.475000 1.065000 ;
      RECT 195.145000  4.375000 195.475000 4.845000 ;
      RECT 195.445000  1.535000 195.715000 2.465000 ;
      RECT 195.445000  2.975000 195.715000 3.905000 ;
      RECT 195.645000  0.425000 195.815000 0.770000 ;
      RECT 195.645000  4.670000 195.815000 5.015000 ;
      RECT 195.885000  1.365000 196.215000 4.075000 ;
      RECT 195.985000  0.595000 196.315000 0.885000 ;
      RECT 195.985000  0.885000 196.215000 1.065000 ;
      RECT 195.985000  4.375000 196.215000 4.555000 ;
      RECT 195.985000  4.555000 196.315000 4.845000 ;
      RECT 196.385000  1.495000 198.615000 1.665000 ;
      RECT 196.385000  1.665000 196.685000 2.465000 ;
      RECT 196.385000  2.635000 202.435000 2.805000 ;
      RECT 196.385000  2.975000 196.685000 3.775000 ;
      RECT 196.385000  3.775000 198.615000 3.945000 ;
      RECT 196.485000  0.425000 196.755000 0.715000 ;
      RECT 196.485000  0.715000 198.615000 0.885000 ;
      RECT 196.485000  4.555000 198.615000 4.725000 ;
      RECT 196.485000  4.725000 196.755000 5.015000 ;
      RECT 196.905000  1.835000 197.175000 2.635000 ;
      RECT 196.905000  2.805000 197.175000 3.605000 ;
      RECT 196.925000  0.085000 197.175000 0.545000 ;
      RECT 196.925000  4.895000 197.175000 5.355000 ;
      RECT 197.345000  0.255000 197.675000 0.715000 ;
      RECT 197.345000  1.665000 197.675000 2.465000 ;
      RECT 197.345000  2.975000 197.675000 3.775000 ;
      RECT 197.345000  4.725000 197.675000 5.185000 ;
      RECT 197.395000  1.055000 198.785000 1.325000 ;
      RECT 197.395000  4.115000 198.785000 4.385000 ;
      RECT 197.845000  0.085000 198.115000 0.545000 ;
      RECT 197.845000  1.835000 198.115000 2.635000 ;
      RECT 197.845000  2.805000 198.115000 3.605000 ;
      RECT 197.845000  4.895000 198.115000 5.355000 ;
      RECT 198.285000  0.255000 198.615000 0.715000 ;
      RECT 198.285000  1.665000 198.615000 2.465000 ;
      RECT 198.285000  2.975000 198.615000 3.775000 ;
      RECT 198.285000  4.725000 198.615000 5.185000 ;
      RECT 198.785000  0.085000 199.035000 0.885000 ;
      RECT 198.785000  1.495000 199.055000 2.635000 ;
      RECT 198.785000  2.805000 199.055000 3.945000 ;
      RECT 198.785000  4.555000 199.035000 5.355000 ;
      RECT 199.265000  0.265000 199.555000 0.810000 ;
      RECT 199.265000  1.470000 199.555000 2.455000 ;
      RECT 199.265000  2.985000 199.555000 3.970000 ;
      RECT 199.265000  4.630000 199.555000 5.175000 ;
      RECT 199.765000  1.495000 200.035000 2.635000 ;
      RECT 199.765000  2.805000 200.035000 3.945000 ;
      RECT 199.785000  0.085000 200.035000 0.885000 ;
      RECT 199.785000  4.555000 200.035000 5.355000 ;
      RECT 200.035000  1.055000 201.425000 1.325000 ;
      RECT 200.035000  4.115000 201.425000 4.385000 ;
      RECT 200.205000  0.255000 200.535000 0.715000 ;
      RECT 200.205000  0.715000 202.335000 0.885000 ;
      RECT 200.205000  1.495000 202.435000 1.665000 ;
      RECT 200.205000  1.665000 200.535000 2.465000 ;
      RECT 200.205000  2.975000 200.535000 3.775000 ;
      RECT 200.205000  3.775000 202.435000 3.945000 ;
      RECT 200.205000  4.555000 202.335000 4.725000 ;
      RECT 200.205000  4.725000 200.535000 5.185000 ;
      RECT 200.705000  0.085000 200.975000 0.545000 ;
      RECT 200.705000  1.835000 200.975000 2.635000 ;
      RECT 200.705000  2.805000 200.975000 3.605000 ;
      RECT 200.705000  4.895000 200.975000 5.355000 ;
      RECT 201.145000  0.255000 201.475000 0.715000 ;
      RECT 201.145000  1.665000 201.475000 2.465000 ;
      RECT 201.145000  2.975000 201.475000 3.775000 ;
      RECT 201.145000  4.725000 201.475000 5.185000 ;
      RECT 201.645000  0.085000 201.895000 0.545000 ;
      RECT 201.645000  1.835000 201.915000 2.635000 ;
      RECT 201.645000  2.805000 201.915000 3.605000 ;
      RECT 201.645000  4.895000 201.895000 5.355000 ;
      RECT 202.065000  0.255000 204.095000 0.425000 ;
      RECT 202.065000  0.425000 202.335000 0.715000 ;
      RECT 202.065000  4.725000 202.335000 5.015000 ;
      RECT 202.065000  5.015000 204.095000 5.185000 ;
      RECT 202.135000  1.665000 202.435000 2.465000 ;
      RECT 202.135000  2.975000 202.435000 3.775000 ;
      RECT 202.505000  0.595000 202.835000 0.885000 ;
      RECT 202.505000  4.555000 202.835000 4.845000 ;
      RECT 202.605000  0.885000 202.835000 1.065000 ;
      RECT 202.605000  1.065000 203.875000 1.365000 ;
      RECT 202.605000  1.365000 202.935000 4.075000 ;
      RECT 202.605000  4.075000 203.875000 4.375000 ;
      RECT 202.605000  4.375000 202.835000 4.555000 ;
      RECT 203.005000  0.425000 203.175000 0.770000 ;
      RECT 203.005000  4.670000 203.175000 5.015000 ;
      RECT 203.105000  1.535000 203.375000 2.465000 ;
      RECT 203.105000  2.975000 203.375000 3.905000 ;
      RECT 203.345000  0.595000 203.675000 1.065000 ;
      RECT 203.345000  4.375000 203.675000 4.845000 ;
      RECT 203.545000  1.365000 203.875000 4.075000 ;
      RECT 203.845000  0.425000 204.095000 0.770000 ;
      RECT 203.845000  4.670000 204.095000 5.015000 ;
      RECT 204.045000  1.065000 205.230000 1.395000 ;
      RECT 204.045000  1.565000 204.345000 2.465000 ;
      RECT 204.045000  2.635000 208.115000 2.805000 ;
      RECT 204.045000  2.975000 204.345000 3.875000 ;
      RECT 204.045000  4.045000 205.230000 4.375000 ;
      RECT 204.590000  1.605000 204.865000 2.635000 ;
      RECT 204.590000  2.805000 204.865000 3.835000 ;
      RECT 204.600000  0.085000 204.890000 0.610000 ;
      RECT 204.600000  4.830000 204.890000 5.355000 ;
      RECT 205.060000  0.280000 205.310000 0.825000 ;
      RECT 205.060000  0.825000 205.230000 1.065000 ;
      RECT 205.060000  1.395000 205.230000 1.605000 ;
      RECT 205.060000  1.605000 205.390000 2.465000 ;
      RECT 205.060000  2.975000 205.390000 3.835000 ;
      RECT 205.060000  3.835000 205.230000 4.045000 ;
      RECT 205.060000  4.375000 205.230000 4.615000 ;
      RECT 205.060000  4.615000 205.310000 5.160000 ;
      RECT 205.400000  0.995000 205.995000 1.325000 ;
      RECT 205.400000  4.115000 205.995000 4.445000 ;
      RECT 205.520000  0.085000 205.810000 0.610000 ;
      RECT 205.520000  4.830000 205.810000 5.355000 ;
      RECT 205.560000  1.605000 205.860000 2.635000 ;
      RECT 205.560000  2.805000 205.860000 3.835000 ;
      RECT 206.165000  0.995000 206.760000 1.325000 ;
      RECT 206.165000  4.115000 206.760000 4.445000 ;
      RECT 206.300000  1.605000 206.600000 2.635000 ;
      RECT 206.300000  2.805000 206.600000 3.835000 ;
      RECT 206.350000  0.085000 206.640000 0.610000 ;
      RECT 206.350000  4.830000 206.640000 5.355000 ;
      RECT 206.770000  1.605000 207.100000 2.465000 ;
      RECT 206.770000  2.975000 207.100000 3.835000 ;
      RECT 206.850000  0.280000 207.100000 0.825000 ;
      RECT 206.850000  4.615000 207.100000 5.160000 ;
      RECT 206.930000  0.825000 207.100000 1.065000 ;
      RECT 206.930000  1.065000 208.115000 1.395000 ;
      RECT 206.930000  1.395000 207.100000 1.605000 ;
      RECT 206.930000  3.835000 207.100000 4.045000 ;
      RECT 206.930000  4.045000 208.115000 4.375000 ;
      RECT 206.930000  4.375000 207.100000 4.615000 ;
      RECT 207.270000  0.085000 207.560000 0.610000 ;
      RECT 207.270000  4.830000 207.560000 5.355000 ;
      RECT 207.295000  1.605000 207.570000 2.635000 ;
      RECT 207.295000  2.805000 207.570000 3.835000 ;
      RECT 207.815000  1.565000 208.115000 2.465000 ;
      RECT 207.815000  2.975000 208.115000 3.875000 ;
      RECT 208.065000  0.255000 210.095000 0.425000 ;
      RECT 208.065000  0.425000 208.315000 0.770000 ;
      RECT 208.065000  4.670000 208.315000 5.015000 ;
      RECT 208.065000  5.015000 210.095000 5.185000 ;
      RECT 208.285000  1.065000 209.555000 1.365000 ;
      RECT 208.285000  1.365000 208.615000 4.075000 ;
      RECT 208.285000  4.075000 209.555000 4.375000 ;
      RECT 208.485000  0.595000 208.815000 1.065000 ;
      RECT 208.485000  4.375000 208.815000 4.845000 ;
      RECT 208.785000  1.535000 209.055000 2.465000 ;
      RECT 208.785000  2.975000 209.055000 3.905000 ;
      RECT 208.985000  0.425000 209.155000 0.770000 ;
      RECT 208.985000  4.670000 209.155000 5.015000 ;
      RECT 209.225000  1.365000 209.555000 4.075000 ;
      RECT 209.325000  0.595000 209.655000 0.885000 ;
      RECT 209.325000  0.885000 209.555000 1.065000 ;
      RECT 209.325000  4.375000 209.555000 4.555000 ;
      RECT 209.325000  4.555000 209.655000 4.845000 ;
      RECT 209.725000  1.495000 211.955000 1.665000 ;
      RECT 209.725000  1.665000 210.025000 2.465000 ;
      RECT 209.725000  2.635000 215.315000 2.805000 ;
      RECT 209.725000  2.975000 210.025000 3.775000 ;
      RECT 209.725000  3.775000 211.955000 3.945000 ;
      RECT 209.825000  0.425000 210.095000 0.715000 ;
      RECT 209.825000  0.715000 211.955000 0.885000 ;
      RECT 209.825000  4.555000 211.955000 4.725000 ;
      RECT 209.825000  4.725000 210.095000 5.015000 ;
      RECT 210.245000  1.835000 210.515000 2.635000 ;
      RECT 210.245000  2.805000 210.515000 3.605000 ;
      RECT 210.265000  0.085000 210.515000 0.545000 ;
      RECT 210.265000  4.895000 210.515000 5.355000 ;
      RECT 210.685000  0.255000 211.015000 0.715000 ;
      RECT 210.685000  1.665000 211.015000 2.465000 ;
      RECT 210.685000  2.975000 211.015000 3.775000 ;
      RECT 210.685000  4.725000 211.015000 5.185000 ;
      RECT 210.735000  1.055000 212.125000 1.325000 ;
      RECT 210.735000  4.115000 212.125000 4.385000 ;
      RECT 211.185000  0.085000 211.455000 0.545000 ;
      RECT 211.185000  1.835000 211.455000 2.635000 ;
      RECT 211.185000  2.805000 211.455000 3.605000 ;
      RECT 211.185000  4.895000 211.455000 5.355000 ;
      RECT 211.625000  0.255000 211.955000 0.715000 ;
      RECT 211.625000  1.665000 211.955000 2.465000 ;
      RECT 211.625000  2.975000 211.955000 3.775000 ;
      RECT 211.625000  4.725000 211.955000 5.185000 ;
      RECT 212.125000  0.085000 212.375000 0.885000 ;
      RECT 212.125000  1.495000 212.395000 2.635000 ;
      RECT 212.125000  2.805000 212.395000 3.945000 ;
      RECT 212.125000  4.555000 212.375000 5.355000 ;
      RECT 212.645000  1.495000 212.915000 2.635000 ;
      RECT 212.645000  2.805000 212.915000 3.945000 ;
      RECT 212.665000  0.085000 212.915000 0.885000 ;
      RECT 212.665000  4.555000 212.915000 5.355000 ;
      RECT 212.915000  1.055000 214.305000 1.325000 ;
      RECT 212.915000  4.115000 214.305000 4.385000 ;
      RECT 213.085000  0.255000 213.415000 0.715000 ;
      RECT 213.085000  0.715000 215.215000 0.885000 ;
      RECT 213.085000  1.495000 215.315000 1.665000 ;
      RECT 213.085000  1.665000 213.415000 2.465000 ;
      RECT 213.085000  2.975000 213.415000 3.775000 ;
      RECT 213.085000  3.775000 215.315000 3.945000 ;
      RECT 213.085000  4.555000 215.215000 4.725000 ;
      RECT 213.085000  4.725000 213.415000 5.185000 ;
      RECT 213.585000  0.085000 213.855000 0.545000 ;
      RECT 213.585000  1.835000 213.855000 2.635000 ;
      RECT 213.585000  2.805000 213.855000 3.605000 ;
      RECT 213.585000  4.895000 213.855000 5.355000 ;
      RECT 214.025000  0.255000 214.355000 0.715000 ;
      RECT 214.025000  1.665000 214.355000 2.465000 ;
      RECT 214.025000  2.975000 214.355000 3.775000 ;
      RECT 214.025000  4.725000 214.355000 5.185000 ;
      RECT 214.525000  0.085000 214.775000 0.545000 ;
      RECT 214.525000  1.835000 214.795000 2.635000 ;
      RECT 214.525000  2.805000 214.795000 3.605000 ;
      RECT 214.525000  4.895000 214.775000 5.355000 ;
      RECT 214.945000  0.255000 216.975000 0.425000 ;
      RECT 214.945000  0.425000 215.215000 0.715000 ;
      RECT 214.945000  4.725000 215.215000 5.015000 ;
      RECT 214.945000  5.015000 216.975000 5.185000 ;
      RECT 215.015000  1.665000 215.315000 2.465000 ;
      RECT 215.015000  2.975000 215.315000 3.775000 ;
      RECT 215.385000  0.595000 215.715000 0.885000 ;
      RECT 215.385000  4.555000 215.715000 4.845000 ;
      RECT 215.485000  0.885000 215.715000 1.065000 ;
      RECT 215.485000  1.065000 216.755000 1.365000 ;
      RECT 215.485000  1.365000 215.815000 4.075000 ;
      RECT 215.485000  4.075000 216.755000 4.375000 ;
      RECT 215.485000  4.375000 215.715000 4.555000 ;
      RECT 215.885000  0.425000 216.055000 0.770000 ;
      RECT 215.885000  4.670000 216.055000 5.015000 ;
      RECT 215.985000  1.535000 216.255000 2.465000 ;
      RECT 215.985000  2.975000 216.255000 3.905000 ;
      RECT 216.225000  0.595000 216.555000 1.065000 ;
      RECT 216.225000  4.375000 216.555000 4.845000 ;
      RECT 216.425000  1.365000 216.755000 4.075000 ;
      RECT 216.725000  0.425000 216.975000 0.770000 ;
      RECT 216.725000  4.670000 216.975000 5.015000 ;
      RECT 216.925000  1.065000 218.110000 1.395000 ;
      RECT 216.925000  1.565000 217.225000 2.465000 ;
      RECT 216.925000  2.635000 220.995000 2.805000 ;
      RECT 216.925000  2.975000 217.225000 3.875000 ;
      RECT 216.925000  4.045000 218.110000 4.375000 ;
      RECT 217.470000  1.605000 217.745000 2.635000 ;
      RECT 217.470000  2.805000 217.745000 3.835000 ;
      RECT 217.480000  0.085000 217.770000 0.610000 ;
      RECT 217.480000  4.830000 217.770000 5.355000 ;
      RECT 217.940000  0.280000 218.190000 0.825000 ;
      RECT 217.940000  0.825000 218.110000 1.065000 ;
      RECT 217.940000  1.395000 218.110000 1.605000 ;
      RECT 217.940000  1.605000 218.270000 2.465000 ;
      RECT 217.940000  2.975000 218.270000 3.835000 ;
      RECT 217.940000  3.835000 218.110000 4.045000 ;
      RECT 217.940000  4.375000 218.110000 4.615000 ;
      RECT 217.940000  4.615000 218.190000 5.160000 ;
      RECT 218.280000  0.995000 218.875000 1.325000 ;
      RECT 218.280000  4.115000 218.875000 4.445000 ;
      RECT 218.400000  0.085000 218.690000 0.610000 ;
      RECT 218.400000  4.830000 218.690000 5.355000 ;
      RECT 218.440000  1.605000 218.740000 2.635000 ;
      RECT 218.440000  2.805000 218.740000 3.835000 ;
      RECT 219.045000  0.995000 219.640000 1.325000 ;
      RECT 219.045000  4.115000 219.640000 4.445000 ;
      RECT 219.180000  1.605000 219.480000 2.635000 ;
      RECT 219.180000  2.805000 219.480000 3.835000 ;
      RECT 219.230000  0.085000 219.520000 0.610000 ;
      RECT 219.230000  4.830000 219.520000 5.355000 ;
      RECT 219.650000  1.605000 219.980000 2.465000 ;
      RECT 219.650000  2.975000 219.980000 3.835000 ;
      RECT 219.730000  0.280000 219.980000 0.825000 ;
      RECT 219.730000  4.615000 219.980000 5.160000 ;
      RECT 219.810000  0.825000 219.980000 1.065000 ;
      RECT 219.810000  1.065000 220.995000 1.395000 ;
      RECT 219.810000  1.395000 219.980000 1.605000 ;
      RECT 219.810000  3.835000 219.980000 4.045000 ;
      RECT 219.810000  4.045000 220.995000 4.375000 ;
      RECT 219.810000  4.375000 219.980000 4.615000 ;
      RECT 220.150000  0.085000 220.440000 0.610000 ;
      RECT 220.150000  4.830000 220.440000 5.355000 ;
      RECT 220.175000  1.605000 220.450000 2.635000 ;
      RECT 220.175000  2.805000 220.450000 3.835000 ;
      RECT 220.695000  1.565000 220.995000 2.465000 ;
      RECT 220.695000  2.975000 220.995000 3.875000 ;
      RECT 220.945000  0.255000 222.975000 0.425000 ;
      RECT 220.945000  0.425000 221.195000 0.770000 ;
      RECT 220.945000  4.670000 221.195000 5.015000 ;
      RECT 220.945000  5.015000 222.975000 5.185000 ;
      RECT 221.165000  1.065000 222.435000 1.365000 ;
      RECT 221.165000  1.365000 221.495000 4.075000 ;
      RECT 221.165000  4.075000 222.435000 4.375000 ;
      RECT 221.365000  0.595000 221.695000 1.065000 ;
      RECT 221.365000  4.375000 221.695000 4.845000 ;
      RECT 221.665000  1.535000 221.935000 2.465000 ;
      RECT 221.665000  2.975000 221.935000 3.905000 ;
      RECT 221.865000  0.425000 222.035000 0.770000 ;
      RECT 221.865000  4.670000 222.035000 5.015000 ;
      RECT 222.105000  1.365000 222.435000 4.075000 ;
      RECT 222.205000  0.595000 222.535000 0.885000 ;
      RECT 222.205000  0.885000 222.435000 1.065000 ;
      RECT 222.205000  4.375000 222.435000 4.555000 ;
      RECT 222.205000  4.555000 222.535000 4.845000 ;
      RECT 222.605000  1.495000 224.835000 1.665000 ;
      RECT 222.605000  1.665000 222.905000 2.465000 ;
      RECT 222.605000  2.635000 225.400000 2.805000 ;
      RECT 222.605000  2.975000 222.905000 3.775000 ;
      RECT 222.605000  3.775000 224.835000 3.945000 ;
      RECT 222.705000  0.425000 222.975000 0.715000 ;
      RECT 222.705000  0.715000 224.835000 0.885000 ;
      RECT 222.705000  4.555000 224.835000 4.725000 ;
      RECT 222.705000  4.725000 222.975000 5.015000 ;
      RECT 223.125000  1.835000 223.395000 2.635000 ;
      RECT 223.125000  2.805000 223.395000 3.605000 ;
      RECT 223.145000  0.085000 223.395000 0.545000 ;
      RECT 223.145000  4.895000 223.395000 5.355000 ;
      RECT 223.565000  0.255000 223.895000 0.715000 ;
      RECT 223.565000  1.665000 223.895000 2.465000 ;
      RECT 223.565000  2.975000 223.895000 3.775000 ;
      RECT 223.565000  4.725000 223.895000 5.185000 ;
      RECT 223.615000  1.055000 225.005000 1.325000 ;
      RECT 223.615000  4.115000 225.005000 4.385000 ;
      RECT 224.065000  0.085000 224.335000 0.545000 ;
      RECT 224.065000  1.835000 224.335000 2.635000 ;
      RECT 224.065000  2.805000 224.335000 3.605000 ;
      RECT 224.065000  4.895000 224.335000 5.355000 ;
      RECT 224.505000  0.255000 224.835000 0.715000 ;
      RECT 224.505000  1.665000 224.835000 2.465000 ;
      RECT 224.505000  2.975000 224.835000 3.775000 ;
      RECT 224.505000  4.725000 224.835000 5.185000 ;
      RECT 225.005000  0.085000 225.255000 0.885000 ;
      RECT 225.005000  1.495000 225.275000 2.635000 ;
      RECT 225.005000  2.805000 225.275000 3.945000 ;
      RECT 225.005000  4.555000 225.255000 5.355000 ;
    LAYER mcon ;
      RECT   0.145000 -0.085000   0.315000 0.085000 ;
      RECT   0.145000  2.635000   0.315000 2.805000 ;
      RECT   0.605000 -0.085000   0.775000 0.085000 ;
      RECT   0.605000  2.635000   0.775000 2.805000 ;
      RECT   1.065000 -0.085000   1.235000 0.085000 ;
      RECT   1.065000  2.635000   1.235000 2.805000 ;
      RECT   1.525000 -0.085000   1.695000 0.085000 ;
      RECT   1.525000  2.635000   1.695000 2.805000 ;
      RECT   1.985000 -0.085000   2.155000 0.085000 ;
      RECT   1.985000  2.635000   2.155000 2.805000 ;
      RECT   2.445000 -0.085000   2.615000 0.085000 ;
      RECT   2.445000  2.635000   2.615000 2.805000 ;
      RECT   2.905000 -0.085000   3.075000 0.085000 ;
      RECT   2.905000  2.635000   3.075000 2.805000 ;
      RECT   3.365000 -0.085000   3.535000 0.085000 ;
      RECT   3.365000  2.635000   3.535000 2.805000 ;
      RECT   3.825000 -0.085000   3.995000 0.085000 ;
      RECT   3.825000  2.635000   3.995000 2.805000 ;
      RECT   4.285000 -0.085000   4.455000 0.085000 ;
      RECT   4.285000  2.635000   4.455000 2.805000 ;
      RECT   4.745000 -0.085000   4.915000 0.085000 ;
      RECT   4.745000  2.635000   4.915000 2.805000 ;
      RECT   5.205000 -0.085000   5.375000 0.085000 ;
      RECT   5.205000  2.635000   5.375000 2.805000 ;
      RECT   5.665000 -0.085000   5.835000 0.085000 ;
      RECT   5.665000  2.635000   5.835000 2.805000 ;
      RECT   6.125000 -0.085000   6.295000 0.085000 ;
      RECT   6.125000  2.635000   6.295000 2.805000 ;
      RECT   6.585000 -0.085000   6.755000 0.085000 ;
      RECT   6.585000  2.635000   6.755000 2.805000 ;
      RECT   7.045000 -0.085000   7.215000 0.085000 ;
      RECT   7.045000  2.635000   7.215000 2.805000 ;
      RECT   7.505000 -0.085000   7.675000 0.085000 ;
      RECT   7.505000  2.635000   7.675000 2.805000 ;
      RECT   7.965000 -0.085000   8.135000 0.085000 ;
      RECT   7.965000  2.635000   8.135000 2.805000 ;
      RECT   8.425000 -0.085000   8.595000 0.085000 ;
      RECT   8.425000  2.635000   8.595000 2.805000 ;
      RECT   8.885000 -0.085000   9.055000 0.085000 ;
      RECT   8.885000  2.635000   9.055000 2.805000 ;
      RECT   9.345000 -0.085000   9.515000 0.085000 ;
      RECT   9.345000  2.635000   9.515000 2.805000 ;
      RECT   9.805000 -0.085000   9.975000 0.085000 ;
      RECT   9.805000  2.635000   9.975000 2.805000 ;
      RECT  10.265000 -0.085000  10.435000 0.085000 ;
      RECT  10.265000  2.635000  10.435000 2.805000 ;
      RECT  10.725000 -0.085000  10.895000 0.085000 ;
      RECT  10.725000  2.635000  10.895000 2.805000 ;
      RECT  11.185000 -0.085000  11.355000 0.085000 ;
      RECT  11.185000  2.635000  11.355000 2.805000 ;
      RECT  11.645000 -0.085000  11.815000 0.085000 ;
      RECT  11.645000  2.635000  11.815000 2.805000 ;
      RECT  12.105000 -0.085000  12.275000 0.085000 ;
      RECT  12.105000  2.635000  12.275000 2.805000 ;
      RECT  12.565000 -0.085000  12.735000 0.085000 ;
      RECT  12.565000  2.635000  12.735000 2.805000 ;
      RECT  13.025000 -0.085000  13.195000 0.085000 ;
      RECT  13.025000  2.635000  13.195000 2.805000 ;
      RECT  13.485000 -0.085000  13.655000 0.085000 ;
      RECT  13.485000  2.635000  13.655000 2.805000 ;
      RECT  13.945000 -0.085000  14.115000 0.085000 ;
      RECT  13.945000  2.635000  14.115000 2.805000 ;
      RECT  14.405000 -0.085000  14.575000 0.085000 ;
      RECT  14.405000  2.635000  14.575000 2.805000 ;
      RECT  14.865000 -0.085000  15.035000 0.085000 ;
      RECT  14.865000  2.635000  15.035000 2.805000 ;
      RECT  15.325000 -0.085000  15.495000 0.085000 ;
      RECT  15.325000  2.635000  15.495000 2.805000 ;
      RECT  15.785000 -0.085000  15.955000 0.085000 ;
      RECT  15.785000  2.635000  15.955000 2.805000 ;
      RECT  16.245000 -0.085000  16.415000 0.085000 ;
      RECT  16.245000  2.635000  16.415000 2.805000 ;
      RECT  16.705000 -0.085000  16.875000 0.085000 ;
      RECT  16.705000  1.785000  16.875000 1.955000 ;
      RECT  16.705000  2.635000  16.875000 2.805000 ;
      RECT  17.165000 -0.085000  17.335000 0.085000 ;
      RECT  17.165000  2.635000  17.335000 2.805000 ;
      RECT  17.625000 -0.085000  17.795000 0.085000 ;
      RECT  17.625000  2.635000  17.795000 2.805000 ;
      RECT  18.085000 -0.085000  18.255000 0.085000 ;
      RECT  18.085000  2.635000  18.255000 2.805000 ;
      RECT  18.545000 -0.085000  18.715000 0.085000 ;
      RECT  18.545000  2.635000  18.715000 2.805000 ;
      RECT  19.005000 -0.085000  19.175000 0.085000 ;
      RECT  19.005000  1.785000  19.175000 1.955000 ;
      RECT  19.005000  2.635000  19.175000 2.805000 ;
      RECT  19.465000 -0.085000  19.635000 0.085000 ;
      RECT  19.465000  2.635000  19.635000 2.805000 ;
      RECT  19.925000 -0.085000  20.095000 0.085000 ;
      RECT  19.925000  2.635000  20.095000 2.805000 ;
      RECT  20.385000 -0.085000  20.555000 0.085000 ;
      RECT  20.385000  2.635000  20.555000 2.805000 ;
      RECT  20.845000 -0.085000  21.015000 0.085000 ;
      RECT  20.845000  1.785000  21.015000 1.955000 ;
      RECT  20.845000  2.635000  21.015000 2.805000 ;
      RECT  21.305000 -0.085000  21.475000 0.085000 ;
      RECT  21.305000  2.635000  21.475000 2.805000 ;
      RECT  21.765000 -0.085000  21.935000 0.085000 ;
      RECT  21.765000  2.635000  21.935000 2.805000 ;
      RECT  22.225000 -0.085000  22.395000 0.085000 ;
      RECT  22.225000  2.635000  22.395000 2.805000 ;
      RECT  22.685000 -0.085000  22.855000 0.085000 ;
      RECT  22.685000  2.635000  22.855000 2.805000 ;
      RECT  23.145000 -0.085000  23.315000 0.085000 ;
      RECT  23.145000  1.785000  23.315000 1.955000 ;
      RECT  23.145000  2.635000  23.315000 2.805000 ;
      RECT  23.605000 -0.085000  23.775000 0.085000 ;
      RECT  23.605000  2.635000  23.775000 2.805000 ;
      RECT  24.065000 -0.085000  24.235000 0.085000 ;
      RECT  24.065000  2.635000  24.235000 2.805000 ;
      RECT  24.525000 -0.085000  24.695000 0.085000 ;
      RECT  24.525000  2.635000  24.695000 2.805000 ;
      RECT  24.985000 -0.085000  25.155000 0.085000 ;
      RECT  24.985000  2.635000  25.155000 2.805000 ;
      RECT  25.445000 -0.085000  25.615000 0.085000 ;
      RECT  25.445000  2.635000  25.615000 2.805000 ;
      RECT  25.905000 -0.085000  26.075000 0.085000 ;
      RECT  25.905000  1.785000  26.075000 1.955000 ;
      RECT  25.905000  2.635000  26.075000 2.805000 ;
      RECT  26.365000 -0.085000  26.535000 0.085000 ;
      RECT  26.365000  2.635000  26.535000 2.805000 ;
      RECT  26.825000 -0.085000  26.995000 0.085000 ;
      RECT  26.825000  2.635000  26.995000 2.805000 ;
      RECT  27.285000 -0.085000  27.455000 0.085000 ;
      RECT  27.285000  2.635000  27.455000 2.805000 ;
      RECT  27.745000 -0.085000  27.915000 0.085000 ;
      RECT  27.745000  2.635000  27.915000 2.805000 ;
      RECT  28.205000 -0.085000  28.375000 0.085000 ;
      RECT  28.205000  2.635000  28.375000 2.805000 ;
      RECT  28.665000 -0.085000  28.835000 0.085000 ;
      RECT  28.665000  2.635000  28.835000 2.805000 ;
      RECT  29.125000 -0.085000  29.295000 0.085000 ;
      RECT  29.125000  1.785000  29.295000 1.955000 ;
      RECT  29.125000  2.635000  29.295000 2.805000 ;
      RECT  29.585000 -0.085000  29.755000 0.085000 ;
      RECT  29.585000  2.635000  29.755000 2.805000 ;
      RECT  30.045000 -0.085000  30.215000 0.085000 ;
      RECT  30.045000  2.635000  30.215000 2.805000 ;
      RECT  30.505000 -0.085000  30.675000 0.085000 ;
      RECT  30.505000  2.635000  30.675000 2.805000 ;
      RECT  30.965000 -0.085000  31.135000 0.085000 ;
      RECT  30.965000  2.635000  31.135000 2.805000 ;
      RECT  31.425000 -0.085000  31.595000 0.085000 ;
      RECT  31.425000  2.635000  31.595000 2.805000 ;
      RECT  31.885000 -0.085000  32.055000 0.085000 ;
      RECT  31.885000  2.635000  32.055000 2.805000 ;
      RECT  32.345000 -0.085000  32.515000 0.085000 ;
      RECT  32.345000  1.785000  32.515000 1.955000 ;
      RECT  32.345000  2.635000  32.515000 2.805000 ;
      RECT  32.805000 -0.085000  32.975000 0.085000 ;
      RECT  32.805000  2.635000  32.975000 2.805000 ;
      RECT  33.265000 -0.085000  33.435000 0.085000 ;
      RECT  33.265000  2.635000  33.435000 2.805000 ;
      RECT  33.725000 -0.085000  33.895000 0.085000 ;
      RECT  33.725000  2.635000  33.895000 2.805000 ;
      RECT  34.185000 -0.085000  34.355000 0.085000 ;
      RECT  34.185000  2.635000  34.355000 2.805000 ;
      RECT  34.645000 -0.085000  34.815000 0.085000 ;
      RECT  34.645000  2.635000  34.815000 2.805000 ;
      RECT  35.105000 -0.085000  35.275000 0.085000 ;
      RECT  35.105000  2.635000  35.275000 2.805000 ;
      RECT  35.565000 -0.085000  35.735000 0.085000 ;
      RECT  35.565000  1.785000  35.735000 1.955000 ;
      RECT  35.565000  2.635000  35.735000 2.805000 ;
      RECT  36.025000 -0.085000  36.195000 0.085000 ;
      RECT  36.025000  2.635000  36.195000 2.805000 ;
      RECT  36.485000 -0.085000  36.655000 0.085000 ;
      RECT  36.485000  2.635000  36.655000 2.805000 ;
      RECT  36.945000 -0.085000  37.115000 0.085000 ;
      RECT  36.945000  2.635000  37.115000 2.805000 ;
      RECT  37.405000 -0.085000  37.575000 0.085000 ;
      RECT  37.405000  2.635000  37.575000 2.805000 ;
      RECT  37.865000 -0.085000  38.035000 0.085000 ;
      RECT  37.865000  2.635000  38.035000 2.805000 ;
      RECT  38.325000 -0.085000  38.495000 0.085000 ;
      RECT  38.325000  2.635000  38.495000 2.805000 ;
      RECT  38.785000 -0.085000  38.955000 0.085000 ;
      RECT  38.785000  2.635000  38.955000 2.805000 ;
      RECT  39.245000 -0.085000  39.415000 0.085000 ;
      RECT  39.245000  2.635000  39.415000 2.805000 ;
      RECT  39.705000 -0.085000  39.875000 0.085000 ;
      RECT  39.705000  2.635000  39.875000 2.805000 ;
      RECT  40.165000 -0.085000  40.335000 0.085000 ;
      RECT  40.165000  2.635000  40.335000 2.805000 ;
      RECT  40.305000  1.785000  40.475000 1.955000 ;
      RECT  40.625000 -0.085000  40.795000 0.085000 ;
      RECT  40.625000  2.635000  40.795000 2.805000 ;
      RECT  41.085000 -0.085000  41.255000 0.085000 ;
      RECT  41.085000  2.635000  41.255000 2.805000 ;
      RECT  41.245000  1.785000  41.415000 1.955000 ;
      RECT  41.545000 -0.085000  41.715000 0.085000 ;
      RECT  41.545000  2.635000  41.715000 2.805000 ;
      RECT  42.005000 -0.085000  42.175000 0.085000 ;
      RECT  42.005000  2.635000  42.175000 2.805000 ;
      RECT  42.465000 -0.085000  42.635000 0.085000 ;
      RECT  42.465000  2.635000  42.635000 2.805000 ;
      RECT  42.925000 -0.085000  43.095000 0.085000 ;
      RECT  42.925000  2.635000  43.095000 2.805000 ;
      RECT  43.385000 -0.085000  43.555000 0.085000 ;
      RECT  43.385000  2.635000  43.555000 2.805000 ;
      RECT  43.845000 -0.085000  44.015000 0.085000 ;
      RECT  43.845000  2.635000  44.015000 2.805000 ;
      RECT  44.305000 -0.085000  44.475000 0.085000 ;
      RECT  44.305000  2.635000  44.475000 2.805000 ;
      RECT  44.765000 -0.085000  44.935000 0.085000 ;
      RECT  44.765000  2.635000  44.935000 2.805000 ;
      RECT  45.225000 -0.085000  45.395000 0.085000 ;
      RECT  45.225000  2.635000  45.395000 2.805000 ;
      RECT  45.685000 -0.085000  45.855000 0.085000 ;
      RECT  45.685000  2.635000  45.855000 2.805000 ;
      RECT  45.985000  1.785000  46.155000 1.955000 ;
      RECT  46.145000 -0.085000  46.315000 0.085000 ;
      RECT  46.145000  2.635000  46.315000 2.805000 ;
      RECT  46.605000 -0.085000  46.775000 0.085000 ;
      RECT  46.605000  2.635000  46.775000 2.805000 ;
      RECT  46.925000  1.785000  47.095000 1.955000 ;
      RECT  47.065000 -0.085000  47.235000 0.085000 ;
      RECT  47.065000  2.635000  47.235000 2.805000 ;
      RECT  47.525000 -0.085000  47.695000 0.085000 ;
      RECT  47.525000  2.635000  47.695000 2.805000 ;
      RECT  47.985000 -0.085000  48.155000 0.085000 ;
      RECT  47.985000  2.635000  48.155000 2.805000 ;
      RECT  48.445000 -0.085000  48.615000 0.085000 ;
      RECT  48.445000  2.635000  48.615000 2.805000 ;
      RECT  48.905000 -0.085000  49.075000 0.085000 ;
      RECT  48.905000  2.635000  49.075000 2.805000 ;
      RECT  49.365000 -0.085000  49.535000 0.085000 ;
      RECT  49.365000  2.635000  49.535000 2.805000 ;
      RECT  49.825000 -0.085000  49.995000 0.085000 ;
      RECT  49.825000  2.635000  49.995000 2.805000 ;
      RECT  50.285000 -0.085000  50.455000 0.085000 ;
      RECT  50.285000  2.635000  50.455000 2.805000 ;
      RECT  50.745000 -0.085000  50.915000 0.085000 ;
      RECT  50.745000  2.635000  50.915000 2.805000 ;
      RECT  51.205000 -0.085000  51.375000 0.085000 ;
      RECT  51.205000  2.635000  51.375000 2.805000 ;
      RECT  51.665000 -0.085000  51.835000 0.085000 ;
      RECT  51.665000  2.635000  51.835000 2.805000 ;
      RECT  52.125000 -0.085000  52.295000 0.085000 ;
      RECT  52.125000  2.635000  52.295000 2.805000 ;
      RECT  52.585000 -0.085000  52.755000 0.085000 ;
      RECT  52.585000  2.635000  52.755000 2.805000 ;
      RECT  53.045000 -0.085000  53.215000 0.085000 ;
      RECT  53.045000  2.635000  53.215000 2.805000 ;
      RECT  53.185000  1.785000  53.355000 1.955000 ;
      RECT  53.505000 -0.085000  53.675000 0.085000 ;
      RECT  53.505000  2.635000  53.675000 2.805000 ;
      RECT  53.965000 -0.085000  54.135000 0.085000 ;
      RECT  53.965000  2.635000  54.135000 2.805000 ;
      RECT  54.125000  1.785000  54.295000 1.955000 ;
      RECT  54.425000 -0.085000  54.595000 0.085000 ;
      RECT  54.425000  2.635000  54.595000 2.805000 ;
      RECT  54.885000 -0.085000  55.055000 0.085000 ;
      RECT  54.885000  2.635000  55.055000 2.805000 ;
      RECT  55.345000 -0.085000  55.515000 0.085000 ;
      RECT  55.345000  2.635000  55.515000 2.805000 ;
      RECT  55.805000 -0.085000  55.975000 0.085000 ;
      RECT  55.805000  2.635000  55.975000 2.805000 ;
      RECT  56.265000 -0.085000  56.435000 0.085000 ;
      RECT  56.265000  2.635000  56.435000 2.805000 ;
      RECT  56.725000 -0.085000  56.895000 0.085000 ;
      RECT  56.725000  2.635000  56.895000 2.805000 ;
      RECT  57.185000 -0.085000  57.355000 0.085000 ;
      RECT  57.185000  2.635000  57.355000 2.805000 ;
      RECT  57.645000 -0.085000  57.815000 0.085000 ;
      RECT  57.645000  2.635000  57.815000 2.805000 ;
      RECT  58.105000 -0.085000  58.275000 0.085000 ;
      RECT  58.105000  2.635000  58.275000 2.805000 ;
      RECT  58.565000 -0.085000  58.735000 0.085000 ;
      RECT  58.565000  2.635000  58.735000 2.805000 ;
      RECT  58.865000  1.785000  59.035000 1.955000 ;
      RECT  59.025000 -0.085000  59.195000 0.085000 ;
      RECT  59.025000  2.635000  59.195000 2.805000 ;
      RECT  59.485000 -0.085000  59.655000 0.085000 ;
      RECT  59.485000  2.635000  59.655000 2.805000 ;
      RECT  59.805000  1.785000  59.975000 1.955000 ;
      RECT  59.945000 -0.085000  60.115000 0.085000 ;
      RECT  59.945000  2.635000  60.115000 2.805000 ;
      RECT  60.405000 -0.085000  60.575000 0.085000 ;
      RECT  60.405000  2.635000  60.575000 2.805000 ;
      RECT  60.865000 -0.085000  61.035000 0.085000 ;
      RECT  60.865000  2.635000  61.035000 2.805000 ;
      RECT  61.325000 -0.085000  61.495000 0.085000 ;
      RECT  61.325000  2.635000  61.495000 2.805000 ;
      RECT  61.785000 -0.085000  61.955000 0.085000 ;
      RECT  61.785000  2.635000  61.955000 2.805000 ;
      RECT  62.245000 -0.085000  62.415000 0.085000 ;
      RECT  62.245000  2.635000  62.415000 2.805000 ;
      RECT  62.705000 -0.085000  62.875000 0.085000 ;
      RECT  62.705000  2.635000  62.875000 2.805000 ;
      RECT  63.165000 -0.085000  63.335000 0.085000 ;
      RECT  63.165000  2.635000  63.335000 2.805000 ;
      RECT  63.625000 -0.085000  63.795000 0.085000 ;
      RECT  63.625000  2.635000  63.795000 2.805000 ;
      RECT  64.085000 -0.085000  64.255000 0.085000 ;
      RECT  64.085000  1.785000  64.255000 1.955000 ;
      RECT  64.085000  2.635000  64.255000 2.805000 ;
      RECT  64.545000 -0.085000  64.715000 0.085000 ;
      RECT  64.545000  2.635000  64.715000 2.805000 ;
      RECT  65.005000 -0.085000  65.175000 0.085000 ;
      RECT  65.005000  2.635000  65.175000 2.805000 ;
      RECT  65.465000 -0.085000  65.635000 0.085000 ;
      RECT  65.465000  2.635000  65.635000 2.805000 ;
      RECT  65.925000 -0.085000  66.095000 0.085000 ;
      RECT  65.925000  2.635000  66.095000 2.805000 ;
      RECT  66.385000 -0.085000  66.555000 0.085000 ;
      RECT  66.385000  1.785000  66.555000 1.955000 ;
      RECT  66.385000  2.635000  66.555000 2.805000 ;
      RECT  66.845000 -0.085000  67.015000 0.085000 ;
      RECT  66.845000  2.635000  67.015000 2.805000 ;
      RECT  67.305000 -0.085000  67.475000 0.085000 ;
      RECT  67.305000  2.635000  67.475000 2.805000 ;
      RECT  67.765000 -0.085000  67.935000 0.085000 ;
      RECT  67.765000  2.635000  67.935000 2.805000 ;
      RECT  68.225000 -0.085000  68.395000 0.085000 ;
      RECT  68.225000  1.785000  68.395000 1.955000 ;
      RECT  68.225000  2.635000  68.395000 2.805000 ;
      RECT  68.685000 -0.085000  68.855000 0.085000 ;
      RECT  68.685000  2.635000  68.855000 2.805000 ;
      RECT  69.145000 -0.085000  69.315000 0.085000 ;
      RECT  69.145000  2.635000  69.315000 2.805000 ;
      RECT  69.605000 -0.085000  69.775000 0.085000 ;
      RECT  69.605000  2.635000  69.775000 2.805000 ;
      RECT  70.065000 -0.085000  70.235000 0.085000 ;
      RECT  70.065000  2.635000  70.235000 2.805000 ;
      RECT  70.525000 -0.085000  70.695000 0.085000 ;
      RECT  70.525000  1.785000  70.695000 1.955000 ;
      RECT  70.525000  2.635000  70.695000 2.805000 ;
      RECT  70.985000 -0.085000  71.155000 0.085000 ;
      RECT  70.985000  2.635000  71.155000 2.805000 ;
      RECT  71.445000 -0.085000  71.615000 0.085000 ;
      RECT  71.445000  2.635000  71.615000 2.805000 ;
      RECT  71.905000 -0.085000  72.075000 0.085000 ;
      RECT  71.905000  2.635000  72.075000 2.805000 ;
      RECT  72.365000 -0.085000  72.535000 0.085000 ;
      RECT  72.365000  1.785000  72.535000 1.955000 ;
      RECT  72.365000  2.635000  72.535000 2.805000 ;
      RECT  72.825000 -0.085000  72.995000 0.085000 ;
      RECT  72.825000  2.635000  72.995000 2.805000 ;
      RECT  73.285000 -0.085000  73.455000 0.085000 ;
      RECT  73.285000  2.635000  73.455000 2.805000 ;
      RECT  73.745000 -0.085000  73.915000 0.085000 ;
      RECT  73.745000  2.635000  73.915000 2.805000 ;
      RECT  74.205000 -0.085000  74.375000 0.085000 ;
      RECT  74.205000  2.635000  74.375000 2.805000 ;
      RECT  74.665000 -0.085000  74.835000 0.085000 ;
      RECT  74.665000  1.785000  74.835000 1.955000 ;
      RECT  74.665000  2.635000  74.835000 2.805000 ;
      RECT  75.125000 -0.085000  75.295000 0.085000 ;
      RECT  75.125000  2.635000  75.295000 2.805000 ;
      RECT  75.585000 -0.085000  75.755000 0.085000 ;
      RECT  75.585000  2.635000  75.755000 2.805000 ;
      RECT  76.045000 -0.085000  76.215000 0.085000 ;
      RECT  76.045000  2.635000  76.215000 2.805000 ;
      RECT  76.505000 -0.085000  76.675000 0.085000 ;
      RECT  76.505000  1.785000  76.675000 1.955000 ;
      RECT  76.505000  2.635000  76.675000 2.805000 ;
      RECT  76.965000 -0.085000  77.135000 0.085000 ;
      RECT  76.965000  2.635000  77.135000 2.805000 ;
      RECT  77.425000 -0.085000  77.595000 0.085000 ;
      RECT  77.425000  2.635000  77.595000 2.805000 ;
      RECT  77.885000 -0.085000  78.055000 0.085000 ;
      RECT  77.885000  2.635000  78.055000 2.805000 ;
      RECT  78.345000 -0.085000  78.515000 0.085000 ;
      RECT  78.345000  2.635000  78.515000 2.805000 ;
      RECT  78.805000 -0.085000  78.975000 0.085000 ;
      RECT  78.805000  1.785000  78.975000 1.955000 ;
      RECT  78.805000  2.635000  78.975000 2.805000 ;
      RECT  79.265000 -0.085000  79.435000 0.085000 ;
      RECT  79.265000  2.635000  79.435000 2.805000 ;
      RECT  79.725000 -0.085000  79.895000 0.085000 ;
      RECT  79.725000  2.635000  79.895000 2.805000 ;
      RECT  80.185000 -0.085000  80.355000 0.085000 ;
      RECT  80.185000  2.635000  80.355000 2.805000 ;
      RECT  80.645000 -0.085000  80.815000 0.085000 ;
      RECT  80.645000  2.635000  80.815000 2.805000 ;
      RECT  81.105000 -0.085000  81.275000 0.085000 ;
      RECT  81.105000  2.635000  81.275000 2.805000 ;
      RECT  81.565000 -0.085000  81.735000 0.085000 ;
      RECT  81.565000  1.785000  81.735000 1.955000 ;
      RECT  81.565000  2.635000  81.735000 2.805000 ;
      RECT  82.025000 -0.085000  82.195000 0.085000 ;
      RECT  82.025000  2.635000  82.195000 2.805000 ;
      RECT  82.485000 -0.085000  82.655000 0.085000 ;
      RECT  82.485000  2.635000  82.655000 2.805000 ;
      RECT  82.945000 -0.085000  83.115000 0.085000 ;
      RECT  82.945000  2.635000  83.115000 2.805000 ;
      RECT  83.405000 -0.085000  83.575000 0.085000 ;
      RECT  83.405000  2.635000  83.575000 2.805000 ;
      RECT  83.865000 -0.085000  84.035000 0.085000 ;
      RECT  83.865000  2.635000  84.035000 2.805000 ;
      RECT  84.325000 -0.085000  84.495000 0.085000 ;
      RECT  84.325000  2.635000  84.495000 2.805000 ;
      RECT  84.785000 -0.085000  84.955000 0.085000 ;
      RECT  84.785000  1.785000  84.955000 1.955000 ;
      RECT  84.785000  2.635000  84.955000 2.805000 ;
      RECT  85.245000 -0.085000  85.415000 0.085000 ;
      RECT  85.245000  2.635000  85.415000 2.805000 ;
      RECT  85.705000 -0.085000  85.875000 0.085000 ;
      RECT  85.705000  2.635000  85.875000 2.805000 ;
      RECT  86.165000 -0.085000  86.335000 0.085000 ;
      RECT  86.165000  2.635000  86.335000 2.805000 ;
      RECT  86.625000 -0.085000  86.795000 0.085000 ;
      RECT  86.625000  2.635000  86.795000 2.805000 ;
      RECT  87.085000 -0.085000  87.255000 0.085000 ;
      RECT  87.085000  2.635000  87.255000 2.805000 ;
      RECT  87.545000 -0.085000  87.715000 0.085000 ;
      RECT  87.545000  2.635000  87.715000 2.805000 ;
      RECT  88.005000 -0.085000  88.175000 0.085000 ;
      RECT  88.005000  1.785000  88.175000 1.955000 ;
      RECT  88.005000  2.635000  88.175000 2.805000 ;
      RECT  88.465000 -0.085000  88.635000 0.085000 ;
      RECT  88.465000  2.635000  88.635000 2.805000 ;
      RECT  88.925000 -0.085000  89.095000 0.085000 ;
      RECT  88.925000  2.635000  89.095000 2.805000 ;
      RECT  89.385000 -0.085000  89.555000 0.085000 ;
      RECT  89.385000  2.635000  89.555000 2.805000 ;
      RECT  89.845000 -0.085000  90.015000 0.085000 ;
      RECT  89.845000  2.635000  90.015000 2.805000 ;
      RECT  90.305000 -0.085000  90.475000 0.085000 ;
      RECT  90.305000  2.635000  90.475000 2.805000 ;
      RECT  90.765000 -0.085000  90.935000 0.085000 ;
      RECT  90.765000  2.635000  90.935000 2.805000 ;
      RECT  91.225000 -0.085000  91.395000 0.085000 ;
      RECT  91.225000  1.785000  91.395000 1.955000 ;
      RECT  91.225000  2.635000  91.395000 2.805000 ;
      RECT  91.685000 -0.085000  91.855000 0.085000 ;
      RECT  91.685000  2.635000  91.855000 2.805000 ;
      RECT  92.145000 -0.085000  92.315000 0.085000 ;
      RECT  92.145000  2.635000  92.315000 2.805000 ;
      RECT  92.605000 -0.085000  92.775000 0.085000 ;
      RECT  92.605000  2.635000  92.775000 2.805000 ;
      RECT  93.065000 -0.085000  93.235000 0.085000 ;
      RECT  93.065000  2.635000  93.235000 2.805000 ;
      RECT  93.525000 -0.085000  93.695000 0.085000 ;
      RECT  93.525000  2.635000  93.695000 2.805000 ;
      RECT  93.985000 -0.085000  94.155000 0.085000 ;
      RECT  93.985000  2.635000  94.155000 2.805000 ;
      RECT  94.445000 -0.085000  94.615000 0.085000 ;
      RECT  94.445000  1.785000  94.615000 1.955000 ;
      RECT  94.445000  2.635000  94.615000 2.805000 ;
      RECT  94.905000 -0.085000  95.075000 0.085000 ;
      RECT  94.905000  2.635000  95.075000 2.805000 ;
      RECT  95.365000 -0.085000  95.535000 0.085000 ;
      RECT  95.365000  2.635000  95.535000 2.805000 ;
      RECT  95.825000 -0.085000  95.995000 0.085000 ;
      RECT  95.825000  2.635000  95.995000 2.805000 ;
      RECT  96.285000 -0.085000  96.455000 0.085000 ;
      RECT  96.285000  2.635000  96.455000 2.805000 ;
      RECT  96.745000 -0.085000  96.915000 0.085000 ;
      RECT  96.745000  2.635000  96.915000 2.805000 ;
      RECT  97.205000 -0.085000  97.375000 0.085000 ;
      RECT  97.205000  2.635000  97.375000 2.805000 ;
      RECT  97.665000 -0.085000  97.835000 0.085000 ;
      RECT  97.665000  1.785000  97.835000 1.955000 ;
      RECT  97.665000  2.635000  97.835000 2.805000 ;
      RECT  98.125000 -0.085000  98.295000 0.085000 ;
      RECT  98.125000  2.635000  98.295000 2.805000 ;
      RECT  98.585000 -0.085000  98.755000 0.085000 ;
      RECT  98.585000  2.635000  98.755000 2.805000 ;
      RECT  99.045000 -0.085000  99.215000 0.085000 ;
      RECT  99.045000  2.635000  99.215000 2.805000 ;
      RECT  99.505000 -0.085000  99.675000 0.085000 ;
      RECT  99.505000  2.635000  99.675000 2.805000 ;
      RECT  99.965000 -0.085000 100.135000 0.085000 ;
      RECT  99.965000  2.635000 100.135000 2.805000 ;
      RECT 100.425000 -0.085000 100.595000 0.085000 ;
      RECT 100.425000  2.635000 100.595000 2.805000 ;
      RECT 100.885000 -0.085000 101.055000 0.085000 ;
      RECT 100.885000  1.785000 101.055000 1.955000 ;
      RECT 100.885000  2.635000 101.055000 2.805000 ;
      RECT 101.345000 -0.085000 101.515000 0.085000 ;
      RECT 101.345000  2.635000 101.515000 2.805000 ;
      RECT 101.805000 -0.085000 101.975000 0.085000 ;
      RECT 101.805000  2.635000 101.975000 2.805000 ;
      RECT 102.265000 -0.085000 102.435000 0.085000 ;
      RECT 102.265000  2.635000 102.435000 2.805000 ;
      RECT 102.725000 -0.085000 102.895000 0.085000 ;
      RECT 102.725000  2.635000 102.895000 2.805000 ;
      RECT 103.185000 -0.085000 103.355000 0.085000 ;
      RECT 103.185000  2.635000 103.355000 2.805000 ;
      RECT 103.645000 -0.085000 103.815000 0.085000 ;
      RECT 103.645000  2.635000 103.815000 2.805000 ;
      RECT 104.105000 -0.085000 104.275000 0.085000 ;
      RECT 104.105000  1.785000 104.275000 1.955000 ;
      RECT 104.105000  2.635000 104.275000 2.805000 ;
      RECT 104.565000 -0.085000 104.735000 0.085000 ;
      RECT 104.565000  2.635000 104.735000 2.805000 ;
      RECT 105.025000 -0.085000 105.195000 0.085000 ;
      RECT 105.025000  2.635000 105.195000 2.805000 ;
      RECT 105.485000 -0.085000 105.655000 0.085000 ;
      RECT 105.485000  2.635000 105.655000 2.805000 ;
      RECT 105.945000 -0.085000 106.115000 0.085000 ;
      RECT 105.945000  2.635000 106.115000 2.805000 ;
      RECT 105.945000  5.355000 106.115000 5.525000 ;
      RECT 106.405000 -0.085000 106.575000 0.085000 ;
      RECT 106.405000  2.635000 106.575000 2.805000 ;
      RECT 106.405000  5.355000 106.575000 5.525000 ;
      RECT 106.865000 -0.085000 107.035000 0.085000 ;
      RECT 106.865000  2.635000 107.035000 2.805000 ;
      RECT 106.865000  5.355000 107.035000 5.525000 ;
      RECT 107.325000 -0.085000 107.495000 0.085000 ;
      RECT 107.325000  2.635000 107.495000 2.805000 ;
      RECT 107.325000  5.355000 107.495000 5.525000 ;
      RECT 107.605000  2.140000 107.775000 2.310000 ;
      RECT 107.605000  3.130000 107.775000 3.300000 ;
      RECT 107.785000 -0.085000 107.955000 0.085000 ;
      RECT 107.785000  5.355000 107.955000 5.525000 ;
      RECT 108.085000  1.785000 108.255000 1.955000 ;
      RECT 108.085000  3.485000 108.255000 3.655000 ;
      RECT 108.245000 -0.085000 108.415000 0.085000 ;
      RECT 108.245000  5.355000 108.415000 5.525000 ;
      RECT 108.555000  2.140000 108.725000 2.310000 ;
      RECT 108.555000  3.130000 108.725000 3.300000 ;
      RECT 108.705000 -0.085000 108.875000 0.085000 ;
      RECT 108.705000  5.355000 108.875000 5.525000 ;
      RECT 109.025000  1.785000 109.195000 1.955000 ;
      RECT 109.025000  3.485000 109.195000 3.655000 ;
      RECT 109.165000 -0.085000 109.335000 0.085000 ;
      RECT 109.165000  5.355000 109.335000 5.525000 ;
      RECT 109.505000  2.140000 109.675000 2.310000 ;
      RECT 109.505000  3.130000 109.675000 3.300000 ;
      RECT 109.625000 -0.085000 109.795000 0.085000 ;
      RECT 109.625000  2.635000 109.795000 2.805000 ;
      RECT 109.625000  5.355000 109.795000 5.525000 ;
      RECT 110.085000 -0.085000 110.255000 0.085000 ;
      RECT 110.085000  2.635000 110.255000 2.805000 ;
      RECT 110.085000  5.355000 110.255000 5.525000 ;
      RECT 110.485000  2.140000 110.655000 2.310000 ;
      RECT 110.485000  3.130000 110.655000 3.300000 ;
      RECT 110.545000 -0.085000 110.715000 0.085000 ;
      RECT 110.545000  2.635000 110.715000 2.805000 ;
      RECT 110.545000  5.355000 110.715000 5.525000 ;
      RECT 111.005000 -0.085000 111.175000 0.085000 ;
      RECT 111.005000  2.635000 111.175000 2.805000 ;
      RECT 111.005000  5.355000 111.175000 5.525000 ;
      RECT 111.425000  2.140000 111.595000 2.310000 ;
      RECT 111.425000  3.130000 111.595000 3.300000 ;
      RECT 111.465000 -0.085000 111.635000 0.085000 ;
      RECT 111.465000  2.635000 111.635000 2.805000 ;
      RECT 111.465000  5.355000 111.635000 5.525000 ;
      RECT 111.925000 -0.085000 112.095000 0.085000 ;
      RECT 111.925000  2.635000 112.095000 2.805000 ;
      RECT 111.925000  5.355000 112.095000 5.525000 ;
      RECT 112.385000 -0.085000 112.555000 0.085000 ;
      RECT 112.385000  2.635000 112.555000 2.805000 ;
      RECT 112.385000  5.355000 112.555000 5.525000 ;
      RECT 112.425000  2.140000 112.595000 2.310000 ;
      RECT 112.425000  3.130000 112.595000 3.300000 ;
      RECT 112.845000 -0.085000 113.015000 0.085000 ;
      RECT 112.845000  2.635000 113.015000 2.805000 ;
      RECT 112.845000  5.355000 113.015000 5.525000 ;
      RECT 113.305000 -0.085000 113.475000 0.085000 ;
      RECT 113.305000  2.635000 113.475000 2.805000 ;
      RECT 113.305000  5.355000 113.475000 5.525000 ;
      RECT 113.365000  2.140000 113.535000 2.310000 ;
      RECT 113.365000  3.130000 113.535000 3.300000 ;
      RECT 113.765000 -0.085000 113.935000 0.085000 ;
      RECT 113.765000  2.635000 113.935000 2.805000 ;
      RECT 113.765000  5.355000 113.935000 5.525000 ;
      RECT 114.225000 -0.085000 114.395000 0.085000 ;
      RECT 114.225000  2.635000 114.395000 2.805000 ;
      RECT 114.225000  5.355000 114.395000 5.525000 ;
      RECT 114.345000  2.140000 114.515000 2.310000 ;
      RECT 114.345000  3.130000 114.515000 3.300000 ;
      RECT 114.685000 -0.085000 114.855000 0.085000 ;
      RECT 114.685000  5.355000 114.855000 5.525000 ;
      RECT 114.825000  1.785000 114.995000 1.955000 ;
      RECT 114.825000  3.485000 114.995000 3.655000 ;
      RECT 115.145000 -0.085000 115.315000 0.085000 ;
      RECT 115.145000  5.355000 115.315000 5.525000 ;
      RECT 115.295000  2.140000 115.465000 2.310000 ;
      RECT 115.295000  3.130000 115.465000 3.300000 ;
      RECT 115.605000 -0.085000 115.775000 0.085000 ;
      RECT 115.605000  5.355000 115.775000 5.525000 ;
      RECT 115.765000  1.785000 115.935000 1.955000 ;
      RECT 115.765000  3.485000 115.935000 3.655000 ;
      RECT 116.065000 -0.085000 116.235000 0.085000 ;
      RECT 116.065000  5.355000 116.235000 5.525000 ;
      RECT 116.245000  2.140000 116.415000 2.310000 ;
      RECT 116.245000  3.130000 116.415000 3.300000 ;
      RECT 116.525000 -0.085000 116.695000 0.085000 ;
      RECT 116.525000  2.635000 116.695000 2.805000 ;
      RECT 116.525000  5.355000 116.695000 5.525000 ;
      RECT 116.985000 -0.085000 117.155000 0.085000 ;
      RECT 116.985000  2.635000 117.155000 2.805000 ;
      RECT 116.985000  5.355000 117.155000 5.525000 ;
      RECT 117.445000 -0.085000 117.615000 0.085000 ;
      RECT 117.445000  2.635000 117.615000 2.805000 ;
      RECT 117.445000  5.355000 117.615000 5.525000 ;
      RECT 117.905000 -0.085000 118.075000 0.085000 ;
      RECT 117.905000  2.635000 118.075000 2.805000 ;
      RECT 117.905000  5.355000 118.075000 5.525000 ;
      RECT 118.365000 -0.085000 118.535000 0.085000 ;
      RECT 118.365000  2.635000 118.535000 2.805000 ;
      RECT 118.365000  5.355000 118.535000 5.525000 ;
      RECT 118.825000 -0.085000 118.995000 0.085000 ;
      RECT 118.825000  2.635000 118.995000 2.805000 ;
      RECT 118.825000  5.355000 118.995000 5.525000 ;
      RECT 119.285000 -0.085000 119.455000 0.085000 ;
      RECT 119.285000  2.635000 119.455000 2.805000 ;
      RECT 119.285000  5.355000 119.455000 5.525000 ;
      RECT 119.745000 -0.085000 119.915000 0.085000 ;
      RECT 119.745000  2.635000 119.915000 2.805000 ;
      RECT 119.745000  5.355000 119.915000 5.525000 ;
      RECT 120.025000  2.140000 120.195000 2.310000 ;
      RECT 120.025000  3.130000 120.195000 3.300000 ;
      RECT 120.205000 -0.085000 120.375000 0.085000 ;
      RECT 120.205000  5.355000 120.375000 5.525000 ;
      RECT 120.505000  1.785000 120.675000 1.955000 ;
      RECT 120.505000  3.485000 120.675000 3.655000 ;
      RECT 120.665000 -0.085000 120.835000 0.085000 ;
      RECT 120.665000  5.355000 120.835000 5.525000 ;
      RECT 120.975000  2.140000 121.145000 2.310000 ;
      RECT 120.975000  3.130000 121.145000 3.300000 ;
      RECT 121.125000 -0.085000 121.295000 0.085000 ;
      RECT 121.125000  5.355000 121.295000 5.525000 ;
      RECT 121.445000  1.785000 121.615000 1.955000 ;
      RECT 121.445000  3.485000 121.615000 3.655000 ;
      RECT 121.585000 -0.085000 121.755000 0.085000 ;
      RECT 121.585000  5.355000 121.755000 5.525000 ;
      RECT 121.925000  2.140000 122.095000 2.310000 ;
      RECT 121.925000  3.130000 122.095000 3.300000 ;
      RECT 122.045000 -0.085000 122.215000 0.085000 ;
      RECT 122.045000  2.635000 122.215000 2.805000 ;
      RECT 122.045000  5.355000 122.215000 5.525000 ;
      RECT 122.505000 -0.085000 122.675000 0.085000 ;
      RECT 122.505000  2.635000 122.675000 2.805000 ;
      RECT 122.505000  5.355000 122.675000 5.525000 ;
      RECT 122.905000  2.140000 123.075000 2.310000 ;
      RECT 122.905000  3.130000 123.075000 3.300000 ;
      RECT 122.965000 -0.085000 123.135000 0.085000 ;
      RECT 122.965000  2.635000 123.135000 2.805000 ;
      RECT 122.965000  5.355000 123.135000 5.525000 ;
      RECT 123.425000 -0.085000 123.595000 0.085000 ;
      RECT 123.425000  2.635000 123.595000 2.805000 ;
      RECT 123.425000  5.355000 123.595000 5.525000 ;
      RECT 123.845000  2.140000 124.015000 2.310000 ;
      RECT 123.845000  3.130000 124.015000 3.300000 ;
      RECT 123.885000 -0.085000 124.055000 0.085000 ;
      RECT 123.885000  2.635000 124.055000 2.805000 ;
      RECT 123.885000  5.355000 124.055000 5.525000 ;
      RECT 124.345000 -0.085000 124.515000 0.085000 ;
      RECT 124.345000  2.635000 124.515000 2.805000 ;
      RECT 124.345000  5.355000 124.515000 5.525000 ;
      RECT 124.805000 -0.085000 124.975000 0.085000 ;
      RECT 124.805000  2.635000 124.975000 2.805000 ;
      RECT 124.805000  5.355000 124.975000 5.525000 ;
      RECT 124.845000  2.140000 125.015000 2.310000 ;
      RECT 124.845000  3.130000 125.015000 3.300000 ;
      RECT 125.265000 -0.085000 125.435000 0.085000 ;
      RECT 125.265000  2.635000 125.435000 2.805000 ;
      RECT 125.265000  5.355000 125.435000 5.525000 ;
      RECT 125.725000 -0.085000 125.895000 0.085000 ;
      RECT 125.725000  2.635000 125.895000 2.805000 ;
      RECT 125.725000  5.355000 125.895000 5.525000 ;
      RECT 125.785000  2.140000 125.955000 2.310000 ;
      RECT 125.785000  3.130000 125.955000 3.300000 ;
      RECT 126.185000 -0.085000 126.355000 0.085000 ;
      RECT 126.185000  2.635000 126.355000 2.805000 ;
      RECT 126.185000  5.355000 126.355000 5.525000 ;
      RECT 126.645000 -0.085000 126.815000 0.085000 ;
      RECT 126.645000  2.635000 126.815000 2.805000 ;
      RECT 126.645000  5.355000 126.815000 5.525000 ;
      RECT 126.765000  2.140000 126.935000 2.310000 ;
      RECT 126.765000  3.130000 126.935000 3.300000 ;
      RECT 127.105000 -0.085000 127.275000 0.085000 ;
      RECT 127.105000  5.355000 127.275000 5.525000 ;
      RECT 127.245000  1.785000 127.415000 1.955000 ;
      RECT 127.245000  3.485000 127.415000 3.655000 ;
      RECT 127.565000 -0.085000 127.735000 0.085000 ;
      RECT 127.565000  5.355000 127.735000 5.525000 ;
      RECT 127.715000  2.140000 127.885000 2.310000 ;
      RECT 127.715000  3.130000 127.885000 3.300000 ;
      RECT 128.025000 -0.085000 128.195000 0.085000 ;
      RECT 128.025000  5.355000 128.195000 5.525000 ;
      RECT 128.185000  1.785000 128.355000 1.955000 ;
      RECT 128.185000  3.485000 128.355000 3.655000 ;
      RECT 128.485000 -0.085000 128.655000 0.085000 ;
      RECT 128.485000  5.355000 128.655000 5.525000 ;
      RECT 128.665000  2.140000 128.835000 2.310000 ;
      RECT 128.665000  3.130000 128.835000 3.300000 ;
      RECT 128.945000 -0.085000 129.115000 0.085000 ;
      RECT 128.945000  2.635000 129.115000 2.805000 ;
      RECT 128.945000  5.355000 129.115000 5.525000 ;
      RECT 129.405000 -0.085000 129.575000 0.085000 ;
      RECT 129.405000  2.635000 129.575000 2.805000 ;
      RECT 129.405000  5.355000 129.575000 5.525000 ;
      RECT 129.865000 -0.085000 130.035000 0.085000 ;
      RECT 129.865000  2.635000 130.035000 2.805000 ;
      RECT 129.865000  5.355000 130.035000 5.525000 ;
      RECT 130.325000 -0.085000 130.495000 0.085000 ;
      RECT 130.325000  2.635000 130.495000 2.805000 ;
      RECT 130.325000  5.355000 130.495000 5.525000 ;
      RECT 130.785000 -0.085000 130.955000 0.085000 ;
      RECT 130.785000  2.635000 130.955000 2.805000 ;
      RECT 130.785000  5.355000 130.955000 5.525000 ;
      RECT 131.245000 -0.085000 131.415000 0.085000 ;
      RECT 131.245000  2.635000 131.415000 2.805000 ;
      RECT 131.245000  5.355000 131.415000 5.525000 ;
      RECT 131.705000 -0.085000 131.875000 0.085000 ;
      RECT 131.705000  1.785000 131.875000 1.955000 ;
      RECT 131.705000  3.485000 131.875000 3.655000 ;
      RECT 131.705000  5.355000 131.875000 5.525000 ;
      RECT 132.165000 -0.085000 132.335000 0.085000 ;
      RECT 132.165000  2.635000 132.335000 2.805000 ;
      RECT 132.165000  5.355000 132.335000 5.525000 ;
      RECT 132.625000 -0.085000 132.795000 0.085000 ;
      RECT 132.625000  2.635000 132.795000 2.805000 ;
      RECT 132.625000  5.355000 132.795000 5.525000 ;
      RECT 133.085000 -0.085000 133.255000 0.085000 ;
      RECT 133.085000  2.635000 133.255000 2.805000 ;
      RECT 133.085000  5.355000 133.255000 5.525000 ;
      RECT 133.545000 -0.085000 133.715000 0.085000 ;
      RECT 133.545000  2.635000 133.715000 2.805000 ;
      RECT 133.545000  5.355000 133.715000 5.525000 ;
      RECT 134.005000 -0.085000 134.175000 0.085000 ;
      RECT 134.005000  1.785000 134.175000 1.955000 ;
      RECT 134.005000  3.485000 134.175000 3.655000 ;
      RECT 134.005000  5.355000 134.175000 5.525000 ;
      RECT 134.465000 -0.085000 134.635000 0.085000 ;
      RECT 134.465000  2.635000 134.635000 2.805000 ;
      RECT 134.465000  5.355000 134.635000 5.525000 ;
      RECT 134.925000 -0.085000 135.095000 0.085000 ;
      RECT 134.925000  2.635000 135.095000 2.805000 ;
      RECT 134.925000  5.355000 135.095000 5.525000 ;
      RECT 135.385000 -0.085000 135.555000 0.085000 ;
      RECT 135.385000  2.635000 135.555000 2.805000 ;
      RECT 135.385000  5.355000 135.555000 5.525000 ;
      RECT 135.845000 -0.085000 136.015000 0.085000 ;
      RECT 135.845000  1.785000 136.015000 1.955000 ;
      RECT 135.845000  3.485000 136.015000 3.655000 ;
      RECT 135.845000  5.355000 136.015000 5.525000 ;
      RECT 136.305000 -0.085000 136.475000 0.085000 ;
      RECT 136.305000  2.635000 136.475000 2.805000 ;
      RECT 136.305000  5.355000 136.475000 5.525000 ;
      RECT 136.765000 -0.085000 136.935000 0.085000 ;
      RECT 136.765000  2.635000 136.935000 2.805000 ;
      RECT 136.765000  5.355000 136.935000 5.525000 ;
      RECT 137.225000 -0.085000 137.395000 0.085000 ;
      RECT 137.225000  2.635000 137.395000 2.805000 ;
      RECT 137.225000  5.355000 137.395000 5.525000 ;
      RECT 137.685000 -0.085000 137.855000 0.085000 ;
      RECT 137.685000  2.635000 137.855000 2.805000 ;
      RECT 137.685000  5.355000 137.855000 5.525000 ;
      RECT 138.145000 -0.085000 138.315000 0.085000 ;
      RECT 138.145000  1.785000 138.315000 1.955000 ;
      RECT 138.145000  3.485000 138.315000 3.655000 ;
      RECT 138.145000  5.355000 138.315000 5.525000 ;
      RECT 138.605000 -0.085000 138.775000 0.085000 ;
      RECT 138.605000  2.635000 138.775000 2.805000 ;
      RECT 138.605000  5.355000 138.775000 5.525000 ;
      RECT 139.065000 -0.085000 139.235000 0.085000 ;
      RECT 139.065000  2.635000 139.235000 2.805000 ;
      RECT 139.065000  5.355000 139.235000 5.525000 ;
      RECT 139.525000 -0.085000 139.695000 0.085000 ;
      RECT 139.525000  2.635000 139.695000 2.805000 ;
      RECT 139.525000  5.355000 139.695000 5.525000 ;
      RECT 139.985000 -0.085000 140.155000 0.085000 ;
      RECT 139.985000  1.785000 140.155000 1.955000 ;
      RECT 139.985000  3.485000 140.155000 3.655000 ;
      RECT 139.985000  5.355000 140.155000 5.525000 ;
      RECT 140.445000 -0.085000 140.615000 0.085000 ;
      RECT 140.445000  2.635000 140.615000 2.805000 ;
      RECT 140.445000  5.355000 140.615000 5.525000 ;
      RECT 140.905000 -0.085000 141.075000 0.085000 ;
      RECT 140.905000  2.635000 141.075000 2.805000 ;
      RECT 140.905000  5.355000 141.075000 5.525000 ;
      RECT 141.365000 -0.085000 141.535000 0.085000 ;
      RECT 141.365000  2.635000 141.535000 2.805000 ;
      RECT 141.365000  5.355000 141.535000 5.525000 ;
      RECT 141.825000 -0.085000 141.995000 0.085000 ;
      RECT 141.825000  2.635000 141.995000 2.805000 ;
      RECT 141.825000  5.355000 141.995000 5.525000 ;
      RECT 142.285000 -0.085000 142.455000 0.085000 ;
      RECT 142.285000  1.785000 142.455000 1.955000 ;
      RECT 142.285000  3.485000 142.455000 3.655000 ;
      RECT 142.285000  5.355000 142.455000 5.525000 ;
      RECT 142.745000 -0.085000 142.915000 0.085000 ;
      RECT 142.745000  2.635000 142.915000 2.805000 ;
      RECT 142.745000  5.355000 142.915000 5.525000 ;
      RECT 143.205000 -0.085000 143.375000 0.085000 ;
      RECT 143.205000  2.635000 143.375000 2.805000 ;
      RECT 143.205000  5.355000 143.375000 5.525000 ;
      RECT 143.665000 -0.085000 143.835000 0.085000 ;
      RECT 143.665000  2.635000 143.835000 2.805000 ;
      RECT 143.665000  5.355000 143.835000 5.525000 ;
      RECT 144.125000 -0.085000 144.295000 0.085000 ;
      RECT 144.125000  1.785000 144.295000 1.955000 ;
      RECT 144.125000  3.485000 144.295000 3.655000 ;
      RECT 144.125000  5.355000 144.295000 5.525000 ;
      RECT 144.585000 -0.085000 144.755000 0.085000 ;
      RECT 144.585000  2.635000 144.755000 2.805000 ;
      RECT 144.585000  5.355000 144.755000 5.525000 ;
      RECT 145.045000 -0.085000 145.215000 0.085000 ;
      RECT 145.045000  2.635000 145.215000 2.805000 ;
      RECT 145.045000  5.355000 145.215000 5.525000 ;
      RECT 145.505000 -0.085000 145.675000 0.085000 ;
      RECT 145.505000  2.635000 145.675000 2.805000 ;
      RECT 145.505000  5.355000 145.675000 5.525000 ;
      RECT 145.965000 -0.085000 146.135000 0.085000 ;
      RECT 145.965000  2.635000 146.135000 2.805000 ;
      RECT 145.965000  5.355000 146.135000 5.525000 ;
      RECT 146.425000 -0.085000 146.595000 0.085000 ;
      RECT 146.425000  1.785000 146.595000 1.955000 ;
      RECT 146.425000  3.485000 146.595000 3.655000 ;
      RECT 146.425000  5.355000 146.595000 5.525000 ;
      RECT 146.885000 -0.085000 147.055000 0.085000 ;
      RECT 146.885000  2.635000 147.055000 2.805000 ;
      RECT 146.885000  5.355000 147.055000 5.525000 ;
      RECT 147.345000 -0.085000 147.515000 0.085000 ;
      RECT 147.345000  2.635000 147.515000 2.805000 ;
      RECT 147.345000  5.355000 147.515000 5.525000 ;
      RECT 147.805000 -0.085000 147.975000 0.085000 ;
      RECT 147.805000  2.635000 147.975000 2.805000 ;
      RECT 147.805000  5.355000 147.975000 5.525000 ;
      RECT 147.835000  2.140000 148.005000 2.310000 ;
      RECT 147.835000  3.130000 148.005000 3.300000 ;
      RECT 148.265000 -0.085000 148.435000 0.085000 ;
      RECT 148.265000  2.635000 148.435000 2.805000 ;
      RECT 148.265000  5.355000 148.435000 5.525000 ;
      RECT 148.725000 -0.085000 148.895000 0.085000 ;
      RECT 148.725000  2.635000 148.895000 2.805000 ;
      RECT 148.725000  5.355000 148.895000 5.525000 ;
      RECT 148.775000  2.140000 148.945000 2.310000 ;
      RECT 148.775000  3.130000 148.945000 3.300000 ;
      RECT 149.185000 -0.085000 149.355000 0.085000 ;
      RECT 149.185000  1.785000 149.355000 1.955000 ;
      RECT 149.185000  3.485000 149.355000 3.655000 ;
      RECT 149.185000  5.355000 149.355000 5.525000 ;
      RECT 149.645000 -0.085000 149.815000 0.085000 ;
      RECT 149.645000  2.635000 149.815000 2.805000 ;
      RECT 149.645000  5.355000 149.815000 5.525000 ;
      RECT 149.770000  2.140000 149.940000 2.310000 ;
      RECT 149.770000  3.130000 149.940000 3.300000 ;
      RECT 150.105000 -0.085000 150.275000 0.085000 ;
      RECT 150.105000  2.635000 150.275000 2.805000 ;
      RECT 150.105000  5.355000 150.275000 5.525000 ;
      RECT 150.565000 -0.085000 150.735000 0.085000 ;
      RECT 150.565000  2.635000 150.735000 2.805000 ;
      RECT 150.565000  5.355000 150.735000 5.525000 ;
      RECT 151.025000 -0.085000 151.195000 0.085000 ;
      RECT 151.025000  2.635000 151.195000 2.805000 ;
      RECT 151.025000  5.355000 151.195000 5.525000 ;
      RECT 151.485000 -0.085000 151.655000 0.085000 ;
      RECT 151.485000  2.635000 151.655000 2.805000 ;
      RECT 151.485000  5.355000 151.655000 5.525000 ;
      RECT 151.820000  2.140000 151.990000 2.310000 ;
      RECT 151.820000  3.130000 151.990000 3.300000 ;
      RECT 151.945000 -0.085000 152.115000 0.085000 ;
      RECT 151.945000  2.635000 152.115000 2.805000 ;
      RECT 151.945000  5.355000 152.115000 5.525000 ;
      RECT 152.405000 -0.085000 152.575000 0.085000 ;
      RECT 152.405000  1.785000 152.575000 1.955000 ;
      RECT 152.405000  3.485000 152.575000 3.655000 ;
      RECT 152.405000  5.355000 152.575000 5.525000 ;
      RECT 152.815000  2.140000 152.985000 2.310000 ;
      RECT 152.815000  3.130000 152.985000 3.300000 ;
      RECT 152.865000 -0.085000 153.035000 0.085000 ;
      RECT 152.865000  2.635000 153.035000 2.805000 ;
      RECT 152.865000  5.355000 153.035000 5.525000 ;
      RECT 153.325000 -0.085000 153.495000 0.085000 ;
      RECT 153.325000  2.635000 153.495000 2.805000 ;
      RECT 153.325000  5.355000 153.495000 5.525000 ;
      RECT 153.755000  2.140000 153.925000 2.310000 ;
      RECT 153.755000  3.130000 153.925000 3.300000 ;
      RECT 153.785000 -0.085000 153.955000 0.085000 ;
      RECT 153.785000  2.635000 153.955000 2.805000 ;
      RECT 153.785000  5.355000 153.955000 5.525000 ;
      RECT 154.245000 -0.085000 154.415000 0.085000 ;
      RECT 154.245000  2.635000 154.415000 2.805000 ;
      RECT 154.245000  5.355000 154.415000 5.525000 ;
      RECT 154.275000  2.140000 154.445000 2.310000 ;
      RECT 154.275000  3.130000 154.445000 3.300000 ;
      RECT 154.705000 -0.085000 154.875000 0.085000 ;
      RECT 154.705000  2.635000 154.875000 2.805000 ;
      RECT 154.705000  5.355000 154.875000 5.525000 ;
      RECT 155.165000 -0.085000 155.335000 0.085000 ;
      RECT 155.165000  2.635000 155.335000 2.805000 ;
      RECT 155.165000  5.355000 155.335000 5.525000 ;
      RECT 155.215000  2.140000 155.385000 2.310000 ;
      RECT 155.215000  3.130000 155.385000 3.300000 ;
      RECT 155.625000 -0.085000 155.795000 0.085000 ;
      RECT 155.625000  1.785000 155.795000 1.955000 ;
      RECT 155.625000  3.485000 155.795000 3.655000 ;
      RECT 155.625000  5.355000 155.795000 5.525000 ;
      RECT 156.085000 -0.085000 156.255000 0.085000 ;
      RECT 156.085000  2.635000 156.255000 2.805000 ;
      RECT 156.085000  5.355000 156.255000 5.525000 ;
      RECT 156.210000  2.140000 156.380000 2.310000 ;
      RECT 156.210000  3.130000 156.380000 3.300000 ;
      RECT 156.545000 -0.085000 156.715000 0.085000 ;
      RECT 156.545000  2.635000 156.715000 2.805000 ;
      RECT 156.545000  5.355000 156.715000 5.525000 ;
      RECT 157.005000 -0.085000 157.175000 0.085000 ;
      RECT 157.005000  2.635000 157.175000 2.805000 ;
      RECT 157.005000  5.355000 157.175000 5.525000 ;
      RECT 157.465000 -0.085000 157.635000 0.085000 ;
      RECT 157.465000  2.635000 157.635000 2.805000 ;
      RECT 157.465000  5.355000 157.635000 5.525000 ;
      RECT 157.925000 -0.085000 158.095000 0.085000 ;
      RECT 157.925000  2.635000 158.095000 2.805000 ;
      RECT 157.925000  5.355000 158.095000 5.525000 ;
      RECT 158.260000  2.140000 158.430000 2.310000 ;
      RECT 158.260000  3.130000 158.430000 3.300000 ;
      RECT 158.385000 -0.085000 158.555000 0.085000 ;
      RECT 158.385000  2.635000 158.555000 2.805000 ;
      RECT 158.385000  5.355000 158.555000 5.525000 ;
      RECT 158.845000 -0.085000 159.015000 0.085000 ;
      RECT 158.845000  1.785000 159.015000 1.955000 ;
      RECT 158.845000  3.485000 159.015000 3.655000 ;
      RECT 158.845000  5.355000 159.015000 5.525000 ;
      RECT 159.255000  2.140000 159.425000 2.310000 ;
      RECT 159.255000  3.130000 159.425000 3.300000 ;
      RECT 159.305000 -0.085000 159.475000 0.085000 ;
      RECT 159.305000  2.635000 159.475000 2.805000 ;
      RECT 159.305000  5.355000 159.475000 5.525000 ;
      RECT 159.765000 -0.085000 159.935000 0.085000 ;
      RECT 159.765000  2.635000 159.935000 2.805000 ;
      RECT 159.765000  5.355000 159.935000 5.525000 ;
      RECT 160.195000  2.140000 160.365000 2.310000 ;
      RECT 160.195000  3.130000 160.365000 3.300000 ;
      RECT 160.225000 -0.085000 160.395000 0.085000 ;
      RECT 160.225000  2.635000 160.395000 2.805000 ;
      RECT 160.225000  5.355000 160.395000 5.525000 ;
      RECT 160.685000 -0.085000 160.855000 0.085000 ;
      RECT 160.685000  2.635000 160.855000 2.805000 ;
      RECT 160.685000  5.355000 160.855000 5.525000 ;
      RECT 160.715000  2.140000 160.885000 2.310000 ;
      RECT 160.715000  3.130000 160.885000 3.300000 ;
      RECT 161.145000 -0.085000 161.315000 0.085000 ;
      RECT 161.145000  2.635000 161.315000 2.805000 ;
      RECT 161.145000  5.355000 161.315000 5.525000 ;
      RECT 161.605000 -0.085000 161.775000 0.085000 ;
      RECT 161.605000  2.635000 161.775000 2.805000 ;
      RECT 161.605000  5.355000 161.775000 5.525000 ;
      RECT 161.655000  2.140000 161.825000 2.310000 ;
      RECT 161.655000  3.130000 161.825000 3.300000 ;
      RECT 162.065000 -0.085000 162.235000 0.085000 ;
      RECT 162.065000  1.785000 162.235000 1.955000 ;
      RECT 162.065000  3.485000 162.235000 3.655000 ;
      RECT 162.065000  5.355000 162.235000 5.525000 ;
      RECT 162.525000 -0.085000 162.695000 0.085000 ;
      RECT 162.525000  2.635000 162.695000 2.805000 ;
      RECT 162.525000  5.355000 162.695000 5.525000 ;
      RECT 162.650000  2.140000 162.820000 2.310000 ;
      RECT 162.650000  3.130000 162.820000 3.300000 ;
      RECT 162.985000 -0.085000 163.155000 0.085000 ;
      RECT 162.985000  2.635000 163.155000 2.805000 ;
      RECT 162.985000  5.355000 163.155000 5.525000 ;
      RECT 163.445000 -0.085000 163.615000 0.085000 ;
      RECT 163.445000  2.635000 163.615000 2.805000 ;
      RECT 163.445000  5.355000 163.615000 5.525000 ;
      RECT 163.905000 -0.085000 164.075000 0.085000 ;
      RECT 163.905000  2.635000 164.075000 2.805000 ;
      RECT 163.905000  5.355000 164.075000 5.525000 ;
      RECT 164.365000 -0.085000 164.535000 0.085000 ;
      RECT 164.365000  2.635000 164.535000 2.805000 ;
      RECT 164.365000  5.355000 164.535000 5.525000 ;
      RECT 164.700000  2.140000 164.870000 2.310000 ;
      RECT 164.700000  3.130000 164.870000 3.300000 ;
      RECT 164.825000 -0.085000 164.995000 0.085000 ;
      RECT 164.825000  2.635000 164.995000 2.805000 ;
      RECT 164.825000  5.355000 164.995000 5.525000 ;
      RECT 165.285000 -0.085000 165.455000 0.085000 ;
      RECT 165.285000  1.785000 165.455000 1.955000 ;
      RECT 165.285000  3.485000 165.455000 3.655000 ;
      RECT 165.285000  5.355000 165.455000 5.525000 ;
      RECT 165.695000  2.140000 165.865000 2.310000 ;
      RECT 165.695000  3.130000 165.865000 3.300000 ;
      RECT 165.745000 -0.085000 165.915000 0.085000 ;
      RECT 165.745000  2.635000 165.915000 2.805000 ;
      RECT 165.745000  5.355000 165.915000 5.525000 ;
      RECT 166.205000 -0.085000 166.375000 0.085000 ;
      RECT 166.205000  2.635000 166.375000 2.805000 ;
      RECT 166.205000  5.355000 166.375000 5.525000 ;
      RECT 166.635000  2.140000 166.805000 2.310000 ;
      RECT 166.635000  3.130000 166.805000 3.300000 ;
      RECT 166.665000 -0.085000 166.835000 0.085000 ;
      RECT 166.665000  2.635000 166.835000 2.805000 ;
      RECT 166.665000  5.355000 166.835000 5.525000 ;
      RECT 167.125000 -0.085000 167.295000 0.085000 ;
      RECT 167.125000  2.635000 167.295000 2.805000 ;
      RECT 167.125000  5.355000 167.295000 5.525000 ;
      RECT 167.155000  2.140000 167.325000 2.310000 ;
      RECT 167.155000  3.130000 167.325000 3.300000 ;
      RECT 167.585000 -0.085000 167.755000 0.085000 ;
      RECT 167.585000  2.635000 167.755000 2.805000 ;
      RECT 167.585000  5.355000 167.755000 5.525000 ;
      RECT 168.045000 -0.085000 168.215000 0.085000 ;
      RECT 168.045000  2.635000 168.215000 2.805000 ;
      RECT 168.045000  5.355000 168.215000 5.525000 ;
      RECT 168.095000  2.140000 168.265000 2.310000 ;
      RECT 168.095000  3.130000 168.265000 3.300000 ;
      RECT 168.505000 -0.085000 168.675000 0.085000 ;
      RECT 168.505000  1.785000 168.675000 1.955000 ;
      RECT 168.505000  3.485000 168.675000 3.655000 ;
      RECT 168.505000  5.355000 168.675000 5.525000 ;
      RECT 168.965000 -0.085000 169.135000 0.085000 ;
      RECT 168.965000  2.635000 169.135000 2.805000 ;
      RECT 168.965000  5.355000 169.135000 5.525000 ;
      RECT 169.090000  2.140000 169.260000 2.310000 ;
      RECT 169.090000  3.130000 169.260000 3.300000 ;
      RECT 169.425000 -0.085000 169.595000 0.085000 ;
      RECT 169.425000  2.635000 169.595000 2.805000 ;
      RECT 169.425000  5.355000 169.595000 5.525000 ;
      RECT 169.885000 -0.085000 170.055000 0.085000 ;
      RECT 169.885000  2.635000 170.055000 2.805000 ;
      RECT 169.885000  5.355000 170.055000 5.525000 ;
      RECT 170.345000 -0.085000 170.515000 0.085000 ;
      RECT 170.345000  2.635000 170.515000 2.805000 ;
      RECT 170.345000  5.355000 170.515000 5.525000 ;
      RECT 170.805000 -0.085000 170.975000 0.085000 ;
      RECT 170.805000  2.635000 170.975000 2.805000 ;
      RECT 170.805000  5.355000 170.975000 5.525000 ;
      RECT 171.140000  2.140000 171.310000 2.310000 ;
      RECT 171.140000  3.130000 171.310000 3.300000 ;
      RECT 171.265000 -0.085000 171.435000 0.085000 ;
      RECT 171.265000  2.635000 171.435000 2.805000 ;
      RECT 171.265000  5.355000 171.435000 5.525000 ;
      RECT 171.725000 -0.085000 171.895000 0.085000 ;
      RECT 171.725000  1.785000 171.895000 1.955000 ;
      RECT 171.725000  3.485000 171.895000 3.655000 ;
      RECT 171.725000  5.355000 171.895000 5.525000 ;
      RECT 172.135000  2.140000 172.305000 2.310000 ;
      RECT 172.135000  3.130000 172.305000 3.300000 ;
      RECT 172.185000 -0.085000 172.355000 0.085000 ;
      RECT 172.185000  2.635000 172.355000 2.805000 ;
      RECT 172.185000  5.355000 172.355000 5.525000 ;
      RECT 172.645000 -0.085000 172.815000 0.085000 ;
      RECT 172.645000  2.635000 172.815000 2.805000 ;
      RECT 172.645000  5.355000 172.815000 5.525000 ;
      RECT 173.075000  2.140000 173.245000 2.310000 ;
      RECT 173.075000  3.130000 173.245000 3.300000 ;
      RECT 173.105000 -0.085000 173.275000 0.085000 ;
      RECT 173.105000  2.635000 173.275000 2.805000 ;
      RECT 173.105000  5.355000 173.275000 5.525000 ;
      RECT 173.565000 -0.085000 173.735000 0.085000 ;
      RECT 173.565000  2.635000 173.735000 2.805000 ;
      RECT 173.565000  5.355000 173.735000 5.525000 ;
      RECT 174.025000 -0.085000 174.195000 0.085000 ;
      RECT 174.025000  2.635000 174.195000 2.805000 ;
      RECT 174.025000  5.355000 174.195000 5.525000 ;
      RECT 174.065000  2.140000 174.235000 2.310000 ;
      RECT 174.065000  3.130000 174.235000 3.300000 ;
      RECT 174.485000 -0.085000 174.655000 0.085000 ;
      RECT 174.485000  2.635000 174.655000 2.805000 ;
      RECT 174.485000  5.355000 174.655000 5.525000 ;
      RECT 174.945000 -0.085000 175.115000 0.085000 ;
      RECT 174.945000  2.635000 175.115000 2.805000 ;
      RECT 174.945000  5.355000 175.115000 5.525000 ;
      RECT 175.005000  2.140000 175.175000 2.310000 ;
      RECT 175.005000  3.130000 175.175000 3.300000 ;
      RECT 175.405000 -0.085000 175.575000 0.085000 ;
      RECT 175.405000  2.635000 175.575000 2.805000 ;
      RECT 175.405000  5.355000 175.575000 5.525000 ;
      RECT 175.865000 -0.085000 176.035000 0.085000 ;
      RECT 175.865000  2.635000 176.035000 2.805000 ;
      RECT 175.865000  5.355000 176.035000 5.525000 ;
      RECT 175.985000  2.140000 176.155000 2.310000 ;
      RECT 175.985000  3.130000 176.155000 3.300000 ;
      RECT 176.325000 -0.085000 176.495000 0.085000 ;
      RECT 176.325000  5.355000 176.495000 5.525000 ;
      RECT 176.465000  1.785000 176.635000 1.955000 ;
      RECT 176.465000  3.485000 176.635000 3.655000 ;
      RECT 176.785000 -0.085000 176.955000 0.085000 ;
      RECT 176.785000  5.355000 176.955000 5.525000 ;
      RECT 176.935000  2.140000 177.105000 2.310000 ;
      RECT 176.935000  3.130000 177.105000 3.300000 ;
      RECT 177.245000 -0.085000 177.415000 0.085000 ;
      RECT 177.245000  5.355000 177.415000 5.525000 ;
      RECT 177.405000  1.785000 177.575000 1.955000 ;
      RECT 177.405000  3.485000 177.575000 3.655000 ;
      RECT 177.705000 -0.085000 177.875000 0.085000 ;
      RECT 177.705000  5.355000 177.875000 5.525000 ;
      RECT 177.885000  2.140000 178.055000 2.310000 ;
      RECT 177.885000  3.130000 178.055000 3.300000 ;
      RECT 178.165000 -0.085000 178.335000 0.085000 ;
      RECT 178.165000  2.635000 178.335000 2.805000 ;
      RECT 178.165000  5.355000 178.335000 5.525000 ;
      RECT 178.625000 -0.085000 178.795000 0.085000 ;
      RECT 178.625000  2.635000 178.795000 2.805000 ;
      RECT 178.625000  5.355000 178.795000 5.525000 ;
      RECT 179.085000 -0.085000 179.255000 0.085000 ;
      RECT 179.085000  2.635000 179.255000 2.805000 ;
      RECT 179.085000  5.355000 179.255000 5.525000 ;
      RECT 179.545000 -0.085000 179.715000 0.085000 ;
      RECT 179.545000  2.635000 179.715000 2.805000 ;
      RECT 179.545000  5.355000 179.715000 5.525000 ;
      RECT 180.005000 -0.085000 180.175000 0.085000 ;
      RECT 180.005000  2.635000 180.175000 2.805000 ;
      RECT 180.005000  5.355000 180.175000 5.525000 ;
      RECT 180.465000 -0.085000 180.635000 0.085000 ;
      RECT 180.465000  2.635000 180.635000 2.805000 ;
      RECT 180.465000  5.355000 180.635000 5.525000 ;
      RECT 180.925000 -0.085000 181.095000 0.085000 ;
      RECT 180.925000  2.635000 181.095000 2.805000 ;
      RECT 180.925000  5.355000 181.095000 5.525000 ;
      RECT 181.385000 -0.085000 181.555000 0.085000 ;
      RECT 181.385000  2.635000 181.555000 2.805000 ;
      RECT 181.385000  5.355000 181.555000 5.525000 ;
      RECT 181.665000  2.140000 181.835000 2.310000 ;
      RECT 181.665000  3.130000 181.835000 3.300000 ;
      RECT 181.845000 -0.085000 182.015000 0.085000 ;
      RECT 181.845000  5.355000 182.015000 5.525000 ;
      RECT 182.145000  1.785000 182.315000 1.955000 ;
      RECT 182.145000  3.485000 182.315000 3.655000 ;
      RECT 182.305000 -0.085000 182.475000 0.085000 ;
      RECT 182.305000  5.355000 182.475000 5.525000 ;
      RECT 182.615000  2.140000 182.785000 2.310000 ;
      RECT 182.615000  3.130000 182.785000 3.300000 ;
      RECT 182.765000 -0.085000 182.935000 0.085000 ;
      RECT 182.765000  5.355000 182.935000 5.525000 ;
      RECT 183.085000  1.785000 183.255000 1.955000 ;
      RECT 183.085000  3.485000 183.255000 3.655000 ;
      RECT 183.225000 -0.085000 183.395000 0.085000 ;
      RECT 183.225000  5.355000 183.395000 5.525000 ;
      RECT 183.565000  2.140000 183.735000 2.310000 ;
      RECT 183.565000  3.130000 183.735000 3.300000 ;
      RECT 183.685000 -0.085000 183.855000 0.085000 ;
      RECT 183.685000  2.635000 183.855000 2.805000 ;
      RECT 183.685000  5.355000 183.855000 5.525000 ;
      RECT 184.145000 -0.085000 184.315000 0.085000 ;
      RECT 184.145000  2.635000 184.315000 2.805000 ;
      RECT 184.145000  5.355000 184.315000 5.525000 ;
      RECT 184.545000  2.140000 184.715000 2.310000 ;
      RECT 184.545000  3.130000 184.715000 3.300000 ;
      RECT 184.605000 -0.085000 184.775000 0.085000 ;
      RECT 184.605000  2.635000 184.775000 2.805000 ;
      RECT 184.605000  5.355000 184.775000 5.525000 ;
      RECT 185.065000 -0.085000 185.235000 0.085000 ;
      RECT 185.065000  2.635000 185.235000 2.805000 ;
      RECT 185.065000  5.355000 185.235000 5.525000 ;
      RECT 185.485000  2.140000 185.655000 2.310000 ;
      RECT 185.485000  3.130000 185.655000 3.300000 ;
      RECT 185.525000 -0.085000 185.695000 0.085000 ;
      RECT 185.525000  2.635000 185.695000 2.805000 ;
      RECT 185.525000  5.355000 185.695000 5.525000 ;
      RECT 185.985000 -0.085000 186.155000 0.085000 ;
      RECT 185.985000  2.635000 186.155000 2.805000 ;
      RECT 185.985000  5.355000 186.155000 5.525000 ;
      RECT 186.445000 -0.085000 186.615000 0.085000 ;
      RECT 186.445000  2.635000 186.615000 2.805000 ;
      RECT 186.445000  5.355000 186.615000 5.525000 ;
      RECT 186.905000 -0.085000 187.075000 0.085000 ;
      RECT 186.905000  2.635000 187.075000 2.805000 ;
      RECT 186.905000  5.355000 187.075000 5.525000 ;
      RECT 186.945000  2.140000 187.115000 2.310000 ;
      RECT 186.945000  3.130000 187.115000 3.300000 ;
      RECT 187.365000 -0.085000 187.535000 0.085000 ;
      RECT 187.365000  2.635000 187.535000 2.805000 ;
      RECT 187.365000  5.355000 187.535000 5.525000 ;
      RECT 187.825000 -0.085000 187.995000 0.085000 ;
      RECT 187.825000  2.635000 187.995000 2.805000 ;
      RECT 187.825000  5.355000 187.995000 5.525000 ;
      RECT 187.885000  2.140000 188.055000 2.310000 ;
      RECT 187.885000  3.130000 188.055000 3.300000 ;
      RECT 188.285000 -0.085000 188.455000 0.085000 ;
      RECT 188.285000  2.635000 188.455000 2.805000 ;
      RECT 188.285000  5.355000 188.455000 5.525000 ;
      RECT 188.745000 -0.085000 188.915000 0.085000 ;
      RECT 188.745000  2.635000 188.915000 2.805000 ;
      RECT 188.745000  5.355000 188.915000 5.525000 ;
      RECT 188.865000  2.140000 189.035000 2.310000 ;
      RECT 188.865000  3.130000 189.035000 3.300000 ;
      RECT 189.205000 -0.085000 189.375000 0.085000 ;
      RECT 189.205000  5.355000 189.375000 5.525000 ;
      RECT 189.345000  1.785000 189.515000 1.955000 ;
      RECT 189.345000  3.485000 189.515000 3.655000 ;
      RECT 189.665000 -0.085000 189.835000 0.085000 ;
      RECT 189.665000  5.355000 189.835000 5.525000 ;
      RECT 189.815000  2.140000 189.985000 2.310000 ;
      RECT 189.815000  3.130000 189.985000 3.300000 ;
      RECT 190.125000 -0.085000 190.295000 0.085000 ;
      RECT 190.125000  5.355000 190.295000 5.525000 ;
      RECT 190.285000  1.785000 190.455000 1.955000 ;
      RECT 190.285000  3.485000 190.455000 3.655000 ;
      RECT 190.585000 -0.085000 190.755000 0.085000 ;
      RECT 190.585000  5.355000 190.755000 5.525000 ;
      RECT 190.765000  2.140000 190.935000 2.310000 ;
      RECT 190.765000  3.130000 190.935000 3.300000 ;
      RECT 191.045000 -0.085000 191.215000 0.085000 ;
      RECT 191.045000  2.635000 191.215000 2.805000 ;
      RECT 191.045000  5.355000 191.215000 5.525000 ;
      RECT 191.505000 -0.085000 191.675000 0.085000 ;
      RECT 191.505000  2.635000 191.675000 2.805000 ;
      RECT 191.505000  5.355000 191.675000 5.525000 ;
      RECT 191.965000 -0.085000 192.135000 0.085000 ;
      RECT 191.965000  2.635000 192.135000 2.805000 ;
      RECT 191.965000  5.355000 192.135000 5.525000 ;
      RECT 192.425000 -0.085000 192.595000 0.085000 ;
      RECT 192.425000  2.635000 192.595000 2.805000 ;
      RECT 192.425000  5.355000 192.595000 5.525000 ;
      RECT 192.885000 -0.085000 193.055000 0.085000 ;
      RECT 192.885000  2.635000 193.055000 2.805000 ;
      RECT 192.885000  5.355000 193.055000 5.525000 ;
      RECT 193.345000 -0.085000 193.515000 0.085000 ;
      RECT 193.345000  2.635000 193.515000 2.805000 ;
      RECT 193.345000  5.355000 193.515000 5.525000 ;
      RECT 193.805000 -0.085000 193.975000 0.085000 ;
      RECT 193.805000  2.635000 193.975000 2.805000 ;
      RECT 193.805000  5.355000 193.975000 5.525000 ;
      RECT 194.265000 -0.085000 194.435000 0.085000 ;
      RECT 194.265000  2.635000 194.435000 2.805000 ;
      RECT 194.265000  5.355000 194.435000 5.525000 ;
      RECT 194.545000  2.140000 194.715000 2.310000 ;
      RECT 194.545000  3.130000 194.715000 3.300000 ;
      RECT 194.725000 -0.085000 194.895000 0.085000 ;
      RECT 194.725000  5.355000 194.895000 5.525000 ;
      RECT 195.025000  1.785000 195.195000 1.955000 ;
      RECT 195.025000  3.485000 195.195000 3.655000 ;
      RECT 195.185000 -0.085000 195.355000 0.085000 ;
      RECT 195.185000  5.355000 195.355000 5.525000 ;
      RECT 195.495000  2.140000 195.665000 2.310000 ;
      RECT 195.495000  3.130000 195.665000 3.300000 ;
      RECT 195.645000 -0.085000 195.815000 0.085000 ;
      RECT 195.645000  5.355000 195.815000 5.525000 ;
      RECT 195.965000  1.785000 196.135000 1.955000 ;
      RECT 195.965000  3.485000 196.135000 3.655000 ;
      RECT 196.105000 -0.085000 196.275000 0.085000 ;
      RECT 196.105000  5.355000 196.275000 5.525000 ;
      RECT 196.445000  2.140000 196.615000 2.310000 ;
      RECT 196.445000  3.130000 196.615000 3.300000 ;
      RECT 196.565000 -0.085000 196.735000 0.085000 ;
      RECT 196.565000  2.635000 196.735000 2.805000 ;
      RECT 196.565000  5.355000 196.735000 5.525000 ;
      RECT 197.025000 -0.085000 197.195000 0.085000 ;
      RECT 197.025000  2.635000 197.195000 2.805000 ;
      RECT 197.025000  5.355000 197.195000 5.525000 ;
      RECT 197.425000  2.140000 197.595000 2.310000 ;
      RECT 197.425000  3.130000 197.595000 3.300000 ;
      RECT 197.485000 -0.085000 197.655000 0.085000 ;
      RECT 197.485000  2.635000 197.655000 2.805000 ;
      RECT 197.485000  5.355000 197.655000 5.525000 ;
      RECT 197.945000 -0.085000 198.115000 0.085000 ;
      RECT 197.945000  2.635000 198.115000 2.805000 ;
      RECT 197.945000  5.355000 198.115000 5.525000 ;
      RECT 198.365000  2.140000 198.535000 2.310000 ;
      RECT 198.365000  3.130000 198.535000 3.300000 ;
      RECT 198.405000 -0.085000 198.575000 0.085000 ;
      RECT 198.405000  2.635000 198.575000 2.805000 ;
      RECT 198.405000  5.355000 198.575000 5.525000 ;
      RECT 198.865000 -0.085000 199.035000 0.085000 ;
      RECT 198.865000  2.635000 199.035000 2.805000 ;
      RECT 198.865000  5.355000 199.035000 5.525000 ;
      RECT 199.325000 -0.085000 199.495000 0.085000 ;
      RECT 199.325000  2.635000 199.495000 2.805000 ;
      RECT 199.325000  5.355000 199.495000 5.525000 ;
      RECT 199.785000 -0.085000 199.955000 0.085000 ;
      RECT 199.785000  2.635000 199.955000 2.805000 ;
      RECT 199.785000  5.355000 199.955000 5.525000 ;
      RECT 200.245000 -0.085000 200.415000 0.085000 ;
      RECT 200.245000  2.635000 200.415000 2.805000 ;
      RECT 200.245000  5.355000 200.415000 5.525000 ;
      RECT 200.285000  2.140000 200.455000 2.310000 ;
      RECT 200.285000  3.130000 200.455000 3.300000 ;
      RECT 200.705000 -0.085000 200.875000 0.085000 ;
      RECT 200.705000  2.635000 200.875000 2.805000 ;
      RECT 200.705000  5.355000 200.875000 5.525000 ;
      RECT 201.165000 -0.085000 201.335000 0.085000 ;
      RECT 201.165000  2.635000 201.335000 2.805000 ;
      RECT 201.165000  5.355000 201.335000 5.525000 ;
      RECT 201.225000  2.140000 201.395000 2.310000 ;
      RECT 201.225000  3.130000 201.395000 3.300000 ;
      RECT 201.625000 -0.085000 201.795000 0.085000 ;
      RECT 201.625000  2.635000 201.795000 2.805000 ;
      RECT 201.625000  5.355000 201.795000 5.525000 ;
      RECT 202.085000 -0.085000 202.255000 0.085000 ;
      RECT 202.085000  2.635000 202.255000 2.805000 ;
      RECT 202.085000  5.355000 202.255000 5.525000 ;
      RECT 202.205000  2.140000 202.375000 2.310000 ;
      RECT 202.205000  3.130000 202.375000 3.300000 ;
      RECT 202.545000 -0.085000 202.715000 0.085000 ;
      RECT 202.545000  5.355000 202.715000 5.525000 ;
      RECT 202.685000  1.785000 202.855000 1.955000 ;
      RECT 202.685000  3.485000 202.855000 3.655000 ;
      RECT 203.005000 -0.085000 203.175000 0.085000 ;
      RECT 203.005000  5.355000 203.175000 5.525000 ;
      RECT 203.155000  2.140000 203.325000 2.310000 ;
      RECT 203.155000  3.130000 203.325000 3.300000 ;
      RECT 203.465000 -0.085000 203.635000 0.085000 ;
      RECT 203.465000  5.355000 203.635000 5.525000 ;
      RECT 203.625000  1.785000 203.795000 1.955000 ;
      RECT 203.625000  3.485000 203.795000 3.655000 ;
      RECT 203.925000 -0.085000 204.095000 0.085000 ;
      RECT 203.925000  5.355000 204.095000 5.525000 ;
      RECT 204.105000  2.140000 204.275000 2.310000 ;
      RECT 204.105000  3.130000 204.275000 3.300000 ;
      RECT 204.385000 -0.085000 204.555000 0.085000 ;
      RECT 204.385000  2.635000 204.555000 2.805000 ;
      RECT 204.385000  5.355000 204.555000 5.525000 ;
      RECT 204.845000 -0.085000 205.015000 0.085000 ;
      RECT 204.845000  2.635000 205.015000 2.805000 ;
      RECT 204.845000  5.355000 205.015000 5.525000 ;
      RECT 205.305000 -0.085000 205.475000 0.085000 ;
      RECT 205.305000  2.635000 205.475000 2.805000 ;
      RECT 205.305000  5.355000 205.475000 5.525000 ;
      RECT 205.765000 -0.085000 205.935000 0.085000 ;
      RECT 205.765000  2.635000 205.935000 2.805000 ;
      RECT 205.765000  5.355000 205.935000 5.525000 ;
      RECT 206.225000 -0.085000 206.395000 0.085000 ;
      RECT 206.225000  2.635000 206.395000 2.805000 ;
      RECT 206.225000  5.355000 206.395000 5.525000 ;
      RECT 206.685000 -0.085000 206.855000 0.085000 ;
      RECT 206.685000  2.635000 206.855000 2.805000 ;
      RECT 206.685000  5.355000 206.855000 5.525000 ;
      RECT 207.145000 -0.085000 207.315000 0.085000 ;
      RECT 207.145000  2.635000 207.315000 2.805000 ;
      RECT 207.145000  5.355000 207.315000 5.525000 ;
      RECT 207.605000 -0.085000 207.775000 0.085000 ;
      RECT 207.605000  2.635000 207.775000 2.805000 ;
      RECT 207.605000  5.355000 207.775000 5.525000 ;
      RECT 207.885000  2.140000 208.055000 2.310000 ;
      RECT 207.885000  3.130000 208.055000 3.300000 ;
      RECT 208.065000 -0.085000 208.235000 0.085000 ;
      RECT 208.065000  5.355000 208.235000 5.525000 ;
      RECT 208.365000  1.785000 208.535000 1.955000 ;
      RECT 208.365000  3.485000 208.535000 3.655000 ;
      RECT 208.525000 -0.085000 208.695000 0.085000 ;
      RECT 208.525000  5.355000 208.695000 5.525000 ;
      RECT 208.835000  2.140000 209.005000 2.310000 ;
      RECT 208.835000  3.130000 209.005000 3.300000 ;
      RECT 208.985000 -0.085000 209.155000 0.085000 ;
      RECT 208.985000  5.355000 209.155000 5.525000 ;
      RECT 209.305000  1.785000 209.475000 1.955000 ;
      RECT 209.305000  3.485000 209.475000 3.655000 ;
      RECT 209.445000 -0.085000 209.615000 0.085000 ;
      RECT 209.445000  5.355000 209.615000 5.525000 ;
      RECT 209.785000  2.140000 209.955000 2.310000 ;
      RECT 209.785000  3.130000 209.955000 3.300000 ;
      RECT 209.905000 -0.085000 210.075000 0.085000 ;
      RECT 209.905000  2.635000 210.075000 2.805000 ;
      RECT 209.905000  5.355000 210.075000 5.525000 ;
      RECT 210.365000 -0.085000 210.535000 0.085000 ;
      RECT 210.365000  2.635000 210.535000 2.805000 ;
      RECT 210.365000  5.355000 210.535000 5.525000 ;
      RECT 210.765000  2.140000 210.935000 2.310000 ;
      RECT 210.765000  3.130000 210.935000 3.300000 ;
      RECT 210.825000 -0.085000 210.995000 0.085000 ;
      RECT 210.825000  2.635000 210.995000 2.805000 ;
      RECT 210.825000  5.355000 210.995000 5.525000 ;
      RECT 211.285000 -0.085000 211.455000 0.085000 ;
      RECT 211.285000  2.635000 211.455000 2.805000 ;
      RECT 211.285000  5.355000 211.455000 5.525000 ;
      RECT 211.705000  2.140000 211.875000 2.310000 ;
      RECT 211.705000  3.130000 211.875000 3.300000 ;
      RECT 211.745000 -0.085000 211.915000 0.085000 ;
      RECT 211.745000  2.635000 211.915000 2.805000 ;
      RECT 211.745000  5.355000 211.915000 5.525000 ;
      RECT 212.205000 -0.085000 212.375000 0.085000 ;
      RECT 212.205000  2.635000 212.375000 2.805000 ;
      RECT 212.205000  5.355000 212.375000 5.525000 ;
      RECT 212.665000 -0.085000 212.835000 0.085000 ;
      RECT 212.665000  2.635000 212.835000 2.805000 ;
      RECT 212.665000  5.355000 212.835000 5.525000 ;
      RECT 213.125000 -0.085000 213.295000 0.085000 ;
      RECT 213.125000  2.635000 213.295000 2.805000 ;
      RECT 213.125000  5.355000 213.295000 5.525000 ;
      RECT 213.165000  2.140000 213.335000 2.310000 ;
      RECT 213.165000  3.130000 213.335000 3.300000 ;
      RECT 213.585000 -0.085000 213.755000 0.085000 ;
      RECT 213.585000  2.635000 213.755000 2.805000 ;
      RECT 213.585000  5.355000 213.755000 5.525000 ;
      RECT 214.045000 -0.085000 214.215000 0.085000 ;
      RECT 214.045000  2.635000 214.215000 2.805000 ;
      RECT 214.045000  5.355000 214.215000 5.525000 ;
      RECT 214.105000  2.140000 214.275000 2.310000 ;
      RECT 214.105000  3.130000 214.275000 3.300000 ;
      RECT 214.505000 -0.085000 214.675000 0.085000 ;
      RECT 214.505000  2.635000 214.675000 2.805000 ;
      RECT 214.505000  5.355000 214.675000 5.525000 ;
      RECT 214.965000 -0.085000 215.135000 0.085000 ;
      RECT 214.965000  2.635000 215.135000 2.805000 ;
      RECT 214.965000  5.355000 215.135000 5.525000 ;
      RECT 215.085000  2.140000 215.255000 2.310000 ;
      RECT 215.085000  3.130000 215.255000 3.300000 ;
      RECT 215.425000 -0.085000 215.595000 0.085000 ;
      RECT 215.425000  5.355000 215.595000 5.525000 ;
      RECT 215.565000  1.785000 215.735000 1.955000 ;
      RECT 215.565000  3.485000 215.735000 3.655000 ;
      RECT 215.885000 -0.085000 216.055000 0.085000 ;
      RECT 215.885000  5.355000 216.055000 5.525000 ;
      RECT 216.035000  2.140000 216.205000 2.310000 ;
      RECT 216.035000  3.130000 216.205000 3.300000 ;
      RECT 216.345000 -0.085000 216.515000 0.085000 ;
      RECT 216.345000  5.355000 216.515000 5.525000 ;
      RECT 216.505000  1.785000 216.675000 1.955000 ;
      RECT 216.505000  3.485000 216.675000 3.655000 ;
      RECT 216.805000 -0.085000 216.975000 0.085000 ;
      RECT 216.805000  5.355000 216.975000 5.525000 ;
      RECT 216.985000  2.140000 217.155000 2.310000 ;
      RECT 216.985000  3.130000 217.155000 3.300000 ;
      RECT 217.265000 -0.085000 217.435000 0.085000 ;
      RECT 217.265000  2.635000 217.435000 2.805000 ;
      RECT 217.265000  5.355000 217.435000 5.525000 ;
      RECT 217.725000 -0.085000 217.895000 0.085000 ;
      RECT 217.725000  2.635000 217.895000 2.805000 ;
      RECT 217.725000  5.355000 217.895000 5.525000 ;
      RECT 218.185000 -0.085000 218.355000 0.085000 ;
      RECT 218.185000  2.635000 218.355000 2.805000 ;
      RECT 218.185000  5.355000 218.355000 5.525000 ;
      RECT 218.645000 -0.085000 218.815000 0.085000 ;
      RECT 218.645000  2.635000 218.815000 2.805000 ;
      RECT 218.645000  5.355000 218.815000 5.525000 ;
      RECT 219.105000 -0.085000 219.275000 0.085000 ;
      RECT 219.105000  2.635000 219.275000 2.805000 ;
      RECT 219.105000  5.355000 219.275000 5.525000 ;
      RECT 219.565000 -0.085000 219.735000 0.085000 ;
      RECT 219.565000  2.635000 219.735000 2.805000 ;
      RECT 219.565000  5.355000 219.735000 5.525000 ;
      RECT 220.025000 -0.085000 220.195000 0.085000 ;
      RECT 220.025000  2.635000 220.195000 2.805000 ;
      RECT 220.025000  5.355000 220.195000 5.525000 ;
      RECT 220.485000 -0.085000 220.655000 0.085000 ;
      RECT 220.485000  2.635000 220.655000 2.805000 ;
      RECT 220.485000  5.355000 220.655000 5.525000 ;
      RECT 220.765000  2.140000 220.935000 2.310000 ;
      RECT 220.765000  3.130000 220.935000 3.300000 ;
      RECT 220.945000 -0.085000 221.115000 0.085000 ;
      RECT 220.945000  5.355000 221.115000 5.525000 ;
      RECT 221.245000  1.785000 221.415000 1.955000 ;
      RECT 221.245000  3.485000 221.415000 3.655000 ;
      RECT 221.405000 -0.085000 221.575000 0.085000 ;
      RECT 221.405000  5.355000 221.575000 5.525000 ;
      RECT 221.715000  2.140000 221.885000 2.310000 ;
      RECT 221.715000  3.130000 221.885000 3.300000 ;
      RECT 221.865000 -0.085000 222.035000 0.085000 ;
      RECT 221.865000  5.355000 222.035000 5.525000 ;
      RECT 222.185000  1.785000 222.355000 1.955000 ;
      RECT 222.185000  3.485000 222.355000 3.655000 ;
      RECT 222.325000 -0.085000 222.495000 0.085000 ;
      RECT 222.325000  5.355000 222.495000 5.525000 ;
      RECT 222.665000  2.140000 222.835000 2.310000 ;
      RECT 222.665000  3.130000 222.835000 3.300000 ;
      RECT 222.785000 -0.085000 222.955000 0.085000 ;
      RECT 222.785000  2.635000 222.955000 2.805000 ;
      RECT 222.785000  5.355000 222.955000 5.525000 ;
      RECT 223.245000 -0.085000 223.415000 0.085000 ;
      RECT 223.245000  2.635000 223.415000 2.805000 ;
      RECT 223.245000  5.355000 223.415000 5.525000 ;
      RECT 223.645000  2.140000 223.815000 2.310000 ;
      RECT 223.645000  3.130000 223.815000 3.300000 ;
      RECT 223.705000 -0.085000 223.875000 0.085000 ;
      RECT 223.705000  2.635000 223.875000 2.805000 ;
      RECT 223.705000  5.355000 223.875000 5.525000 ;
      RECT 224.165000 -0.085000 224.335000 0.085000 ;
      RECT 224.165000  2.635000 224.335000 2.805000 ;
      RECT 224.165000  5.355000 224.335000 5.525000 ;
      RECT 224.585000  2.140000 224.755000 2.310000 ;
      RECT 224.585000  3.130000 224.755000 3.300000 ;
      RECT 224.625000 -0.085000 224.795000 0.085000 ;
      RECT 224.625000  2.635000 224.795000 2.805000 ;
      RECT 224.625000  5.355000 224.795000 5.525000 ;
      RECT 225.085000 -0.085000 225.255000 0.085000 ;
      RECT 225.085000  2.635000 225.255000 2.805000 ;
      RECT 225.085000  5.355000 225.255000 5.525000 ;
    LAYER met1 ;
      RECT   0.000000 -0.240000 225.400000 0.240000 ;
      RECT   0.000000  2.480000 225.400000 2.960000 ;
      RECT  16.645000  1.755000  16.935000 1.800000 ;
      RECT  16.645000  1.800000  23.375000 1.940000 ;
      RECT  16.645000  1.940000  16.935000 1.985000 ;
      RECT  18.945000  1.755000  19.235000 1.800000 ;
      RECT  18.945000  1.940000  19.235000 1.985000 ;
      RECT  20.785000  1.755000  21.075000 1.800000 ;
      RECT  20.785000  1.940000  21.075000 1.985000 ;
      RECT  23.085000  1.755000  23.375000 1.800000 ;
      RECT  23.085000  1.940000  23.375000 1.985000 ;
      RECT  25.845000  1.755000  26.135000 1.800000 ;
      RECT  25.845000  1.800000  35.795000 1.940000 ;
      RECT  25.845000  1.940000  26.135000 1.985000 ;
      RECT  29.065000  1.755000  29.355000 1.800000 ;
      RECT  29.065000  1.940000  29.355000 1.985000 ;
      RECT  32.285000  1.755000  32.575000 1.800000 ;
      RECT  32.285000  1.940000  32.575000 1.985000 ;
      RECT  35.505000  1.755000  35.795000 1.800000 ;
      RECT  35.505000  1.940000  35.795000 1.985000 ;
      RECT  40.245000  1.755000  40.535000 1.800000 ;
      RECT  40.245000  1.800000  60.035000 1.940000 ;
      RECT  40.245000  1.940000  40.535000 1.985000 ;
      RECT  41.185000  1.755000  41.475000 1.800000 ;
      RECT  41.185000  1.940000  41.475000 1.985000 ;
      RECT  45.925000  1.755000  46.215000 1.800000 ;
      RECT  45.925000  1.940000  46.215000 1.985000 ;
      RECT  46.865000  1.755000  47.155000 1.800000 ;
      RECT  46.865000  1.940000  47.155000 1.985000 ;
      RECT  53.125000  1.755000  53.415000 1.800000 ;
      RECT  53.125000  1.940000  53.415000 1.985000 ;
      RECT  54.065000  1.755000  54.355000 1.800000 ;
      RECT  54.065000  1.940000  54.355000 1.985000 ;
      RECT  58.805000  1.755000  59.095000 1.800000 ;
      RECT  58.805000  1.940000  59.095000 1.985000 ;
      RECT  59.745000  1.755000  60.035000 1.800000 ;
      RECT  59.745000  1.940000  60.035000 1.985000 ;
      RECT  64.025000  1.755000  64.315000 1.800000 ;
      RECT  64.025000  1.800000  79.035000 1.940000 ;
      RECT  64.025000  1.940000  64.315000 1.985000 ;
      RECT  66.325000  1.755000  66.615000 1.800000 ;
      RECT  66.325000  1.940000  66.615000 1.985000 ;
      RECT  68.165000  1.755000  68.455000 1.800000 ;
      RECT  68.165000  1.940000  68.455000 1.985000 ;
      RECT  70.465000  1.755000  70.755000 1.800000 ;
      RECT  70.465000  1.940000  70.755000 1.985000 ;
      RECT  72.305000  1.755000  72.595000 1.800000 ;
      RECT  72.305000  1.940000  72.595000 1.985000 ;
      RECT  74.605000  1.755000  74.895000 1.800000 ;
      RECT  74.605000  1.940000  74.895000 1.985000 ;
      RECT  76.445000  1.755000  76.735000 1.800000 ;
      RECT  76.445000  1.940000  76.735000 1.985000 ;
      RECT  78.745000  1.755000  79.035000 1.800000 ;
      RECT  78.745000  1.940000  79.035000 1.985000 ;
      RECT  81.505000  1.755000  81.795000 1.800000 ;
      RECT  81.505000  1.800000 104.335000 1.940000 ;
      RECT  81.505000  1.940000  81.795000 1.985000 ;
      RECT  84.725000  1.755000  85.015000 1.800000 ;
      RECT  84.725000  1.940000  85.015000 1.985000 ;
      RECT  87.945000  1.755000  88.235000 1.800000 ;
      RECT  87.945000  1.940000  88.235000 1.985000 ;
      RECT  91.165000  1.755000  91.455000 1.800000 ;
      RECT  91.165000  1.940000  91.455000 1.985000 ;
      RECT  94.385000  1.755000  94.675000 1.800000 ;
      RECT  94.385000  1.940000  94.675000 1.985000 ;
      RECT  97.605000  1.755000  97.895000 1.800000 ;
      RECT  97.605000  1.940000  97.895000 1.985000 ;
      RECT 100.825000  1.755000 101.115000 1.800000 ;
      RECT 100.825000  1.940000 101.115000 1.985000 ;
      RECT 104.045000  1.755000 104.335000 1.800000 ;
      RECT 104.045000  1.940000 104.335000 1.985000 ;
      RECT 105.800000  5.200000 225.400000 5.680000 ;
      RECT 107.545000  2.110000 107.835000 2.155000 ;
      RECT 107.545000  2.155000 111.655000 2.295000 ;
      RECT 107.545000  2.295000 107.835000 2.340000 ;
      RECT 107.545000  3.100000 107.835000 3.145000 ;
      RECT 107.545000  3.145000 111.655000 3.285000 ;
      RECT 107.545000  3.285000 107.835000 3.330000 ;
      RECT 108.025000  1.755000 108.315000 1.800000 ;
      RECT 108.025000  1.800000 128.415000 1.940000 ;
      RECT 108.025000  1.940000 108.315000 1.985000 ;
      RECT 108.025000  3.455000 108.315000 3.500000 ;
      RECT 108.025000  3.500000 128.415000 3.640000 ;
      RECT 108.025000  3.640000 108.315000 3.685000 ;
      RECT 108.495000  2.110000 108.785000 2.155000 ;
      RECT 108.495000  2.295000 108.785000 2.340000 ;
      RECT 108.495000  3.100000 108.785000 3.145000 ;
      RECT 108.495000  3.285000 108.785000 3.330000 ;
      RECT 108.965000  1.755000 109.255000 1.800000 ;
      RECT 108.965000  1.940000 109.255000 1.985000 ;
      RECT 108.965000  3.455000 109.255000 3.500000 ;
      RECT 108.965000  3.640000 109.255000 3.685000 ;
      RECT 109.445000  2.110000 109.735000 2.155000 ;
      RECT 109.445000  2.295000 109.735000 2.340000 ;
      RECT 109.445000  3.100000 109.735000 3.145000 ;
      RECT 109.445000  3.285000 109.735000 3.330000 ;
      RECT 110.425000  2.110000 110.715000 2.155000 ;
      RECT 110.425000  2.295000 110.715000 2.340000 ;
      RECT 110.425000  3.100000 110.715000 3.145000 ;
      RECT 110.425000  3.285000 110.715000 3.330000 ;
      RECT 111.365000  2.110000 111.655000 2.155000 ;
      RECT 111.365000  2.295000 111.655000 2.340000 ;
      RECT 111.365000  3.100000 111.655000 3.145000 ;
      RECT 111.365000  3.285000 111.655000 3.330000 ;
      RECT 112.365000  2.110000 112.655000 2.155000 ;
      RECT 112.365000  2.155000 116.475000 2.295000 ;
      RECT 112.365000  2.295000 112.655000 2.340000 ;
      RECT 112.365000  3.100000 112.655000 3.145000 ;
      RECT 112.365000  3.145000 116.475000 3.285000 ;
      RECT 112.365000  3.285000 112.655000 3.330000 ;
      RECT 113.305000  2.110000 113.595000 2.155000 ;
      RECT 113.305000  2.295000 113.595000 2.340000 ;
      RECT 113.305000  3.100000 113.595000 3.145000 ;
      RECT 113.305000  3.285000 113.595000 3.330000 ;
      RECT 114.285000  2.110000 114.575000 2.155000 ;
      RECT 114.285000  2.295000 114.575000 2.340000 ;
      RECT 114.285000  3.100000 114.575000 3.145000 ;
      RECT 114.285000  3.285000 114.575000 3.330000 ;
      RECT 114.765000  1.755000 115.055000 1.800000 ;
      RECT 114.765000  1.940000 115.055000 1.985000 ;
      RECT 114.765000  3.455000 115.055000 3.500000 ;
      RECT 114.765000  3.640000 115.055000 3.685000 ;
      RECT 115.235000  2.110000 115.525000 2.155000 ;
      RECT 115.235000  2.295000 115.525000 2.340000 ;
      RECT 115.235000  3.100000 115.525000 3.145000 ;
      RECT 115.235000  3.285000 115.525000 3.330000 ;
      RECT 115.705000  1.755000 115.995000 1.800000 ;
      RECT 115.705000  1.940000 115.995000 1.985000 ;
      RECT 115.705000  3.455000 115.995000 3.500000 ;
      RECT 115.705000  3.640000 115.995000 3.685000 ;
      RECT 116.185000  2.110000 116.475000 2.155000 ;
      RECT 116.185000  2.295000 116.475000 2.340000 ;
      RECT 116.185000  3.100000 116.475000 3.145000 ;
      RECT 116.185000  3.285000 116.475000 3.330000 ;
      RECT 119.965000  2.110000 120.255000 2.155000 ;
      RECT 119.965000  2.155000 124.075000 2.295000 ;
      RECT 119.965000  2.295000 120.255000 2.340000 ;
      RECT 119.965000  3.100000 120.255000 3.145000 ;
      RECT 119.965000  3.145000 124.075000 3.285000 ;
      RECT 119.965000  3.285000 120.255000 3.330000 ;
      RECT 120.445000  1.755000 120.735000 1.800000 ;
      RECT 120.445000  1.940000 120.735000 1.985000 ;
      RECT 120.445000  3.455000 120.735000 3.500000 ;
      RECT 120.445000  3.640000 120.735000 3.685000 ;
      RECT 120.915000  2.110000 121.205000 2.155000 ;
      RECT 120.915000  2.295000 121.205000 2.340000 ;
      RECT 120.915000  3.100000 121.205000 3.145000 ;
      RECT 120.915000  3.285000 121.205000 3.330000 ;
      RECT 121.385000  1.755000 121.675000 1.800000 ;
      RECT 121.385000  1.940000 121.675000 1.985000 ;
      RECT 121.385000  3.455000 121.675000 3.500000 ;
      RECT 121.385000  3.640000 121.675000 3.685000 ;
      RECT 121.865000  2.110000 122.155000 2.155000 ;
      RECT 121.865000  2.295000 122.155000 2.340000 ;
      RECT 121.865000  3.100000 122.155000 3.145000 ;
      RECT 121.865000  3.285000 122.155000 3.330000 ;
      RECT 122.845000  2.110000 123.135000 2.155000 ;
      RECT 122.845000  2.295000 123.135000 2.340000 ;
      RECT 122.845000  3.100000 123.135000 3.145000 ;
      RECT 122.845000  3.285000 123.135000 3.330000 ;
      RECT 123.785000  2.110000 124.075000 2.155000 ;
      RECT 123.785000  2.295000 124.075000 2.340000 ;
      RECT 123.785000  3.100000 124.075000 3.145000 ;
      RECT 123.785000  3.285000 124.075000 3.330000 ;
      RECT 124.785000  2.110000 125.075000 2.155000 ;
      RECT 124.785000  2.155000 128.895000 2.295000 ;
      RECT 124.785000  2.295000 125.075000 2.340000 ;
      RECT 124.785000  3.100000 125.075000 3.145000 ;
      RECT 124.785000  3.145000 128.895000 3.285000 ;
      RECT 124.785000  3.285000 125.075000 3.330000 ;
      RECT 125.725000  2.110000 126.015000 2.155000 ;
      RECT 125.725000  2.295000 126.015000 2.340000 ;
      RECT 125.725000  3.100000 126.015000 3.145000 ;
      RECT 125.725000  3.285000 126.015000 3.330000 ;
      RECT 126.705000  2.110000 126.995000 2.155000 ;
      RECT 126.705000  2.295000 126.995000 2.340000 ;
      RECT 126.705000  3.100000 126.995000 3.145000 ;
      RECT 126.705000  3.285000 126.995000 3.330000 ;
      RECT 127.185000  1.755000 127.475000 1.800000 ;
      RECT 127.185000  1.940000 127.475000 1.985000 ;
      RECT 127.185000  3.455000 127.475000 3.500000 ;
      RECT 127.185000  3.640000 127.475000 3.685000 ;
      RECT 127.655000  2.110000 127.945000 2.155000 ;
      RECT 127.655000  2.295000 127.945000 2.340000 ;
      RECT 127.655000  3.100000 127.945000 3.145000 ;
      RECT 127.655000  3.285000 127.945000 3.330000 ;
      RECT 128.125000  1.755000 128.415000 1.800000 ;
      RECT 128.125000  1.940000 128.415000 1.985000 ;
      RECT 128.125000  3.455000 128.415000 3.500000 ;
      RECT 128.125000  3.640000 128.415000 3.685000 ;
      RECT 128.605000  2.110000 128.895000 2.155000 ;
      RECT 128.605000  2.295000 128.895000 2.340000 ;
      RECT 128.605000  3.100000 128.895000 3.145000 ;
      RECT 128.605000  3.285000 128.895000 3.330000 ;
      RECT 131.645000  1.755000 131.935000 1.800000 ;
      RECT 131.645000  1.800000 146.655000 1.940000 ;
      RECT 131.645000  1.940000 131.935000 1.985000 ;
      RECT 131.645000  3.455000 131.935000 3.500000 ;
      RECT 131.645000  3.500000 146.655000 3.640000 ;
      RECT 131.645000  3.640000 131.935000 3.685000 ;
      RECT 133.945000  1.755000 134.235000 1.800000 ;
      RECT 133.945000  1.940000 134.235000 1.985000 ;
      RECT 133.945000  3.455000 134.235000 3.500000 ;
      RECT 133.945000  3.640000 134.235000 3.685000 ;
      RECT 135.785000  1.755000 136.075000 1.800000 ;
      RECT 135.785000  1.940000 136.075000 1.985000 ;
      RECT 135.785000  3.455000 136.075000 3.500000 ;
      RECT 135.785000  3.640000 136.075000 3.685000 ;
      RECT 138.085000  1.755000 138.375000 1.800000 ;
      RECT 138.085000  1.940000 138.375000 1.985000 ;
      RECT 138.085000  3.455000 138.375000 3.500000 ;
      RECT 138.085000  3.640000 138.375000 3.685000 ;
      RECT 139.925000  1.755000 140.215000 1.800000 ;
      RECT 139.925000  1.940000 140.215000 1.985000 ;
      RECT 139.925000  3.455000 140.215000 3.500000 ;
      RECT 139.925000  3.640000 140.215000 3.685000 ;
      RECT 142.225000  1.755000 142.515000 1.800000 ;
      RECT 142.225000  1.940000 142.515000 1.985000 ;
      RECT 142.225000  3.455000 142.515000 3.500000 ;
      RECT 142.225000  3.640000 142.515000 3.685000 ;
      RECT 144.065000  1.755000 144.355000 1.800000 ;
      RECT 144.065000  1.940000 144.355000 1.985000 ;
      RECT 144.065000  3.455000 144.355000 3.500000 ;
      RECT 144.065000  3.640000 144.355000 3.685000 ;
      RECT 146.365000  1.755000 146.655000 1.800000 ;
      RECT 146.365000  1.940000 146.655000 1.985000 ;
      RECT 146.365000  3.455000 146.655000 3.500000 ;
      RECT 146.365000  3.640000 146.655000 3.685000 ;
      RECT 147.775000  2.110000 148.065000 2.155000 ;
      RECT 147.775000  2.155000 150.000000 2.295000 ;
      RECT 147.775000  2.295000 148.065000 2.340000 ;
      RECT 147.775000  3.100000 148.065000 3.145000 ;
      RECT 147.775000  3.145000 150.000000 3.285000 ;
      RECT 147.775000  3.285000 148.065000 3.330000 ;
      RECT 148.715000  2.110000 149.005000 2.155000 ;
      RECT 148.715000  2.295000 149.005000 2.340000 ;
      RECT 148.715000  3.100000 149.005000 3.145000 ;
      RECT 148.715000  3.285000 149.005000 3.330000 ;
      RECT 149.125000  1.755000 149.415000 1.800000 ;
      RECT 149.125000  1.800000 171.955000 1.940000 ;
      RECT 149.125000  1.940000 149.415000 1.985000 ;
      RECT 149.125000  3.455000 149.415000 3.500000 ;
      RECT 149.125000  3.500000 171.955000 3.640000 ;
      RECT 149.125000  3.640000 149.415000 3.685000 ;
      RECT 149.710000  2.110000 150.000000 2.155000 ;
      RECT 149.710000  2.295000 150.000000 2.340000 ;
      RECT 149.710000  3.100000 150.000000 3.145000 ;
      RECT 149.710000  3.285000 150.000000 3.330000 ;
      RECT 151.760000  2.110000 152.050000 2.155000 ;
      RECT 151.760000  2.155000 153.985000 2.295000 ;
      RECT 151.760000  2.295000 152.050000 2.340000 ;
      RECT 151.760000  3.100000 152.050000 3.145000 ;
      RECT 151.760000  3.145000 153.985000 3.285000 ;
      RECT 151.760000  3.285000 152.050000 3.330000 ;
      RECT 152.345000  1.755000 152.635000 1.800000 ;
      RECT 152.345000  1.940000 152.635000 1.985000 ;
      RECT 152.345000  3.455000 152.635000 3.500000 ;
      RECT 152.345000  3.640000 152.635000 3.685000 ;
      RECT 152.755000  2.110000 153.045000 2.155000 ;
      RECT 152.755000  2.295000 153.045000 2.340000 ;
      RECT 152.755000  3.100000 153.045000 3.145000 ;
      RECT 152.755000  3.285000 153.045000 3.330000 ;
      RECT 153.695000  2.110000 153.985000 2.155000 ;
      RECT 153.695000  2.295000 153.985000 2.340000 ;
      RECT 153.695000  3.100000 153.985000 3.145000 ;
      RECT 153.695000  3.285000 153.985000 3.330000 ;
      RECT 154.215000  2.110000 154.505000 2.155000 ;
      RECT 154.215000  2.155000 156.440000 2.295000 ;
      RECT 154.215000  2.295000 154.505000 2.340000 ;
      RECT 154.215000  3.100000 154.505000 3.145000 ;
      RECT 154.215000  3.145000 156.440000 3.285000 ;
      RECT 154.215000  3.285000 154.505000 3.330000 ;
      RECT 155.155000  2.110000 155.445000 2.155000 ;
      RECT 155.155000  2.295000 155.445000 2.340000 ;
      RECT 155.155000  3.100000 155.445000 3.145000 ;
      RECT 155.155000  3.285000 155.445000 3.330000 ;
      RECT 155.565000  1.755000 155.855000 1.800000 ;
      RECT 155.565000  1.940000 155.855000 1.985000 ;
      RECT 155.565000  3.455000 155.855000 3.500000 ;
      RECT 155.565000  3.640000 155.855000 3.685000 ;
      RECT 156.150000  2.110000 156.440000 2.155000 ;
      RECT 156.150000  2.295000 156.440000 2.340000 ;
      RECT 156.150000  3.100000 156.440000 3.145000 ;
      RECT 156.150000  3.285000 156.440000 3.330000 ;
      RECT 158.200000  2.110000 158.490000 2.155000 ;
      RECT 158.200000  2.155000 160.425000 2.295000 ;
      RECT 158.200000  2.295000 158.490000 2.340000 ;
      RECT 158.200000  3.100000 158.490000 3.145000 ;
      RECT 158.200000  3.145000 160.425000 3.285000 ;
      RECT 158.200000  3.285000 158.490000 3.330000 ;
      RECT 158.785000  1.755000 159.075000 1.800000 ;
      RECT 158.785000  1.940000 159.075000 1.985000 ;
      RECT 158.785000  3.455000 159.075000 3.500000 ;
      RECT 158.785000  3.640000 159.075000 3.685000 ;
      RECT 159.195000  2.110000 159.485000 2.155000 ;
      RECT 159.195000  2.295000 159.485000 2.340000 ;
      RECT 159.195000  3.100000 159.485000 3.145000 ;
      RECT 159.195000  3.285000 159.485000 3.330000 ;
      RECT 160.135000  2.110000 160.425000 2.155000 ;
      RECT 160.135000  2.295000 160.425000 2.340000 ;
      RECT 160.135000  3.100000 160.425000 3.145000 ;
      RECT 160.135000  3.285000 160.425000 3.330000 ;
      RECT 160.655000  2.110000 160.945000 2.155000 ;
      RECT 160.655000  2.155000 162.880000 2.295000 ;
      RECT 160.655000  2.295000 160.945000 2.340000 ;
      RECT 160.655000  3.100000 160.945000 3.145000 ;
      RECT 160.655000  3.145000 162.880000 3.285000 ;
      RECT 160.655000  3.285000 160.945000 3.330000 ;
      RECT 161.595000  2.110000 161.885000 2.155000 ;
      RECT 161.595000  2.295000 161.885000 2.340000 ;
      RECT 161.595000  3.100000 161.885000 3.145000 ;
      RECT 161.595000  3.285000 161.885000 3.330000 ;
      RECT 162.005000  1.755000 162.295000 1.800000 ;
      RECT 162.005000  1.940000 162.295000 1.985000 ;
      RECT 162.005000  3.455000 162.295000 3.500000 ;
      RECT 162.005000  3.640000 162.295000 3.685000 ;
      RECT 162.590000  2.110000 162.880000 2.155000 ;
      RECT 162.590000  2.295000 162.880000 2.340000 ;
      RECT 162.590000  3.100000 162.880000 3.145000 ;
      RECT 162.590000  3.285000 162.880000 3.330000 ;
      RECT 164.640000  2.110000 164.930000 2.155000 ;
      RECT 164.640000  2.155000 166.865000 2.295000 ;
      RECT 164.640000  2.295000 164.930000 2.340000 ;
      RECT 164.640000  3.100000 164.930000 3.145000 ;
      RECT 164.640000  3.145000 166.865000 3.285000 ;
      RECT 164.640000  3.285000 164.930000 3.330000 ;
      RECT 165.225000  1.755000 165.515000 1.800000 ;
      RECT 165.225000  1.940000 165.515000 1.985000 ;
      RECT 165.225000  3.455000 165.515000 3.500000 ;
      RECT 165.225000  3.640000 165.515000 3.685000 ;
      RECT 165.635000  2.110000 165.925000 2.155000 ;
      RECT 165.635000  2.295000 165.925000 2.340000 ;
      RECT 165.635000  3.100000 165.925000 3.145000 ;
      RECT 165.635000  3.285000 165.925000 3.330000 ;
      RECT 166.575000  2.110000 166.865000 2.155000 ;
      RECT 166.575000  2.295000 166.865000 2.340000 ;
      RECT 166.575000  3.100000 166.865000 3.145000 ;
      RECT 166.575000  3.285000 166.865000 3.330000 ;
      RECT 167.095000  2.110000 167.385000 2.155000 ;
      RECT 167.095000  2.155000 169.320000 2.295000 ;
      RECT 167.095000  2.295000 167.385000 2.340000 ;
      RECT 167.095000  3.100000 167.385000 3.145000 ;
      RECT 167.095000  3.145000 169.320000 3.285000 ;
      RECT 167.095000  3.285000 167.385000 3.330000 ;
      RECT 168.035000  2.110000 168.325000 2.155000 ;
      RECT 168.035000  2.295000 168.325000 2.340000 ;
      RECT 168.035000  3.100000 168.325000 3.145000 ;
      RECT 168.035000  3.285000 168.325000 3.330000 ;
      RECT 168.445000  1.755000 168.735000 1.800000 ;
      RECT 168.445000  1.940000 168.735000 1.985000 ;
      RECT 168.445000  3.455000 168.735000 3.500000 ;
      RECT 168.445000  3.640000 168.735000 3.685000 ;
      RECT 169.030000  2.110000 169.320000 2.155000 ;
      RECT 169.030000  2.295000 169.320000 2.340000 ;
      RECT 169.030000  3.100000 169.320000 3.145000 ;
      RECT 169.030000  3.285000 169.320000 3.330000 ;
      RECT 171.080000  2.110000 171.370000 2.155000 ;
      RECT 171.080000  2.155000 173.305000 2.295000 ;
      RECT 171.080000  2.295000 171.370000 2.340000 ;
      RECT 171.080000  3.100000 171.370000 3.145000 ;
      RECT 171.080000  3.145000 173.305000 3.285000 ;
      RECT 171.080000  3.285000 171.370000 3.330000 ;
      RECT 171.665000  1.755000 171.955000 1.800000 ;
      RECT 171.665000  1.940000 171.955000 1.985000 ;
      RECT 171.665000  3.455000 171.955000 3.500000 ;
      RECT 171.665000  3.640000 171.955000 3.685000 ;
      RECT 172.075000  2.110000 172.365000 2.155000 ;
      RECT 172.075000  2.295000 172.365000 2.340000 ;
      RECT 172.075000  3.100000 172.365000 3.145000 ;
      RECT 172.075000  3.285000 172.365000 3.330000 ;
      RECT 173.015000  2.110000 173.305000 2.155000 ;
      RECT 173.015000  2.295000 173.305000 2.340000 ;
      RECT 173.015000  3.100000 173.305000 3.145000 ;
      RECT 173.015000  3.285000 173.305000 3.330000 ;
      RECT 174.005000  2.110000 174.295000 2.155000 ;
      RECT 174.005000  2.155000 178.115000 2.295000 ;
      RECT 174.005000  2.295000 174.295000 2.340000 ;
      RECT 174.005000  3.100000 174.295000 3.145000 ;
      RECT 174.005000  3.145000 178.115000 3.285000 ;
      RECT 174.005000  3.285000 174.295000 3.330000 ;
      RECT 174.945000  2.110000 175.235000 2.155000 ;
      RECT 174.945000  2.295000 175.235000 2.340000 ;
      RECT 174.945000  3.100000 175.235000 3.145000 ;
      RECT 174.945000  3.285000 175.235000 3.330000 ;
      RECT 175.925000  2.110000 176.215000 2.155000 ;
      RECT 175.925000  2.295000 176.215000 2.340000 ;
      RECT 175.925000  3.100000 176.215000 3.145000 ;
      RECT 175.925000  3.285000 176.215000 3.330000 ;
      RECT 176.405000  1.755000 176.695000 1.800000 ;
      RECT 176.405000  1.800000 222.415000 1.940000 ;
      RECT 176.405000  1.940000 176.695000 1.985000 ;
      RECT 176.405000  3.455000 176.695000 3.500000 ;
      RECT 176.405000  3.500000 222.415000 3.640000 ;
      RECT 176.405000  3.640000 176.695000 3.685000 ;
      RECT 176.875000  2.110000 177.165000 2.155000 ;
      RECT 176.875000  2.295000 177.165000 2.340000 ;
      RECT 176.875000  3.100000 177.165000 3.145000 ;
      RECT 176.875000  3.285000 177.165000 3.330000 ;
      RECT 177.345000  1.755000 177.635000 1.800000 ;
      RECT 177.345000  1.940000 177.635000 1.985000 ;
      RECT 177.345000  3.455000 177.635000 3.500000 ;
      RECT 177.345000  3.640000 177.635000 3.685000 ;
      RECT 177.825000  2.110000 178.115000 2.155000 ;
      RECT 177.825000  2.295000 178.115000 2.340000 ;
      RECT 177.825000  3.100000 178.115000 3.145000 ;
      RECT 177.825000  3.285000 178.115000 3.330000 ;
      RECT 181.605000  2.110000 181.895000 2.155000 ;
      RECT 181.605000  2.155000 185.715000 2.295000 ;
      RECT 181.605000  2.295000 181.895000 2.340000 ;
      RECT 181.605000  3.100000 181.895000 3.145000 ;
      RECT 181.605000  3.145000 185.715000 3.285000 ;
      RECT 181.605000  3.285000 181.895000 3.330000 ;
      RECT 182.085000  1.755000 182.375000 1.800000 ;
      RECT 182.085000  1.940000 182.375000 1.985000 ;
      RECT 182.085000  3.455000 182.375000 3.500000 ;
      RECT 182.085000  3.640000 182.375000 3.685000 ;
      RECT 182.555000  2.110000 182.845000 2.155000 ;
      RECT 182.555000  2.295000 182.845000 2.340000 ;
      RECT 182.555000  3.100000 182.845000 3.145000 ;
      RECT 182.555000  3.285000 182.845000 3.330000 ;
      RECT 183.025000  1.755000 183.315000 1.800000 ;
      RECT 183.025000  1.940000 183.315000 1.985000 ;
      RECT 183.025000  3.455000 183.315000 3.500000 ;
      RECT 183.025000  3.640000 183.315000 3.685000 ;
      RECT 183.505000  2.110000 183.795000 2.155000 ;
      RECT 183.505000  2.295000 183.795000 2.340000 ;
      RECT 183.505000  3.100000 183.795000 3.145000 ;
      RECT 183.505000  3.285000 183.795000 3.330000 ;
      RECT 184.485000  2.110000 184.775000 2.155000 ;
      RECT 184.485000  2.295000 184.775000 2.340000 ;
      RECT 184.485000  3.100000 184.775000 3.145000 ;
      RECT 184.485000  3.285000 184.775000 3.330000 ;
      RECT 185.425000  2.110000 185.715000 2.155000 ;
      RECT 185.425000  2.295000 185.715000 2.340000 ;
      RECT 185.425000  3.100000 185.715000 3.145000 ;
      RECT 185.425000  3.285000 185.715000 3.330000 ;
      RECT 186.885000  2.110000 187.175000 2.155000 ;
      RECT 186.885000  2.155000 190.995000 2.295000 ;
      RECT 186.885000  2.295000 187.175000 2.340000 ;
      RECT 186.885000  3.100000 187.175000 3.145000 ;
      RECT 186.885000  3.145000 190.995000 3.285000 ;
      RECT 186.885000  3.285000 187.175000 3.330000 ;
      RECT 187.825000  2.110000 188.115000 2.155000 ;
      RECT 187.825000  2.295000 188.115000 2.340000 ;
      RECT 187.825000  3.100000 188.115000 3.145000 ;
      RECT 187.825000  3.285000 188.115000 3.330000 ;
      RECT 188.805000  2.110000 189.095000 2.155000 ;
      RECT 188.805000  2.295000 189.095000 2.340000 ;
      RECT 188.805000  3.100000 189.095000 3.145000 ;
      RECT 188.805000  3.285000 189.095000 3.330000 ;
      RECT 189.285000  1.755000 189.575000 1.800000 ;
      RECT 189.285000  1.940000 189.575000 1.985000 ;
      RECT 189.285000  3.455000 189.575000 3.500000 ;
      RECT 189.285000  3.640000 189.575000 3.685000 ;
      RECT 189.755000  2.110000 190.045000 2.155000 ;
      RECT 189.755000  2.295000 190.045000 2.340000 ;
      RECT 189.755000  3.100000 190.045000 3.145000 ;
      RECT 189.755000  3.285000 190.045000 3.330000 ;
      RECT 190.225000  1.755000 190.515000 1.800000 ;
      RECT 190.225000  1.940000 190.515000 1.985000 ;
      RECT 190.225000  3.455000 190.515000 3.500000 ;
      RECT 190.225000  3.640000 190.515000 3.685000 ;
      RECT 190.705000  2.110000 190.995000 2.155000 ;
      RECT 190.705000  2.295000 190.995000 2.340000 ;
      RECT 190.705000  3.100000 190.995000 3.145000 ;
      RECT 190.705000  3.285000 190.995000 3.330000 ;
      RECT 194.485000  2.110000 194.775000 2.155000 ;
      RECT 194.485000  2.155000 198.595000 2.295000 ;
      RECT 194.485000  2.295000 194.775000 2.340000 ;
      RECT 194.485000  3.100000 194.775000 3.145000 ;
      RECT 194.485000  3.145000 198.595000 3.285000 ;
      RECT 194.485000  3.285000 194.775000 3.330000 ;
      RECT 194.965000  1.755000 195.255000 1.800000 ;
      RECT 194.965000  1.940000 195.255000 1.985000 ;
      RECT 194.965000  3.455000 195.255000 3.500000 ;
      RECT 194.965000  3.640000 195.255000 3.685000 ;
      RECT 195.435000  2.110000 195.725000 2.155000 ;
      RECT 195.435000  2.295000 195.725000 2.340000 ;
      RECT 195.435000  3.100000 195.725000 3.145000 ;
      RECT 195.435000  3.285000 195.725000 3.330000 ;
      RECT 195.905000  1.755000 196.195000 1.800000 ;
      RECT 195.905000  1.940000 196.195000 1.985000 ;
      RECT 195.905000  3.455000 196.195000 3.500000 ;
      RECT 195.905000  3.640000 196.195000 3.685000 ;
      RECT 196.385000  2.110000 196.675000 2.155000 ;
      RECT 196.385000  2.295000 196.675000 2.340000 ;
      RECT 196.385000  3.100000 196.675000 3.145000 ;
      RECT 196.385000  3.285000 196.675000 3.330000 ;
      RECT 197.365000  2.110000 197.655000 2.155000 ;
      RECT 197.365000  2.295000 197.655000 2.340000 ;
      RECT 197.365000  3.100000 197.655000 3.145000 ;
      RECT 197.365000  3.285000 197.655000 3.330000 ;
      RECT 198.305000  2.110000 198.595000 2.155000 ;
      RECT 198.305000  2.295000 198.595000 2.340000 ;
      RECT 198.305000  3.100000 198.595000 3.145000 ;
      RECT 198.305000  3.285000 198.595000 3.330000 ;
      RECT 200.225000  2.110000 200.515000 2.155000 ;
      RECT 200.225000  2.155000 204.335000 2.295000 ;
      RECT 200.225000  2.295000 200.515000 2.340000 ;
      RECT 200.225000  3.100000 200.515000 3.145000 ;
      RECT 200.225000  3.145000 204.335000 3.285000 ;
      RECT 200.225000  3.285000 200.515000 3.330000 ;
      RECT 201.165000  2.110000 201.455000 2.155000 ;
      RECT 201.165000  2.295000 201.455000 2.340000 ;
      RECT 201.165000  3.100000 201.455000 3.145000 ;
      RECT 201.165000  3.285000 201.455000 3.330000 ;
      RECT 202.145000  2.110000 202.435000 2.155000 ;
      RECT 202.145000  2.295000 202.435000 2.340000 ;
      RECT 202.145000  3.100000 202.435000 3.145000 ;
      RECT 202.145000  3.285000 202.435000 3.330000 ;
      RECT 202.625000  1.755000 202.915000 1.800000 ;
      RECT 202.625000  1.940000 202.915000 1.985000 ;
      RECT 202.625000  3.455000 202.915000 3.500000 ;
      RECT 202.625000  3.640000 202.915000 3.685000 ;
      RECT 203.095000  2.110000 203.385000 2.155000 ;
      RECT 203.095000  2.295000 203.385000 2.340000 ;
      RECT 203.095000  3.100000 203.385000 3.145000 ;
      RECT 203.095000  3.285000 203.385000 3.330000 ;
      RECT 203.565000  1.755000 203.855000 1.800000 ;
      RECT 203.565000  1.940000 203.855000 1.985000 ;
      RECT 203.565000  3.455000 203.855000 3.500000 ;
      RECT 203.565000  3.640000 203.855000 3.685000 ;
      RECT 204.045000  2.110000 204.335000 2.155000 ;
      RECT 204.045000  2.295000 204.335000 2.340000 ;
      RECT 204.045000  3.100000 204.335000 3.145000 ;
      RECT 204.045000  3.285000 204.335000 3.330000 ;
      RECT 207.825000  2.110000 208.115000 2.155000 ;
      RECT 207.825000  2.155000 211.935000 2.295000 ;
      RECT 207.825000  2.295000 208.115000 2.340000 ;
      RECT 207.825000  3.100000 208.115000 3.145000 ;
      RECT 207.825000  3.145000 211.935000 3.285000 ;
      RECT 207.825000  3.285000 208.115000 3.330000 ;
      RECT 208.305000  1.755000 208.595000 1.800000 ;
      RECT 208.305000  1.940000 208.595000 1.985000 ;
      RECT 208.305000  3.455000 208.595000 3.500000 ;
      RECT 208.305000  3.640000 208.595000 3.685000 ;
      RECT 208.775000  2.110000 209.065000 2.155000 ;
      RECT 208.775000  2.295000 209.065000 2.340000 ;
      RECT 208.775000  3.100000 209.065000 3.145000 ;
      RECT 208.775000  3.285000 209.065000 3.330000 ;
      RECT 209.245000  1.755000 209.535000 1.800000 ;
      RECT 209.245000  1.940000 209.535000 1.985000 ;
      RECT 209.245000  3.455000 209.535000 3.500000 ;
      RECT 209.245000  3.640000 209.535000 3.685000 ;
      RECT 209.725000  2.110000 210.015000 2.155000 ;
      RECT 209.725000  2.295000 210.015000 2.340000 ;
      RECT 209.725000  3.100000 210.015000 3.145000 ;
      RECT 209.725000  3.285000 210.015000 3.330000 ;
      RECT 210.705000  2.110000 210.995000 2.155000 ;
      RECT 210.705000  2.295000 210.995000 2.340000 ;
      RECT 210.705000  3.100000 210.995000 3.145000 ;
      RECT 210.705000  3.285000 210.995000 3.330000 ;
      RECT 211.645000  2.110000 211.935000 2.155000 ;
      RECT 211.645000  2.295000 211.935000 2.340000 ;
      RECT 211.645000  3.100000 211.935000 3.145000 ;
      RECT 211.645000  3.285000 211.935000 3.330000 ;
      RECT 213.105000  2.110000 213.395000 2.155000 ;
      RECT 213.105000  2.155000 217.215000 2.295000 ;
      RECT 213.105000  2.295000 213.395000 2.340000 ;
      RECT 213.105000  3.100000 213.395000 3.145000 ;
      RECT 213.105000  3.145000 217.215000 3.285000 ;
      RECT 213.105000  3.285000 213.395000 3.330000 ;
      RECT 214.045000  2.110000 214.335000 2.155000 ;
      RECT 214.045000  2.295000 214.335000 2.340000 ;
      RECT 214.045000  3.100000 214.335000 3.145000 ;
      RECT 214.045000  3.285000 214.335000 3.330000 ;
      RECT 215.025000  2.110000 215.315000 2.155000 ;
      RECT 215.025000  2.295000 215.315000 2.340000 ;
      RECT 215.025000  3.100000 215.315000 3.145000 ;
      RECT 215.025000  3.285000 215.315000 3.330000 ;
      RECT 215.505000  1.755000 215.795000 1.800000 ;
      RECT 215.505000  1.940000 215.795000 1.985000 ;
      RECT 215.505000  3.455000 215.795000 3.500000 ;
      RECT 215.505000  3.640000 215.795000 3.685000 ;
      RECT 215.975000  2.110000 216.265000 2.155000 ;
      RECT 215.975000  2.295000 216.265000 2.340000 ;
      RECT 215.975000  3.100000 216.265000 3.145000 ;
      RECT 215.975000  3.285000 216.265000 3.330000 ;
      RECT 216.445000  1.755000 216.735000 1.800000 ;
      RECT 216.445000  1.940000 216.735000 1.985000 ;
      RECT 216.445000  3.455000 216.735000 3.500000 ;
      RECT 216.445000  3.640000 216.735000 3.685000 ;
      RECT 216.925000  2.110000 217.215000 2.155000 ;
      RECT 216.925000  2.295000 217.215000 2.340000 ;
      RECT 216.925000  3.100000 217.215000 3.145000 ;
      RECT 216.925000  3.285000 217.215000 3.330000 ;
      RECT 220.705000  2.110000 220.995000 2.155000 ;
      RECT 220.705000  2.155000 224.815000 2.295000 ;
      RECT 220.705000  2.295000 220.995000 2.340000 ;
      RECT 220.705000  3.100000 220.995000 3.145000 ;
      RECT 220.705000  3.145000 224.815000 3.285000 ;
      RECT 220.705000  3.285000 220.995000 3.330000 ;
      RECT 221.185000  1.755000 221.475000 1.800000 ;
      RECT 221.185000  1.940000 221.475000 1.985000 ;
      RECT 221.185000  3.455000 221.475000 3.500000 ;
      RECT 221.185000  3.640000 221.475000 3.685000 ;
      RECT 221.655000  2.110000 221.945000 2.155000 ;
      RECT 221.655000  2.295000 221.945000 2.340000 ;
      RECT 221.655000  3.100000 221.945000 3.145000 ;
      RECT 221.655000  3.285000 221.945000 3.330000 ;
      RECT 222.125000  1.755000 222.415000 1.800000 ;
      RECT 222.125000  1.940000 222.415000 1.985000 ;
      RECT 222.125000  3.455000 222.415000 3.500000 ;
      RECT 222.125000  3.640000 222.415000 3.685000 ;
      RECT 222.605000  2.110000 222.895000 2.155000 ;
      RECT 222.605000  2.295000 222.895000 2.340000 ;
      RECT 222.605000  3.100000 222.895000 3.145000 ;
      RECT 222.605000  3.285000 222.895000 3.330000 ;
      RECT 223.585000  2.110000 223.875000 2.155000 ;
      RECT 223.585000  2.295000 223.875000 2.340000 ;
      RECT 223.585000  3.100000 223.875000 3.145000 ;
      RECT 223.585000  3.285000 223.875000 3.330000 ;
      RECT 224.525000  2.110000 224.815000 2.155000 ;
      RECT 224.525000  2.295000 224.815000 2.340000 ;
      RECT 224.525000  3.100000 224.815000 3.145000 ;
      RECT 224.525000  3.285000 224.815000 3.330000 ;
    LAYER nwell ;
      RECT  -0.190000 1.305000 225.590000 2.910000 ;
      RECT 105.610000 2.910000 225.590000 4.135000 ;
    LAYER pwell ;
      RECT   0.420000 -0.085000   0.640000 0.085000 ;
      RECT   5.480000 -0.085000   5.700000 0.085000 ;
      RECT  11.460000 -0.085000  11.680000 0.085000 ;
      RECT  15.785000 -0.085000  15.955000 0.085000 ;
      RECT  24.525000 -0.085000  24.695000 0.085000 ;
      RECT  30.505000 -0.085000  30.675000 0.085000 ;
      RECT  30.965000 -0.085000  31.135000 0.085000 ;
      RECT  36.945000 -0.085000  37.115000 0.085000 ;
      RECT  37.405000 -0.085000  37.575000 0.085000 ;
      RECT  49.825000 -0.085000  49.995000 0.085000 ;
      RECT  50.285000 -0.085000  50.455000 0.085000 ;
      RECT  62.705000 -0.085000  62.875000 0.085000 ;
      RECT  63.165000 -0.085000  63.335000 0.085000 ;
      RECT  67.305000 -0.085000  67.475000 0.085000 ;
      RECT  71.445000 -0.085000  71.615000 0.085000 ;
      RECT  75.585000 -0.085000  75.755000 0.085000 ;
      RECT  79.725000 -0.085000  79.895000 0.085000 ;
      RECT  80.185000 -0.085000  80.355000 0.085000 ;
      RECT  86.165000 -0.085000  86.335000 0.085000 ;
      RECT  86.625000 -0.085000  86.795000 0.085000 ;
      RECT  92.605000 -0.085000  92.775000 0.085000 ;
      RECT  93.065000 -0.085000  93.235000 0.085000 ;
      RECT  99.045000 -0.085000  99.215000 0.085000 ;
      RECT  99.505000 -0.085000  99.675000 0.085000 ;
      RECT 105.485000 -0.085000 105.655000 0.085000 ;
      RECT 105.945000 -0.085000 106.115000 0.085000 ;
      RECT 111.925000 -0.085000 112.095000 0.085000 ;
      RECT 124.345000 -0.085000 124.515000 0.085000 ;
      RECT 130.785000 -0.085000 130.955000 0.085000 ;
      RECT 134.925000 -0.085000 135.095000 0.085000 ;
      RECT 139.065000 -0.085000 139.235000 0.085000 ;
      RECT 143.205000 -0.085000 143.375000 0.085000 ;
      RECT 147.345000 -0.085000 147.515000 0.085000 ;
      RECT 147.805000 -0.085000 147.975000 0.085000 ;
      RECT 153.785000 -0.085000 153.955000 0.085000 ;
      RECT 154.245000 -0.085000 154.415000 0.085000 ;
      RECT 160.225000 -0.085000 160.395000 0.085000 ;
      RECT 160.685000 -0.085000 160.855000 0.085000 ;
      RECT 166.665000 -0.085000 166.835000 0.085000 ;
      RECT 167.125000 -0.085000 167.295000 0.085000 ;
      RECT 173.105000 -0.085000 173.275000 0.085000 ;
      RECT 173.565000 -0.085000 173.735000 0.085000 ;
      RECT 185.985000 -0.085000 186.155000 0.085000 ;
      RECT 186.445000 -0.085000 186.615000 0.085000 ;
      RECT 198.865000 -0.085000 199.035000 0.085000 ;
      RECT 199.325000  0.320000 199.495000 0.845000 ;
      RECT 199.785000 -0.085000 199.955000 0.085000 ;
      RECT 212.205000 -0.085000 212.375000 0.085000 ;
      RECT 212.665000 -0.085000 212.835000 0.085000 ;
      RECT 225.085000 -0.085000 225.255000 0.085000 ;
    LAYER pwell ;
      RECT 105.945000 5.355000 106.115000 5.525000 ;
      RECT 111.925000 5.355000 112.095000 5.525000 ;
      RECT 124.345000 5.355000 124.515000 5.525000 ;
      RECT 130.785000 5.355000 130.955000 5.525000 ;
      RECT 134.925000 5.355000 135.095000 5.525000 ;
      RECT 139.065000 5.355000 139.235000 5.525000 ;
      RECT 143.205000 5.355000 143.375000 5.525000 ;
      RECT 147.345000 5.355000 147.515000 5.525000 ;
      RECT 147.805000 5.355000 147.975000 5.525000 ;
      RECT 153.785000 5.355000 153.955000 5.525000 ;
      RECT 154.245000 5.355000 154.415000 5.525000 ;
      RECT 160.225000 5.355000 160.395000 5.525000 ;
      RECT 160.685000 5.355000 160.855000 5.525000 ;
      RECT 166.665000 5.355000 166.835000 5.525000 ;
      RECT 167.125000 5.355000 167.295000 5.525000 ;
      RECT 173.105000 5.355000 173.275000 5.525000 ;
      RECT 173.565000 5.355000 173.735000 5.525000 ;
      RECT 185.985000 5.355000 186.155000 5.525000 ;
      RECT 186.445000 5.355000 186.615000 5.525000 ;
      RECT 198.865000 5.355000 199.035000 5.525000 ;
      RECT 199.325000 4.595000 199.495000 5.120000 ;
      RECT 199.785000 5.355000 199.955000 5.525000 ;
      RECT 212.205000 5.355000 212.375000 5.525000 ;
      RECT 212.665000 5.355000 212.835000 5.525000 ;
      RECT 225.085000 5.355000 225.255000 5.525000 ;
  END
END sky130_fd_sc_hdll__muxb
END LIBRARY
