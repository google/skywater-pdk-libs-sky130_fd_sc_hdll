* File: sky130_fd_sc_hdll__mux2_2.pex.spice
* Created: Wed Sep  2 08:34:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUX2_2%A_79_21# 1 2 7 9 10 12 13 15 16 18 22 23 24
+ 25 26 28 29 31 33 35 38 40 49
c111 26 0 1.7675e-19 $X=1.265 $Y=1.92
r112 48 49 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r113 47 48 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.94 $Y2=1.202
r114 46 47 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r115 39 49 11.6613 $w=3.72e-07 $l=9e-08 $layer=POLY_cond $X=1.055 $Y=1.202
+ $X2=0.965 $Y2=1.202
r116 38 41 8.49766 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.117 $Y=1.16
+ $X2=1.117 $Y2=1.325
r117 38 40 8.49766 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.117 $Y=1.16
+ $X2=1.117 $Y2=0.995
r118 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.055
+ $Y=1.16 $X2=1.055 $Y2=1.16
r119 33 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.62 $Y=0.43
+ $X2=1.62 $Y2=0.72
r120 33 35 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.705 $Y=0.43
+ $X2=2.165 $Y2=0.43
r121 29 31 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=1.625 $Y=2.34
+ $X2=2.695 $Y2=2.34
r122 28 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.54 $Y=2.255
+ $X2=1.625 $Y2=2.34
r123 27 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.54 $Y=2.005
+ $X2=1.54 $Y2=2.255
r124 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.455 $Y=1.92
+ $X2=1.54 $Y2=2.005
r125 25 26 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.92
+ $X2=1.265 $Y2=1.92
r126 23 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=0.72
+ $X2=1.62 $Y2=0.72
r127 23 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.535 $Y=0.72
+ $X2=1.265 $Y2=0.72
r128 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=1.835
+ $X2=1.265 $Y2=1.92
r129 22 41 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.18 $Y=1.835
+ $X2=1.18 $Y2=1.325
r130 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=0.805
+ $X2=1.265 $Y2=0.72
r131 19 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.18 $Y=0.805
+ $X2=1.18 $Y2=0.995
r132 16 49 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r133 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r134 13 48 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r135 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r136 10 47 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r137 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r138 7 46 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r139 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r140 2 31 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=2.55
+ $Y=1.845 $X2=2.695 $Y2=2.34
r141 1 35 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=2.03
+ $Y=0.235 $X2=2.165 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_2%A_280_21# 1 2 9 12 13 15 18 19 22 23 24 29
+ 33 36
c90 24 0 1.25191e-19 $X=1.965 $Y=1.92
r91 27 36 2.99104 $w=3.17e-07 $l=1.14039e-07 $layer=LI1_cond $X=4.11 $Y=1.835
+ $X2=4.042 $Y2=1.92
r92 27 29 65.2283 $w=2.48e-07 $l=1.415e-06 $layer=LI1_cond $X=4.11 $Y=1.835
+ $X2=4.11 $Y2=0.42
r93 23 36 3.66292 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.85 $Y=1.92
+ $X2=4.042 $Y2=1.92
r94 23 24 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=3.85 $Y=1.92
+ $X2=1.965 $Y2=1.92
r95 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.88 $Y=1.835
+ $X2=1.965 $Y2=1.92
r96 21 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=1.665
+ $X2=1.88 $Y2=1.58
r97 21 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.88 $Y=1.665
+ $X2=1.88 $Y2=1.835
r98 19 39 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.535 $Y=1.16
+ $X2=1.535 $Y2=1.325
r99 19 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.535 $Y=1.16
+ $X2=1.535 $Y2=0.995
r100 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.535
+ $Y=1.16 $X2=1.535 $Y2=1.16
r101 16 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.545 $Y=1.58
+ $X2=1.88 $Y2=1.58
r102 16 18 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=1.545 $Y=1.495
+ $X2=1.545 $Y2=1.16
r103 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.5 $Y=1.77
+ $X2=1.5 $Y2=2.165
r104 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.5 $Y=1.67 $X2=1.5
+ $Y2=1.77
r105 12 39 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=1.5 $Y=1.67 $X2=1.5
+ $Y2=1.325
r106 9 38 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.475 $Y=0.445
+ $X2=1.475 $Y2=0.995
r107 2 36 300 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_PDIFF $count=2 $X=3.91
+ $Y=1.845 $X2=4.065 $Y2=2
r108 1 29 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.235 $X2=4.07 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_2%A0 3 4 6 7 9 10 11 12 18 20 31 34
r55 23 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.905
+ $Y=1.45 $X2=2.905 $Y2=1.45
r56 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=0.93
+ $X2=2.015 $Y2=0.765
r57 12 34 2.83935 $w=3.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=1.452
+ $X2=2.905 $Y2=1.452
r58 11 34 12.5266 $w=3.43e-07 $l=3.75e-07 $layer=LI1_cond $X=2.53 $Y=1.452
+ $X2=2.905 $Y2=1.452
r59 11 31 0.167021 $w=3.43e-07 $l=5e-09 $layer=LI1_cond $X=2.53 $Y=1.452
+ $X2=2.525 $Y2=1.452
r60 9 10 10.4488 $w=3.73e-07 $l=3.4e-07 $layer=LI1_cond $X=2.107 $Y=0.85
+ $X2=2.107 $Y2=1.19
r61 9 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=0.93 $X2=2.015 $Y2=0.93
r62 8 10 2.76586 $w=3.73e-07 $l=9e-08 $layer=LI1_cond $X=2.107 $Y=1.28 $X2=2.107
+ $Y2=1.19
r63 7 31 7.68295 $w=3.43e-07 $l=2.3e-07 $layer=LI1_cond $X=2.295 $Y=1.452
+ $X2=2.525 $Y2=1.452
r64 7 8 14.6175 $w=1.68e-07 $l=2.60154e-07 $layer=LI1_cond $X=2.295 $Y=1.452
+ $X2=2.107 $Y2=1.28
r65 4 23 66.0793 $w=2.47e-07 $l=3.37046e-07 $layer=POLY_cond $X=2.94 $Y=1.77
+ $X2=2.905 $Y2=1.45
r66 4 6 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.94 $Y=1.77 $X2=2.94
+ $Y2=2.165
r67 3 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.955 $Y=0.445
+ $X2=1.955 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_2%A1 3 6 7 9 10 13 15 16 25
r48 20 22 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.435 $Y=0.94
+ $X2=2.46 $Y2=0.94
r49 16 25 4.51862 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=2.972 $Y=0.94
+ $X2=2.972 $Y2=0.775
r50 16 25 0.27051 $w=2.03e-07 $l=5e-09 $layer=LI1_cond $X=2.972 $Y=0.77
+ $X2=2.972 $Y2=0.775
r51 15 16 14.0665 $w=2.03e-07 $l=2.6e-07 $layer=LI1_cond $X=2.972 $Y=0.51
+ $X2=2.972 $Y2=0.77
r52 13 22 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=2.615 $Y=0.94
+ $X2=2.46 $Y2=0.94
r53 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.615
+ $Y=0.94 $X2=2.615 $Y2=0.94
r54 10 16 2.79333 $w=3.3e-07 $l=1.02e-07 $layer=LI1_cond $X=2.87 $Y=0.94
+ $X2=2.972 $Y2=0.94
r55 10 12 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.87 $Y=0.94
+ $X2=2.615 $Y2=0.94
r56 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.46 $Y=1.77 $X2=2.46
+ $Y2=2.165
r57 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.46 $Y=1.67 $X2=2.46
+ $Y2=1.77
r58 5 22 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=2.46 $Y=1.075 $X2=2.46
+ $Y2=0.94
r59 5 6 197.288 $w=2e-07 $l=5.95e-07 $layer=POLY_cond $X=2.46 $Y=1.075 $X2=2.46
+ $Y2=1.67
r60 1 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.435 $Y=0.805
+ $X2=2.435 $Y2=0.94
r61 1 3 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.435 $Y=0.805
+ $X2=2.435 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_2%S 3 6 7 9 11 12 14 17 19 20 21 32
r48 31 32 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.82 $Y=1.16
+ $X2=3.845 $Y2=1.16
r49 29 31 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=3.45 $Y=1.16
+ $X2=3.82 $Y2=1.16
r50 27 29 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=3.35 $Y=1.16 $X2=3.45
+ $Y2=1.16
r51 25 27 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.325 $Y=1.16
+ $X2=3.35 $Y2=1.16
r52 20 21 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.45 $Y=1.16
+ $X2=3.45 $Y2=1.53
r53 20 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.45
+ $Y=1.16 $X2=3.45 $Y2=1.16
r54 19 20 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=3.45 $Y=0.85
+ $X2=3.45 $Y2=1.16
r55 15 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=0.995
+ $X2=3.845 $Y2=1.16
r56 15 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.845 $Y=0.995
+ $X2=3.845 $Y2=0.445
r57 12 14 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.82 $Y=1.77
+ $X2=3.82 $Y2=2.165
r58 11 12 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.82 $Y=1.67 $X2=3.82
+ $Y2=1.77
r59 10 31 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.82 $Y=1.325
+ $X2=3.82 $Y2=1.16
r60 10 11 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=3.82 $Y=1.325
+ $X2=3.82 $Y2=1.67
r61 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.35 $Y=1.77 $X2=3.35
+ $Y2=2.165
r62 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.35 $Y=1.67 $X2=3.35
+ $Y2=1.77
r63 5 27 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=1.325 $X2=3.35
+ $Y2=1.16
r64 5 6 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=3.35 $Y=1.325 $X2=3.35
+ $Y2=1.67
r65 1 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.325 $Y=0.995
+ $X2=3.325 $Y2=1.16
r66 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.325 $Y=0.995
+ $X2=3.325 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_2%VPWR 1 2 3 10 12 16 20 24 27 28 29 39 40 46
c61 16 0 1.7675e-19 $X=1.115 $Y=2.72
r62 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r64 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r65 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 34 37 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 33 36 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r69 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r70 31 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72 $X2=1.2
+ $Y2=2.72
r71 31 33 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 29 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r73 29 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 27 36 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.46 $Y=2.72 $X2=3.45
+ $Y2=2.72
r75 27 28 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.46 $Y=2.72 $X2=3.57
+ $Y2=2.72
r76 26 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.68 $Y=2.72 $X2=4.37
+ $Y2=2.72
r77 26 28 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.68 $Y=2.72 $X2=3.57
+ $Y2=2.72
r78 22 28 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=2.635
+ $X2=3.57 $Y2=2.72
r79 22 24 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=3.57 $Y=2.635
+ $X2=3.57 $Y2=2.34
r80 18 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r81 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.34
r82 17 43 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r83 16 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72 $X2=1.2
+ $Y2=2.72
r84 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r85 12 15 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r86 10 43 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r87 10 15 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r88 3 24 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.845 $X2=3.585 $Y2=2.34
r89 2 20 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r90 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r91 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_2%X 1 2 9 11 13 14
r24 14 20 8.00308 $w=3.58e-07 $l=2.5e-07 $layer=LI1_cond $X=0.695 $Y=2.21
+ $X2=0.695 $Y2=1.96
r25 13 20 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=0.695 $Y=1.87
+ $X2=0.695 $Y2=1.96
r26 11 13 3.04117 $w=3.58e-07 $l=9.5e-08 $layer=LI1_cond $X=0.695 $Y=1.775
+ $X2=0.695 $Y2=1.87
r27 11 12 6.29484 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.695 $Y=1.775
+ $X2=0.695 $Y2=1.595
r28 9 12 47.513 $w=2.83e-07 $l=1.175e-06 $layer=LI1_cond $X=0.657 $Y=0.42
+ $X2=0.657 $Y2=1.595
r29 2 20 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
r30 1 9 182 $w=1.7e-07 $l=2.56271e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.715 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_2%VGND 1 2 3 10 12 16 19 20 21 23 36 37 44
r65 44 47 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.175
+ $Y2=0.38
r66 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r67 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r68 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r69 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r70 31 34 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=3.45
+ $Y2=0
r71 31 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r72 30 33 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=3.45
+ $Y2=0
r73 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r74 28 44 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.175
+ $Y2=0
r75 28 30 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r76 27 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r77 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r78 24 40 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r79 24 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r80 23 44 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.175
+ $Y2=0
r81 23 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.69
+ $Y2=0
r82 21 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r83 21 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r84 19 33 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.45
+ $Y2=0
r85 19 20 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.585
+ $Y2=0
r86 18 36 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=4.37
+ $Y2=0
r87 18 20 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.585
+ $Y2=0
r88 14 20 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0
r89 14 16 18.5773 $w=1.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0.42
r90 10 40 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.172 $Y2=0
r91 10 12 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.217 $Y2=0.38
r92 3 16 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=3.4
+ $Y=0.235 $X2=3.585 $Y2=0.42
r93 2 47 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.38
r94 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

