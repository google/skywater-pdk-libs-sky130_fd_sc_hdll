* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__ebufn_8 A TE_B VGND VNB VPB VPWR Z
X0 a_437_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X1 a_437_309# a_124_297# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_124_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Z a_124_297# a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Z a_124_297# a_437_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_485_47# a_321_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND a_321_47# a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Z a_124_297# a_437_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 Z a_124_297# a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR TE_B a_437_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X10 VGND A a_124_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_485_47# a_124_297# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_485_47# a_321_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_124_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_485_47# a_124_297# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_437_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X16 a_437_309# a_124_297# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 VGND TE_B a_321_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_485_47# a_321_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Z a_124_297# a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VPWR TE_B a_321_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 a_437_309# a_124_297# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_485_47# a_124_297# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR TE_B a_437_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X24 VPWR A a_124_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 a_437_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X26 a_485_47# a_321_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR TE_B a_437_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X28 Z a_124_297# a_437_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_485_47# a_124_297# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 Z a_124_297# a_437_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 Z a_124_297# a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_437_309# a_124_297# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 VGND a_321_47# a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 VGND a_321_47# a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_437_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X36 VGND a_321_47# a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VPWR TE_B a_437_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
.ends
