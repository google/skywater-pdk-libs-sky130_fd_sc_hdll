* File: sky130_fd_sc_hdll__mux2_1.pex.spice
* Created: Thu Aug 27 19:10:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUX2_1%A_79_21# 1 2 7 9 10 12 15 18 19 21 22 24 26
c70 26 0 1.9931e-19 $X=1.525 $Y=0.54
r71 26 28 9.72055 $w=4.33e-07 $l=3.45e-07 $layer=LI1_cond $X=1.525 $Y=0.54
+ $X2=1.87 $Y2=0.54
r72 22 24 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.61 $Y=2.04
+ $X2=2.535 $Y2=2.04
r73 21 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.525 $Y=1.955
+ $X2=1.61 $Y2=2.04
r74 20 26 6.26295 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=1.525 $Y=0.825
+ $X2=1.525 $Y2=0.54
r75 20 21 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=1.525 $Y=0.825
+ $X2=1.525 $Y2=1.955
r76 18 26 7.20249 $w=4.33e-07 $l=2.40832e-07 $layer=LI1_cond $X=1.435 $Y=0.74
+ $X2=1.525 $Y2=0.54
r77 18 19 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.435 $Y=0.74
+ $X2=0.685 $Y2=0.74
r78 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r79 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=0.825
+ $X2=0.685 $Y2=0.74
r80 13 15 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.6 $Y=0.825
+ $X2=0.6 $Y2=1.16
r81 10 16 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.565 $Y2=1.16
r82 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r83 7 16 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.565 $Y2=1.16
r84 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
r85 2 24 300 $w=1.7e-07 $l=8.05528e-07 $layer=licon1_PDIFF $count=2 $X=1.81
+ $Y=1.87 $X2=2.535 $Y2=2.04
r86 1 28 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=1.735
+ $Y=0.235 $X2=1.87 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_1%S 2 3 5 8 10 12 15 18 19 20 21 22 24 25 28
+ 29 44
c91 8 0 4.11942e-20 $X=1.15 $Y=0.445
r92 37 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.83
+ $Y=1.545 $X2=3.83 $Y2=1.545
r93 29 44 3.50239 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=3.89 $Y=1.535 $X2=3.83
+ $Y2=1.535
r94 28 44 20.8976 $w=1.88e-07 $l=3.58e-07 $layer=LI1_cond $X=3.472 $Y=1.535
+ $X2=3.83 $Y2=1.535
r95 25 35 40.3353 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.16
+ $X2=1.085 $Y2=1.325
r96 25 34 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.16
+ $X2=1.085 $Y2=0.995
r97 24 27 7.79239 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.132 $Y=1.16
+ $X2=1.132 $Y2=1.325
r98 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.16 $X2=1.08 $Y2=1.16
r99 21 28 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.33 $Y=1.63 $X2=3.33
+ $Y2=1.535
r100 21 22 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.33 $Y=1.63
+ $X2=3.33 $Y2=2.295
r101 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=2.38
+ $X2=3.33 $Y2=2.295
r102 19 20 128.85 $w=1.68e-07 $l=1.975e-06 $layer=LI1_cond $X=3.245 $Y=2.38
+ $X2=1.27 $Y2=2.38
r103 18 20 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.17 $Y=2.295
+ $X2=1.27 $Y2=2.38
r104 18 27 53.7909 $w=1.98e-07 $l=9.7e-07 $layer=LI1_cond $X=1.17 $Y=2.295
+ $X2=1.17 $Y2=1.325
r105 13 37 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.94 $Y=1.38
+ $X2=3.855 $Y2=1.545
r106 13 15 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=3.94 $Y=1.38
+ $X2=3.94 $Y2=0.445
r107 10 37 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=3.915 $Y=1.795
+ $X2=3.855 $Y2=1.545
r108 10 12 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.915 $Y=1.795
+ $X2=3.915 $Y2=2.08
r109 8 34 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.15 $Y=0.445
+ $X2=1.15 $Y2=0.995
r110 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.125 $Y=1.795
+ $X2=1.125 $Y2=2.08
r111 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.125 $Y=1.695 $X2=1.125
+ $Y2=1.795
r112 2 35 122.684 $w=2e-07 $l=3.7e-07 $layer=POLY_cond $X=1.125 $Y=1.695
+ $X2=1.125 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_1%A1 3 5 7 10 11 13 14 16 17
c62 13 0 1.9722e-19 $X=2.855 $Y=1.7
c63 10 0 4.11942e-20 $X=1.865 $Y=0.98
r64 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.94
+ $Y=1.545 $X2=2.94 $Y2=1.545
r65 16 26 18.5962 $w=2.18e-07 $l=3.55e-07 $layer=LI1_cond $X=2.965 $Y=1.19
+ $X2=2.965 $Y2=1.545
r66 16 17 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.965 $Y=1.19
+ $X2=2.965 $Y2=0.85
r67 15 26 3.66686 $w=2.18e-07 $l=7e-08 $layer=LI1_cond $X=2.965 $Y=1.615
+ $X2=2.965 $Y2=1.545
r68 13 15 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.855 $Y=1.7
+ $X2=2.965 $Y2=1.615
r69 13 14 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.855 $Y=1.7
+ $X2=1.95 $Y2=1.7
r70 11 20 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.865 $Y=0.98
+ $X2=1.66 $Y2=0.98
r71 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=0.98 $X2=1.865 $Y2=0.98
r72 8 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.865 $Y=1.615
+ $X2=1.95 $Y2=1.7
r73 8 10 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.865 $Y=1.615
+ $X2=1.865 $Y2=0.98
r74 5 25 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.975 $Y=1.795
+ $X2=2.94 $Y2=1.545
r75 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.975 $Y=1.795
+ $X2=2.975 $Y2=2.08
r76 1 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=0.815
+ $X2=1.66 $Y2=0.98
r77 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.66 $Y=0.815 $X2=1.66
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_1%A0 1 3 4 5 8 11 12 15 16
r47 15 18 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=0.98
+ $X2=2.505 $Y2=1.145
r48 15 17 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=0.98
+ $X2=2.505 $Y2=0.815
r49 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=0.98 $X2=2.48 $Y2=0.98
r50 12 16 7.44655 $w=3.23e-07 $l=2.1e-07 $layer=LI1_cond $X=2.452 $Y=1.19
+ $X2=2.452 $Y2=0.98
r51 11 18 165.789 $w=2e-07 $l=5e-07 $layer=POLY_cond $X=2.445 $Y=1.645 $X2=2.445
+ $Y2=1.145
r52 8 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.42 $Y=0.445
+ $X2=2.42 $Y2=0.815
r53 4 11 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=2.345 $Y=1.72
+ $X2=2.445 $Y2=1.645
r54 4 5 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.345 $Y=1.72 $X2=1.81
+ $Y2=1.72
r55 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.72 $Y=1.795
+ $X2=1.81 $Y2=1.72
r56 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.72 $Y=1.795
+ $X2=1.72 $Y2=2.08
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_1%A_657_21# 1 2 9 12 13 15 16 19 23 26 27 31
c49 12 0 1.9722e-19 $X=3.385 $Y=1.695
r50 29 31 5.81843 $w=4.08e-07 $l=2.07e-07 $layer=LI1_cond $X=4.15 $Y=2.08
+ $X2=4.357 $Y2=2.08
r51 26 31 2.88189 $w=2.85e-07 $l=2.05e-07 $layer=LI1_cond $X=4.357 $Y=1.875
+ $X2=4.357 $Y2=2.08
r52 25 27 3.52026 $w=2.65e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.357 $Y=1.065
+ $X2=4.267 $Y2=0.98
r53 25 26 32.7536 $w=2.83e-07 $l=8.1e-07 $layer=LI1_cond $X=4.357 $Y=1.065
+ $X2=4.357 $Y2=1.875
r54 21 27 3.52026 $w=2.65e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.157 $Y=0.895
+ $X2=4.267 $Y2=0.98
r55 21 23 20.6969 $w=2.43e-07 $l=4.4e-07 $layer=LI1_cond $X=4.157 $Y=0.895
+ $X2=4.157 $Y2=0.455
r56 19 35 32.4954 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.45 $Y=0.98
+ $X2=3.45 $Y2=1.115
r57 19 34 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.45 $Y=0.98
+ $X2=3.45 $Y2=0.845
r58 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.45
+ $Y=0.98 $X2=3.45 $Y2=0.98
r59 16 27 2.98021 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=4.035 $Y=0.98
+ $X2=4.267 $Y2=0.98
r60 16 18 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.035 $Y=0.98
+ $X2=3.45 $Y2=0.98
r61 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.385 $Y=1.795
+ $X2=3.385 $Y2=2.08
r62 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.385 $Y=1.695 $X2=3.385
+ $Y2=1.795
r63 12 35 192.315 $w=2e-07 $l=5.8e-07 $layer=POLY_cond $X=3.385 $Y=1.695
+ $X2=3.385 $Y2=1.115
r64 9 34 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.36 $Y=0.445 $X2=3.36
+ $Y2=0.845
r65 2 29 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.87 $X2=4.15 $Y2=2.04
r66 1 23 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.15 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_1%X 1 2 10 12 13 14
r16 14 27 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=0.257 $Y=2.21
+ $X2=0.257 $Y2=2.34
r17 13 14 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=1.87
+ $X2=0.257 $Y2=2.21
r18 11 12 46.0977 $w=2.53e-07 $l=1.02e-06 $layer=LI1_cond $X=0.217 $Y=1.495
+ $X2=0.217 $Y2=0.475
r19 10 11 6.36149 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.257 $Y=1.66
+ $X2=0.257 $Y2=1.495
r20 8 13 7.15547 $w=3.33e-07 $l=2.08e-07 $layer=LI1_cond $X=0.257 $Y=1.662
+ $X2=0.257 $Y2=1.87
r21 8 10 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=0.257 $Y=1.662
+ $X2=0.257 $Y2=1.66
r22 2 27 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r23 2 10 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r24 1 12 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_1%VPWR 1 2 11 17 20 21 22 32 33 36
r40 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r42 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r43 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 27 30 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r45 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 26 29 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 24 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.73 $Y2=2.72
r49 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 22 37 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 20 29 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 20 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.67 $Y2=2.72
r53 19 32 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=4.37 $Y2=2.72
r54 19 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.67 $Y2=2.72
r55 15 21 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=2.635
+ $X2=3.67 $Y2=2.72
r56 15 17 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.67 $Y=2.635
+ $X2=3.67 $Y2=2.04
r57 11 14 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.73 $Y=1.66
+ $X2=0.73 $Y2=2.34
r58 9 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635 $X2=0.73
+ $Y2=2.72
r59 9 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.34
r60 2 17 600 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.87 $X2=3.67 $Y2=2.04
r61 1 14 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r62 1 11 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r51 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r52 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r53 33 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r54 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r55 30 39 11.4944 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.507
+ $Y2=0
r56 30 32 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=4.37
+ $Y2=0
r57 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r58 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r59 26 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r60 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r61 25 28 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r62 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r63 23 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r64 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r65 22 39 11.4944 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.507
+ $Y2=0
r66 22 28 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=2.99
+ $Y2=0
r67 17 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r68 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r69 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r70 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r71 11 39 2.14989 $w=5.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.507 $Y=0.085
+ $X2=3.507 $Y2=0
r72 11 13 8.59318 $w=5.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.507 $Y=0.085
+ $X2=3.507 $Y2=0.455
r73 7 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r74 7 9 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.38
r75 2 13 182 $w=1.7e-07 $l=3.37528e-07 $layer=licon1_NDIFF $count=1 $X=3.435
+ $Y=0.235 $X2=3.68 $Y2=0.455
r76 1 9 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

