* File: sky130_fd_sc_hdll__a222oi_1.pex.spice
* Created: Thu Aug 27 18:53:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%C1 1 3 4 6 7 11 13
r24 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.38
+ $Y=1.165 $X2=0.38 $Y2=1.165
r25 7 11 5.12197 $w=3.13e-07 $l=1.4e-07 $layer=LI1_cond $X=0.24 $Y=1.157
+ $X2=0.38 $Y2=1.157
r26 7 13 0.548782 $w=3.13e-07 $l=1.5e-08 $layer=LI1_cond $X=0.24 $Y=1.157
+ $X2=0.225 $Y2=1.157
r27 4 10 40.2858 $w=4.33e-07 $l=2.38642e-07 $layer=POLY_cond $X=0.52 $Y=1
+ $X2=0.35 $Y2=1.165
r28 4 6 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1 $X2=0.52
+ $Y2=0.555
r29 1 10 44.1536 $w=4.33e-07 $l=3.09112e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.35 $Y2=1.165
r30 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%C2 1 3 4 6 7
r25 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.165 $X2=0.94 $Y2=1.165
r26 4 10 47.2445 $w=2.96e-07 $l=2.45e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.165
r27 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r28 1 10 38.5718 $w=2.96e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.88 $Y=1
+ $X2=0.965 $Y2=1.165
r29 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.88 $Y=1 $X2=0.88
+ $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%B2 1 3 4 6 7 15
r26 7 15 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.05 $Y=1.165
+ $X2=2.075 $Y2=1.165
r27 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.05
+ $Y=1.165 $X2=2.05 $Y2=1.165
r28 4 10 38.5876 $w=3.28e-07 $l=2.11069e-07 $layer=POLY_cond $X=2.17 $Y=1
+ $X2=2.065 $Y2=1.165
r29 4 6 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.17 $Y=1 $X2=2.17
+ $Y2=0.555
r30 1 10 45.7447 $w=3.28e-07 $l=2.82179e-07 $layer=POLY_cond $X=2.145 $Y=1.41
+ $X2=2.065 $Y2=1.165
r31 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.145 $Y=1.41
+ $X2=2.145 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%B1 1 3 4 6 7 13
r27 7 13 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=2.555 $Y=1.165
+ $X2=2.545 $Y2=1.165
r28 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.165 $X2=2.59 $Y2=1.165
r29 4 10 49.6426 $w=2.64e-07 $l=2.54804e-07 $layer=POLY_cond $X=2.615 $Y=1.41
+ $X2=2.595 $Y2=1.165
r30 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.615 $Y=1.41
+ $X2=2.615 $Y2=1.985
r31 1 10 39.0383 $w=2.64e-07 $l=1.94808e-07 $layer=POLY_cond $X=2.53 $Y=1
+ $X2=2.595 $Y2=1.165
r32 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.53 $Y=1 $X2=2.53
+ $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%A1 1 3 4 6 7 15
r26 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.165 $X2=3.12 $Y2=1.165
r27 7 15 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.02 $Y=1.165
+ $X2=3.065 $Y2=1.165
r28 4 10 47.2445 $w=2.96e-07 $l=2.73359e-07 $layer=POLY_cond $X=3.085 $Y=1.41
+ $X2=3.145 $Y2=1.165
r29 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.085 $Y=1.41
+ $X2=3.085 $Y2=1.985
r30 1 10 38.5718 $w=2.96e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.06 $Y=1
+ $X2=3.145 $Y2=1.165
r31 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.06 $Y=1 $X2=3.06
+ $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%A2 1 3 4 6 7 15
r22 11 15 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.65 $Y=1.165
+ $X2=3.82 $Y2=1.165
r23 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.65
+ $Y=1.165 $X2=3.65 $Y2=1.165
r24 7 15 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=3.88 $Y=1.165 $X2=3.82
+ $Y2=1.165
r25 4 10 47.2445 $w=2.96e-07 $l=2.73359e-07 $layer=POLY_cond $X=3.615 $Y=1.41
+ $X2=3.675 $Y2=1.165
r26 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.615 $Y=1.41
+ $X2=3.615 $Y2=1.985
r27 1 10 38.5718 $w=2.96e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.59 $Y=1
+ $X2=3.675 $Y2=1.165
r28 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.59 $Y=1 $X2=3.59
+ $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%Y 1 2 3 4 15 19 20 21 25 27 29 30 31 36
+ 43
r62 31 43 2.75204 $w=5.63e-07 $l=1.3e-07 $layer=LI1_cond $X=2.692 $Y=0.51
+ $X2=2.692 $Y2=0.38
r63 29 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=0.51
+ $X2=0.26 $Y2=0.38
r64 28 30 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=1.53 $Y=1.485
+ $X2=1.53 $Y2=1.175
r65 26 30 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=1.53 $Y=0.815
+ $X2=1.53 $Y2=1.175
r66 26 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.53 $Y=0.815
+ $X2=1.53 $Y2=0.73
r67 23 29 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.26 $Y=0.645
+ $X2=0.26 $Y2=0.51
r68 22 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.655 $Y=0.73
+ $X2=1.53 $Y2=0.73
r69 21 31 4.6573 $w=5.63e-07 $l=2.2e-07 $layer=LI1_cond $X=2.692 $Y=0.73
+ $X2=2.692 $Y2=0.51
r70 21 22 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.41 $Y=0.73
+ $X2=1.655 $Y2=0.73
r71 20 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.425 $Y=0.73
+ $X2=0.26 $Y2=0.645
r72 19 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.405 $Y=0.73
+ $X2=1.53 $Y2=0.73
r73 19 20 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=1.405 $Y=0.73
+ $X2=0.425 $Y2=0.73
r74 16 25 3.08873 $w=3.1e-07 $l=1.25e-07 $layer=LI1_cond $X=0.345 $Y=1.64
+ $X2=0.22 $Y2=1.64
r75 16 18 31.7851 $w=3.08e-07 $l=8.55e-07 $layer=LI1_cond $X=0.345 $Y=1.64
+ $X2=1.2 $Y2=1.64
r76 15 28 6.91877 $w=3.1e-07 $l=2.08327e-07 $layer=LI1_cond $X=1.405 $Y=1.64
+ $X2=1.53 $Y2=1.485
r77 15 18 7.62099 $w=3.08e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=1.64
+ $X2=1.2 $Y2=1.64
r78 4 18 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.63
r79 3 25 300 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.765
r80 2 43 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=2.605
+ $Y=0.235 $X2=2.81 $Y2=0.38
r81 1 36 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%A_117_297# 1 2 10 15 16
r22 15 16 10.0337 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.38 $Y=2.3 $X2=2.17
+ $Y2=2.3
r23 10 12 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.73 $Y=2.3 $X2=0.73
+ $Y2=2.38
r24 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.38
+ $X2=0.73 $Y2=2.38
r25 8 16 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=0.895 $Y=2.38
+ $X2=2.17 $Y2=2.38
r26 2 15 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.485 $X2=2.38 $Y2=2.3
r27 1 10 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%A_357_297# 1 2 3 10 16 21 23
r32 17 21 4.66096 $w=2.82e-07 $l=1.47054e-07 $layer=LI1_cond $X=2.935 $Y=1.617
+ $X2=2.81 $Y2=1.665
r33 16 23 3.58503 $w=2.35e-07 $l=1.3e-07 $layer=LI1_cond $X=3.765 $Y=1.617
+ $X2=3.895 $Y2=1.617
r34 16 17 40.7033 $w=2.33e-07 $l=8.3e-07 $layer=LI1_cond $X=3.765 $Y=1.617
+ $X2=2.935 $Y2=1.617
r35 10 21 4.66096 $w=2.82e-07 $l=1.25e-07 $layer=LI1_cond $X=2.685 $Y=1.665
+ $X2=2.81 $Y2=1.665
r36 10 12 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=2.685 $Y=1.665
+ $X2=1.91 $Y2=1.665
r37 3 23 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=3.705
+ $Y=1.485 $X2=3.85 $Y2=1.665
r38 2 21 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=2.705
+ $Y=1.485 $X2=2.85 $Y2=1.665
r39 1 12 600 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=1.785
+ $Y=1.485 $X2=1.91 $Y2=1.665
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%VPWR 1 6 9 10 11 21 22
r41 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r42 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r43 18 19 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 14 18 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 11 19 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 11 14 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r47 9 18 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=2.72
+ $X2=2.99 $Y2=2.72
r48 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=2.72
+ $X2=3.32 $Y2=2.72
r49 8 21 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.91 $Y2=2.72
r50 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.32 $Y2=2.72
r51 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=2.635 $X2=3.32
+ $Y2=2.72
r52 4 6 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=3.32 $Y=2.635 $X2=3.32
+ $Y2=1.99
r53 1 6 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=3.175
+ $Y=1.485 $X2=3.32 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HDLL__A222OI_1%VGND 1 2 7 9 11 18 29 35 38 40
r46 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r47 33 35 8.3097 $w=5.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.61 $Y=0.19
+ $X2=1.705 $Y2=0.19
r48 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r49 31 33 2.82709 $w=5.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.48 $Y=0.19
+ $X2=1.61 $Y2=0.19
r50 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r51 27 31 7.17647 $w=5.48e-07 $l=3.3e-07 $layer=LI1_cond $X=1.15 $Y=0.19
+ $X2=1.48 $Y2=0.19
r52 27 29 11.1368 $w=5.48e-07 $l=2.25e-07 $layer=LI1_cond $X=1.15 $Y=0.19
+ $X2=0.925 $Y2=0.19
r53 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 25 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r55 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r56 22 25 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r57 22 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r58 21 24 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r59 21 35 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.705
+ $Y2=0
r60 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r61 18 37 5.32272 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.847
+ $Y2=0
r62 18 24 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.45
+ $Y2=0
r63 16 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r64 15 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=0.925
+ $Y2=0
r65 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r66 11 16 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r67 11 40 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r68 7 37 3.1353 $w=4.1e-07 $l=1.22327e-07 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.847 $Y2=0
r69 7 9 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.76 $Y=0.085
+ $X2=3.76 $Y2=0.38
r70 2 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.665
+ $Y=0.235 $X2=3.8 $Y2=0.38
r71 1 31 91 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_NDIFF $count=2 $X=0.955
+ $Y=0.235 $X2=1.48 $Y2=0.38
.ends

