* File: sky130_fd_sc_hdll__dfrtp_2.pxi.spice
* Created: Thu Aug 27 19:04:31 2020
* 
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%CLK N_CLK_c_195_n N_CLK_c_199_n N_CLK_c_200_n
+ N_CLK_M1006_g N_CLK_c_196_n N_CLK_M1024_g CLK CLK
+ PM_SKY130_FD_SC_HDLL__DFRTP_2%CLK
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%A_27_47# N_A_27_47#_M1024_s N_A_27_47#_M1006_s
+ N_A_27_47#_c_253_n N_A_27_47#_c_254_n N_A_27_47#_M1027_g N_A_27_47#_M1003_g
+ N_A_27_47#_c_233_n N_A_27_47#_M1015_g N_A_27_47#_c_235_n N_A_27_47#_c_236_n
+ N_A_27_47#_c_257_n N_A_27_47#_c_258_n N_A_27_47#_M1004_g N_A_27_47#_c_259_n
+ N_A_27_47#_c_260_n N_A_27_47#_M1018_g N_A_27_47#_M1020_g N_A_27_47#_c_238_n
+ N_A_27_47#_c_239_n N_A_27_47#_c_240_n N_A_27_47#_c_241_n N_A_27_47#_c_242_n
+ N_A_27_47#_c_262_n N_A_27_47#_c_263_n N_A_27_47#_c_243_n N_A_27_47#_c_244_n
+ N_A_27_47#_c_245_n N_A_27_47#_c_246_n N_A_27_47#_c_247_n N_A_27_47#_c_320_p
+ N_A_27_47#_c_248_n N_A_27_47#_c_249_n N_A_27_47#_c_250_n N_A_27_47#_c_251_n
+ N_A_27_47#_c_252_n PM_SKY130_FD_SC_HDLL__DFRTP_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%D N_D_c_474_n N_D_c_475_n N_D_M1000_g
+ N_D_M1008_g D N_D_c_472_n N_D_c_473_n PM_SKY130_FD_SC_HDLL__DFRTP_2%D
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%A_211_363# N_A_211_363#_M1003_d
+ N_A_211_363#_M1027_d N_A_211_363#_c_530_n N_A_211_363#_M1028_g
+ N_A_211_363#_M1019_g N_A_211_363#_c_523_n N_A_211_363#_M1014_g
+ N_A_211_363#_c_531_n N_A_211_363#_M1029_g N_A_211_363#_c_524_n
+ N_A_211_363#_c_525_n N_A_211_363#_c_526_n N_A_211_363#_c_534_n
+ N_A_211_363#_c_535_n N_A_211_363#_c_527_n N_A_211_363#_c_536_n
+ N_A_211_363#_c_537_n N_A_211_363#_c_538_n N_A_211_363#_c_539_n
+ N_A_211_363#_c_540_n N_A_211_363#_c_528_n N_A_211_363#_c_541_n
+ N_A_211_363#_c_529_n N_A_211_363#_c_543_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_2%A_211_363#
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%A_751_289# N_A_751_289#_M1011_d
+ N_A_751_289#_M1017_d N_A_751_289#_c_739_n N_A_751_289#_M1010_g
+ N_A_751_289#_M1005_g N_A_751_289#_c_741_n N_A_751_289#_c_762_n
+ N_A_751_289#_c_738_n N_A_751_289#_c_764_n N_A_751_289#_c_751_n
+ N_A_751_289#_c_770_n N_A_751_289#_c_754_n N_A_751_289#_c_788_p
+ N_A_751_289#_c_755_n N_A_751_289#_c_743_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_2%A_751_289#
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%RESET_B N_RESET_B_M1007_g N_RESET_B_c_848_n
+ N_RESET_B_c_860_n N_RESET_B_M1023_g N_RESET_B_M1021_g N_RESET_B_c_850_n
+ N_RESET_B_c_862_n N_RESET_B_M1025_g N_RESET_B_c_851_n N_RESET_B_c_852_n
+ N_RESET_B_c_853_n N_RESET_B_c_854_n RESET_B N_RESET_B_c_855_n
+ N_RESET_B_c_856_n N_RESET_B_c_857_n N_RESET_B_c_858_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_2%RESET_B
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%A_534_47# N_A_534_47#_M1015_d
+ N_A_534_47#_M1028_d N_A_534_47#_M1011_g N_A_534_47#_c_995_n
+ N_A_534_47#_c_996_n N_A_534_47#_M1017_g N_A_534_47#_c_1006_n
+ N_A_534_47#_c_1007_n N_A_534_47#_c_997_n N_A_534_47#_c_990_n
+ N_A_534_47#_c_991_n N_A_534_47#_c_992_n N_A_534_47#_c_993_n
+ N_A_534_47#_c_994_n PM_SKY130_FD_SC_HDLL__DFRTP_2%A_534_47#
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%A_1323_21# N_A_1323_21#_M1022_d
+ N_A_1323_21#_M1025_d N_A_1323_21#_M1009_g N_A_1323_21#_c_1118_n
+ N_A_1323_21#_c_1132_n N_A_1323_21#_M1001_g N_A_1323_21#_c_1119_n
+ N_A_1323_21#_M1016_g N_A_1323_21#_c_1133_n N_A_1323_21#_M1002_g
+ N_A_1323_21#_c_1134_n N_A_1323_21#_M1012_g N_A_1323_21#_c_1120_n
+ N_A_1323_21#_M1026_g N_A_1323_21#_c_1121_n N_A_1323_21#_c_1156_n
+ N_A_1323_21#_c_1237_p N_A_1323_21#_c_1202_p N_A_1323_21#_c_1135_n
+ N_A_1323_21#_c_1136_n N_A_1323_21#_c_1122_n N_A_1323_21#_c_1123_n
+ N_A_1323_21#_c_1124_n N_A_1323_21#_c_1125_n N_A_1323_21#_c_1126_n
+ N_A_1323_21#_c_1127_n N_A_1323_21#_c_1128_n N_A_1323_21#_c_1129_n
+ N_A_1323_21#_c_1130_n PM_SKY130_FD_SC_HDLL__DFRTP_2%A_1323_21#
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%A_1128_47# N_A_1128_47#_M1014_d
+ N_A_1128_47#_M1018_d N_A_1128_47#_c_1268_n N_A_1128_47#_M1013_g
+ N_A_1128_47#_M1022_g N_A_1128_47#_c_1275_n N_A_1128_47#_c_1278_n
+ N_A_1128_47#_c_1267_n N_A_1128_47#_c_1270_n N_A_1128_47#_c_1271_n
+ N_A_1128_47#_c_1272_n N_A_1128_47#_c_1273_n N_A_1128_47#_c_1274_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_2%A_1128_47#
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%VPWR N_VPWR_M1006_d N_VPWR_M1000_s
+ N_VPWR_M1010_d N_VPWR_M1017_s N_VPWR_M1001_d N_VPWR_M1013_d N_VPWR_M1002_d
+ N_VPWR_M1012_d N_VPWR_c_1371_n N_VPWR_c_1372_n N_VPWR_c_1373_n N_VPWR_c_1374_n
+ N_VPWR_c_1375_n N_VPWR_c_1376_n N_VPWR_c_1377_n N_VPWR_c_1378_n
+ N_VPWR_c_1379_n N_VPWR_c_1380_n N_VPWR_c_1381_n N_VPWR_c_1382_n
+ N_VPWR_c_1383_n N_VPWR_c_1384_n N_VPWR_c_1385_n N_VPWR_c_1386_n VPWR
+ N_VPWR_c_1387_n N_VPWR_c_1388_n N_VPWR_c_1389_n N_VPWR_c_1390_n
+ N_VPWR_c_1391_n N_VPWR_c_1392_n N_VPWR_c_1393_n N_VPWR_c_1370_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_2%VPWR
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%A_436_413# N_A_436_413#_M1008_d
+ N_A_436_413#_M1000_d N_A_436_413#_c_1526_n N_A_436_413#_c_1534_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_2%A_436_413#
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%A_649_413# N_A_649_413#_M1004_d
+ N_A_649_413#_M1023_d N_A_649_413#_c_1558_n N_A_649_413#_c_1559_n
+ N_A_649_413#_c_1560_n N_A_649_413#_c_1561_n
+ PM_SKY130_FD_SC_HDLL__DFRTP_2%A_649_413#
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%Q N_Q_M1016_d N_Q_M1002_s N_Q_c_1600_n
+ N_Q_c_1601_n Q Q Q Q PM_SKY130_FD_SC_HDLL__DFRTP_2%Q
x_PM_SKY130_FD_SC_HDLL__DFRTP_2%VGND N_VGND_M1024_d N_VGND_M1008_s
+ N_VGND_M1007_d N_VGND_M1009_d N_VGND_M1016_s N_VGND_M1026_s N_VGND_c_1629_n
+ N_VGND_c_1630_n N_VGND_c_1631_n N_VGND_c_1632_n N_VGND_c_1633_n
+ N_VGND_c_1634_n N_VGND_c_1635_n N_VGND_c_1636_n N_VGND_c_1637_n
+ N_VGND_c_1638_n N_VGND_c_1639_n VGND N_VGND_c_1640_n N_VGND_c_1641_n
+ N_VGND_c_1642_n N_VGND_c_1643_n N_VGND_c_1644_n N_VGND_c_1645_n
+ N_VGND_c_1646_n PM_SKY130_FD_SC_HDLL__DFRTP_2%VGND
cc_1 VNB N_CLK_c_195_n 0.0612188f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.325
cc_2 VNB N_CLK_c_196_n 0.0173562f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_3 VNB CLK 0.0160726f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_27_47#_M1003_g 0.0398926f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_5 VNB N_A_27_47#_c_233_n 0.00940056f $X=-0.19 $Y=-0.24 $X2=0.352 $Y2=1.16
cc_6 VNB N_A_27_47#_M1015_g 0.0216328f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_7 VNB N_A_27_47#_c_235_n 0.0166446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_236_n 0.00209111f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_9 VNB N_A_27_47#_M1020_g 0.0295774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_238_n 0.00876829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_239_n 0.0122713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_240_n 0.0111414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_241_n 0.00233121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_242_n 0.00783792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_243_n 0.0241996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_244_n 0.00242452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_245_n 0.0304994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_246_n 0.00143056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_247_n 0.00705679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_248_n 0.0128491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_249_n 0.00850994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_250_n 0.0267639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_251_n 0.0243368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_252_n 0.00481911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_D_M1008_g 0.0473066f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_26 VNB N_D_c_472_n 0.0175222f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_27 VNB N_D_c_473_n 0.0117199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_211_363#_M1019_g 0.0242299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_211_363#_c_523_n 0.0181936f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_30 VNB N_A_211_363#_c_524_n 0.00301844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_211_363#_c_525_n 0.00523438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_211_363#_c_526_n 0.0373752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_211_363#_c_527_n 0.00348148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_211_363#_c_528_n 0.0280171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_211_363#_c_529_n 0.0129087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_751_289#_M1005_g 0.0473898f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_751_289#_c_738_n 0.0068767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_RESET_B_c_848_n 0.010178f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_39 VNB N_RESET_B_M1021_g 0.03034f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_40 VNB N_RESET_B_c_850_n 0.00107309f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_41 VNB N_RESET_B_c_851_n 0.00475244f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_42 VNB N_RESET_B_c_852_n 0.0126778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_RESET_B_c_853_n 0.0239364f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_44 VNB N_RESET_B_c_854_n 0.00118946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_c_855_n 0.0287326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_RESET_B_c_856_n 0.0180244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_857_n 0.0255139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_RESET_B_c_858_n 0.0109903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_534_47#_M1011_g 0.0198132f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_50 VNB N_A_534_47#_c_990_n 0.0122396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_534_47#_c_991_n 0.00579517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_534_47#_c_992_n 0.00381677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_534_47#_c_993_n 0.00185456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_534_47#_c_994_n 0.03171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1323_21#_M1009_g 0.0235966f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_56 VNB N_A_1323_21#_c_1118_n 0.0119026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1323_21#_c_1119_n 0.020444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1323_21#_c_1120_n 0.020726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1323_21#_c_1121_n 0.00212051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1323_21#_c_1122_n 0.00309251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1323_21#_c_1123_n 0.0145092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1323_21#_c_1124_n 2.46176e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1323_21#_c_1125_n 0.021055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1323_21#_c_1126_n 6.38325e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1323_21#_c_1127_n 0.00574148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1323_21#_c_1128_n 0.00784546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1323_21#_c_1129_n 0.0560539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1323_21#_c_1130_n 0.0443114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1128_47#_M1022_g 0.0509803f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1128_47#_c_1267_n 0.0075193f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_71 VNB N_VPWR_c_1370_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_436_413#_c_1526_n 0.00396469f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_73 VNB Q 0.0301873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1629_n 0.0197352f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_75 VNB N_VGND_c_1630_n 0.0083472f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_76 VNB N_VGND_c_1631_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1632_n 0.00469188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1633_n 0.00647875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1634_n 0.0114954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1635_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1636_n 0.0495892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1637_n 0.00323844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1638_n 0.0442527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1639_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1640_n 0.014742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1641_n 0.0720206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1642_n 0.0199439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1643_n 0.0085923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1644_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1645_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1646_n 0.482071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VPB N_CLK_c_195_n 0.00482568f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.325
cc_93 VPB N_CLK_c_199_n 0.014844f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_94 VPB N_CLK_c_200_n 0.0466088f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_95 VPB CLK 0.0154183f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_96 VPB N_A_27_47#_c_253_n 0.018961f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_97 VPB N_A_27_47#_c_254_n 0.025741f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_98 VPB N_A_27_47#_c_235_n 0.0167098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_27_47#_c_236_n 0.0066803f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_100 VPB N_A_27_47#_c_257_n 0.029683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_27_47#_c_258_n 0.0247481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_27_47#_c_259_n 0.0295268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_27_47#_c_260_n 0.0241122f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_27_47#_c_238_n 0.0127828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_47#_c_262_n 0.00133165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_27_47#_c_263_n 0.0297432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_27_47#_c_244_n 4.26143e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_27_47#_c_247_n 0.00369171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_27_47#_c_249_n 2.26672e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_27_47#_c_250_n 0.0124295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_252_n 6.80124e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_D_c_474_n 0.0154669f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_113 VPB N_D_c_475_n 0.0279937f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_114 VPB D 0.0110956f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_115 VPB N_D_c_472_n 0.00480826f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_116 VPB N_D_c_473_n 0.0413087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_211_363#_c_530_n 0.0530318f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_118 VPB N_A_211_363#_c_531_n 0.0547481f $X=-0.19 $Y=1.305 $X2=0.352 $Y2=1.16
cc_119 VPB N_A_211_363#_c_524_n 0.00372121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_211_363#_c_525_n 0.00412205f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_211_363#_c_534_n 0.00249202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_211_363#_c_535_n 0.00178621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_211_363#_c_536_n 0.0100109f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_211_363#_c_537_n 0.00230751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_211_363#_c_538_n 0.0163244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_211_363#_c_539_n 0.00140509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_211_363#_c_540_n 0.00284223f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_211_363#_c_541_n 0.00955918f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_211_363#_c_529_n 0.0113234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_211_363#_c_543_n 0.00625748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_751_289#_c_739_n 0.0620472f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_132 VPB N_A_751_289#_M1005_g 0.00822468f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_751_289#_c_741_n 0.013925f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_134 VPB N_A_751_289#_c_738_n 0.00189073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_751_289#_c_743_n 5.23824e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_RESET_B_c_848_n 0.0368117f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_137 VPB N_RESET_B_c_860_n 0.0266961f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_138 VPB N_RESET_B_c_850_n 0.0350735f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_139 VPB N_RESET_B_c_862_n 0.0251347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_RESET_B_c_858_n 0.00382208f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_534_47#_c_995_n 0.0300431f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_142 VPB N_A_534_47#_c_996_n 0.0188583f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_143 VPB N_A_534_47#_c_997_n 0.00699003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_534_47#_c_991_n 0.00744183f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_534_47#_c_992_n 0.00396196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_534_47#_c_993_n 0.00113493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_534_47#_c_994_n 0.0256017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_1323_21#_c_1118_n 0.0375913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_1323_21#_c_1132_n 0.0235314f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_150 VPB N_A_1323_21#_c_1133_n 0.0195301f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_151 VPB N_A_1323_21#_c_1134_n 0.0194452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_1323_21#_c_1135_n 0.00709871f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_1323_21#_c_1136_n 0.00336491f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_1323_21#_c_1124_n 0.0146808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_1323_21#_c_1130_n 0.0223386f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_1128_47#_c_1268_n 0.0598568f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_157 VPB N_A_1128_47#_M1022_g 0.0112371f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_1128_47#_c_1270_n 0.0037881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_1128_47#_c_1271_n 0.00376023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_1128_47#_c_1272_n 0.00187849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_1128_47#_c_1273_n 0.0341344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_1128_47#_c_1274_n 0.00364602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1371_n 0.00126291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1372_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1373_n 0.00286019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1374_n 0.00785764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1375_n 0.00234526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1376_n 0.00824014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1377_n 0.00356354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1378_n 0.0118247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1379_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1380_n 0.0241628f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1381_n 0.0032427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1382_n 0.0525704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1383_n 0.00513379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1384_n 0.0480155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1385_n 0.00359728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1386_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1387_n 0.0146985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1388_n 0.0184687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1389_n 0.0138694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1390_n 0.0216041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1391_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1392_n 0.0067475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1393_n 0.00960541f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1370_n 0.0665812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_436_413#_c_1526_n 0.00787003f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.445
cc_188 VPB N_A_649_413#_c_1558_n 4.90981e-19 $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_189 VPB N_A_649_413#_c_1559_n 0.00902117f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.665
cc_190 VPB N_A_649_413#_c_1560_n 0.00246066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_649_413#_c_1561_n 7.36897e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB Q 0.00732327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB Q 0.0121091f $X=-0.19 $Y=1.305 $X2=0.352 $Y2=1.16
cc_194 N_CLK_c_199_n N_A_27_47#_c_253_n 0.00262901f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_195 N_CLK_c_200_n N_A_27_47#_c_253_n 0.00668506f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_196 CLK N_A_27_47#_c_253_n 8.03089e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_197 N_CLK_c_200_n N_A_27_47#_c_254_n 0.0192779f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_198 N_CLK_c_195_n N_A_27_47#_M1003_g 0.00192687f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_199 N_CLK_c_196_n N_A_27_47#_M1003_g 0.0154184f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_200 N_CLK_c_195_n N_A_27_47#_c_241_n 0.0108877f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_201 N_CLK_c_196_n N_A_27_47#_c_241_n 0.00652815f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_202 CLK N_A_27_47#_c_241_n 0.00736322f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_203 N_CLK_c_195_n N_A_27_47#_c_242_n 0.0070116f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_204 CLK N_A_27_47#_c_242_n 0.0220292f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_205 N_CLK_c_200_n N_A_27_47#_c_262_n 0.0171402f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_206 CLK N_A_27_47#_c_262_n 0.00731943f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_207 N_CLK_c_195_n N_A_27_47#_c_263_n 4.93713e-19 $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_208 N_CLK_c_200_n N_A_27_47#_c_263_n 0.00841026f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_209 CLK N_A_27_47#_c_263_n 0.0231715f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_210 CLK N_A_27_47#_c_244_n 0.00762548f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_211 N_CLK_c_195_n N_A_27_47#_c_247_n 0.0029245f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_212 N_CLK_c_199_n N_A_27_47#_c_247_n 4.50807e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_213 N_CLK_c_200_n N_A_27_47#_c_247_n 0.00460739f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_214 CLK N_A_27_47#_c_247_n 0.0396442f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_215 N_CLK_c_195_n N_A_27_47#_c_250_n 0.0139997f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_216 CLK N_A_27_47#_c_250_n 0.00161375f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_217 N_CLK_c_200_n N_VPWR_c_1371_n 0.0125197f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_218 N_CLK_c_200_n N_VPWR_c_1387_n 0.00304525f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_219 N_CLK_c_200_n N_VPWR_c_1370_n 0.00454898f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_220 N_CLK_c_195_n N_VGND_c_1640_n 6.41851e-19 $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_221 N_CLK_c_196_n N_VGND_c_1640_n 0.00198377f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_222 N_CLK_c_196_n N_VGND_c_1643_n 0.0142867f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_223 N_CLK_c_196_n N_VGND_c_1646_n 0.00367064f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_233_n N_D_M1008_g 0.0069239f $X=2.567 $Y=1.245 $X2=0 $Y2=0
cc_225 N_A_27_47#_M1015_g N_D_M1008_g 0.0114163f $X=2.595 $Y=0.415 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_243_n N_D_M1008_g 0.00433004f $X=2.42 $Y=1.19 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_251_n N_D_M1008_g 0.0202027f $X=2.535 $Y=0.93 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_252_n N_D_M1008_g 0.00110511f $X=2.535 $Y=0.93 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_243_n N_D_c_472_n 0.0442169f $X=2.42 $Y=1.19 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_236_n N_D_c_473_n 0.0069239f $X=2.67 $Y=1.32 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_243_n N_D_c_473_n 0.00279795f $X=2.42 $Y=1.19 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_250_n N_D_c_473_n 0.00387403f $X=0.99 $Y=1.235 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_236_n N_A_211_363#_c_530_n 0.0220389f $X=2.67 $Y=1.32 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_257_n N_A_211_363#_c_530_n 0.0178804f $X=3.155 $Y=1.89 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_258_n N_A_211_363#_c_530_n 0.0156562f $X=3.155 $Y=1.99 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_251_n N_A_211_363#_c_530_n 6.13774e-19 $X=2.535 $Y=0.93
+ $X2=0 $Y2=0
cc_237 N_A_27_47#_c_252_n N_A_211_363#_c_530_n 0.00148383f $X=2.535 $Y=0.93
+ $X2=0 $Y2=0
cc_238 N_A_27_47#_M1015_g N_A_211_363#_M1019_g 0.0170554f $X=2.595 $Y=0.415
+ $X2=0 $Y2=0
cc_239 N_A_27_47#_M1020_g N_A_211_363#_c_523_n 0.0133187f $X=6.11 $Y=0.415 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_259_n N_A_211_363#_c_531_n 0.0187963f $X=6.02 $Y=1.89 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_260_n N_A_211_363#_c_531_n 0.0193363f $X=6.02 $Y=1.99 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_235_n N_A_211_363#_c_524_n 0.0110718f $X=3.055 $Y=1.32 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_257_n N_A_211_363#_c_524_n 0.00429121f $X=3.155 $Y=1.89
+ $X2=0 $Y2=0
cc_244 N_A_27_47#_c_245_n N_A_211_363#_c_524_n 0.0112341f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_246_n N_A_211_363#_c_524_n 0.00245105f $X=2.71 $Y=1.19 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_251_n N_A_211_363#_c_524_n 0.00150259f $X=2.535 $Y=0.93
+ $X2=0 $Y2=0
cc_247 N_A_27_47#_c_252_n N_A_211_363#_c_524_n 0.0281131f $X=2.535 $Y=0.93 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_M1020_g N_A_211_363#_c_525_n 3.86971e-19 $X=6.11 $Y=0.415
+ $X2=0 $Y2=0
cc_249 N_A_27_47#_c_238_n N_A_211_363#_c_525_n 0.0071137f $X=6.112 $Y=1.395
+ $X2=0 $Y2=0
cc_250 N_A_27_47#_c_239_n N_A_211_363#_c_525_n 0.00110845f $X=6.17 $Y=1.08 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_245_n N_A_211_363#_c_525_n 0.0128498f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_320_p N_A_211_363#_c_525_n 6.5357e-19 $X=6.105 $Y=1.19 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_249_n N_A_211_363#_c_525_n 0.0451388f $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_M1020_g N_A_211_363#_c_526_n 0.021218f $X=6.11 $Y=0.415 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_245_n N_A_211_363#_c_526_n 0.00202654f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_249_n N_A_211_363#_c_526_n 0.00186694f $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_259_n N_A_211_363#_c_534_n 0.013719f $X=6.02 $Y=1.89 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_238_n N_A_211_363#_c_534_n 7.12282e-19 $X=6.112 $Y=1.395
+ $X2=0 $Y2=0
cc_259 N_A_27_47#_c_245_n N_A_211_363#_c_534_n 0.00477835f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_320_p N_A_211_363#_c_534_n 7.00605e-19 $X=6.105 $Y=1.19
+ $X2=0 $Y2=0
cc_261 N_A_27_47#_c_249_n N_A_211_363#_c_534_n 0.0132445f $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_235_n N_A_211_363#_c_527_n 0.00115186f $X=3.055 $Y=1.32
+ $X2=0 $Y2=0
cc_263 N_A_27_47#_c_245_n N_A_211_363#_c_527_n 0.00894827f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_251_n N_A_211_363#_c_527_n 7.0175e-19 $X=2.535 $Y=0.93 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_252_n N_A_211_363#_c_527_n 0.0180079f $X=2.535 $Y=0.93 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_243_n N_A_211_363#_c_536_n 0.0464444f $X=2.42 $Y=1.19 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_246_n N_A_211_363#_c_536_n 0.0107245f $X=2.71 $Y=1.19 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_252_n N_A_211_363#_c_536_n 0.00257362f $X=2.535 $Y=0.93
+ $X2=0 $Y2=0
cc_269 N_A_27_47#_c_254_n N_A_211_363#_c_537_n 0.00479165f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_270 N_A_27_47#_c_262_n N_A_211_363#_c_537_n 0.00546643f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_243_n N_A_211_363#_c_537_n 0.0161767f $X=2.42 $Y=1.19 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_247_n N_A_211_363#_c_537_n 0.00111166f $X=0.745 $Y=1.19
+ $X2=0 $Y2=0
cc_273 N_A_27_47#_c_235_n N_A_211_363#_c_538_n 3.59761e-19 $X=3.055 $Y=1.32
+ $X2=0 $Y2=0
cc_274 N_A_27_47#_c_257_n N_A_211_363#_c_538_n 0.00285737f $X=3.155 $Y=1.89
+ $X2=0 $Y2=0
cc_275 N_A_27_47#_c_258_n N_A_211_363#_c_538_n 0.00164817f $X=3.155 $Y=1.99
+ $X2=0 $Y2=0
cc_276 N_A_27_47#_c_259_n N_A_211_363#_c_538_n 0.00335603f $X=6.02 $Y=1.89 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_260_n N_A_211_363#_c_538_n 0.00369059f $X=6.02 $Y=1.99 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_245_n N_A_211_363#_c_538_n 0.129135f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_320_p N_A_211_363#_c_538_n 0.0129049f $X=6.105 $Y=1.19 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_249_n N_A_211_363#_c_538_n 5.22408e-19 $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_258_n N_A_211_363#_c_539_n 3.51991e-19 $X=3.155 $Y=1.99
+ $X2=0 $Y2=0
cc_282 N_A_27_47#_c_245_n N_A_211_363#_c_539_n 0.0108696f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_246_n N_A_211_363#_c_539_n 0.00221839f $X=2.71 $Y=1.19 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_260_n N_A_211_363#_c_540_n 4.36466e-19 $X=6.02 $Y=1.99 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_235_n N_A_211_363#_c_528_n 0.0230522f $X=3.055 $Y=1.32 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_245_n N_A_211_363#_c_528_n 0.0025822f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_251_n N_A_211_363#_c_528_n 0.0175107f $X=2.535 $Y=0.93 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_252_n N_A_211_363#_c_528_n 7.93384e-19 $X=2.535 $Y=0.93
+ $X2=0 $Y2=0
cc_289 N_A_27_47#_c_259_n N_A_211_363#_c_541_n 0.00599608f $X=6.02 $Y=1.89 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_238_n N_A_211_363#_c_541_n 0.00436301f $X=6.112 $Y=1.395
+ $X2=0 $Y2=0
cc_291 N_A_27_47#_c_320_p N_A_211_363#_c_541_n 5.03987e-19 $X=6.105 $Y=1.19
+ $X2=0 $Y2=0
cc_292 N_A_27_47#_c_249_n N_A_211_363#_c_541_n 0.0130457f $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_254_n N_A_211_363#_c_529_n 0.0065704f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_M1003_g N_A_211_363#_c_529_n 0.0217374f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_241_n N_A_211_363#_c_529_n 0.0103201f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_262_n N_A_211_363#_c_529_n 0.00841124f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_243_n N_A_211_363#_c_529_n 0.0193232f $X=2.42 $Y=1.19 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_244_n N_A_211_363#_c_529_n 0.00224499f $X=0.89 $Y=1.19 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_247_n N_A_211_363#_c_529_n 0.0568565f $X=0.745 $Y=1.19 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_235_n N_A_211_363#_c_543_n 8.09221e-19 $X=3.055 $Y=1.32
+ $X2=0 $Y2=0
cc_301 N_A_27_47#_c_236_n N_A_211_363#_c_543_n 0.00575298f $X=2.67 $Y=1.32 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_257_n N_A_211_363#_c_543_n 0.00348747f $X=3.155 $Y=1.89
+ $X2=0 $Y2=0
cc_303 N_A_27_47#_c_245_n N_A_211_363#_c_543_n 0.0042506f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_246_n N_A_211_363#_c_543_n 0.00149973f $X=2.71 $Y=1.19 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_252_n N_A_211_363#_c_543_n 0.0114129f $X=2.535 $Y=0.93 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_257_n N_A_751_289#_c_739_n 0.0107188f $X=3.155 $Y=1.89 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_258_n N_A_751_289#_c_739_n 0.00903797f $X=3.155 $Y=1.99
+ $X2=0 $Y2=0
cc_308 N_A_27_47#_c_235_n N_A_751_289#_M1005_g 0.00258973f $X=3.055 $Y=1.32
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_c_245_n N_A_751_289#_M1005_g 0.00261559f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_257_n N_A_751_289#_c_741_n 6.92247e-19 $X=3.155 $Y=1.89
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_c_245_n N_A_751_289#_c_741_n 0.00817769f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_245_n N_A_751_289#_c_738_n 0.0134253f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_259_n N_A_751_289#_c_751_n 0.00211497f $X=6.02 $Y=1.89 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_260_n N_A_751_289#_c_751_n 4.46283e-19 $X=6.02 $Y=1.99 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_245_n N_A_751_289#_c_751_n 0.00274109f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_260_n N_A_751_289#_c_754_n 0.00558596f $X=6.02 $Y=1.99 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_245_n N_A_751_289#_c_755_n 0.00116222f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_245_n N_RESET_B_c_848_n 0.00186512f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_245_n N_RESET_B_c_851_n 0.0683084f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_245_n N_RESET_B_c_852_n 0.00859934f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_245_n N_RESET_B_c_853_n 0.0965654f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_320_p N_RESET_B_c_853_n 0.0249445f $X=6.105 $Y=1.19 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_249_n N_RESET_B_c_853_n 0.0195295f $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_245_n N_RESET_B_c_855_n 0.00219045f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_259_n N_A_534_47#_c_995_n 0.00471069f $X=6.02 $Y=1.89 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_245_n N_A_534_47#_c_995_n 0.00392735f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_259_n N_A_534_47#_c_996_n 0.0138529f $X=6.02 $Y=1.89 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_260_n N_A_534_47#_c_996_n 0.0125159f $X=6.02 $Y=1.99 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_258_n N_A_534_47#_c_1006_n 0.0176799f $X=3.155 $Y=1.99 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_246_n N_A_534_47#_c_1007_n 4.77127e-19 $X=2.71 $Y=1.19 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_235_n N_A_534_47#_c_997_n 0.00143343f $X=3.055 $Y=1.32 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_257_n N_A_534_47#_c_997_n 0.0118934f $X=3.155 $Y=1.89 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_258_n N_A_534_47#_c_997_n 0.00704505f $X=3.155 $Y=1.99 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_245_n N_A_534_47#_c_997_n 4.47339e-19 $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_245_n N_A_534_47#_c_990_n 0.0136728f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_245_n N_A_534_47#_c_991_n 0.0392271f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_235_n N_A_534_47#_c_992_n 0.00519898f $X=3.055 $Y=1.32 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_245_n N_A_534_47#_c_992_n 0.0158094f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_245_n N_A_534_47#_c_993_n 0.0100049f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_245_n N_A_534_47#_c_994_n 0.00541754f $X=5.96 $Y=1.19 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_M1020_g N_A_1323_21#_M1009_g 0.021318f $X=6.11 $Y=0.415 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_249_n N_A_1323_21#_M1009_g 6.57524e-19 $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_248_n N_A_1323_21#_c_1118_n 0.0031393f $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_239_n N_A_1323_21#_c_1129_n 0.00393729f $X=6.17 $Y=1.08
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_M1020_g N_A_1128_47#_c_1275_n 0.0116653f $X=6.11 $Y=0.415
+ $X2=0 $Y2=0
cc_346 N_A_27_47#_c_239_n N_A_1128_47#_c_1275_n 4.18304e-19 $X=6.17 $Y=1.08
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_c_249_n N_A_1128_47#_c_1275_n 0.0230263f $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_260_n N_A_1128_47#_c_1278_n 0.00711942f $X=6.02 $Y=1.99
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_M1020_g N_A_1128_47#_c_1267_n 0.00375536f $X=6.11 $Y=0.415
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_239_n N_A_1128_47#_c_1267_n 0.00139891f $X=6.17 $Y=1.08
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_320_p N_A_1128_47#_c_1267_n 0.00142991f $X=6.105 $Y=1.19
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_c_249_n N_A_1128_47#_c_1267_n 0.046143f $X=6.17 $Y=1.11 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_259_n N_A_1128_47#_c_1271_n 0.00281119f $X=6.02 $Y=1.89
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_238_n N_A_1128_47#_c_1271_n 0.00198112f $X=6.112 $Y=1.395
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_c_249_n N_A_1128_47#_c_1271_n 8.51835e-19 $X=6.17 $Y=1.11
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_c_262_n N_VPWR_M1006_d 0.001889f $X=0.66 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_357 N_A_27_47#_c_254_n N_VPWR_c_1371_n 0.00960497f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_262_n N_VPWR_c_1371_n 0.0213487f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_359 N_A_27_47#_c_263_n N_VPWR_c_1371_n 0.0254007f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_360 N_A_27_47#_c_260_n N_VPWR_c_1374_n 0.00107286f $X=6.02 $Y=1.99 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_254_n N_VPWR_c_1380_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_258_n N_VPWR_c_1382_n 0.00431663f $X=3.155 $Y=1.99 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_260_n N_VPWR_c_1384_n 0.00632161f $X=6.02 $Y=1.99 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_262_n N_VPWR_c_1387_n 0.00180073f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_263_n N_VPWR_c_1387_n 0.0181185f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_366 N_A_27_47#_c_254_n N_VPWR_c_1370_n 0.00986661f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_258_n N_VPWR_c_1370_n 0.00673557f $X=3.155 $Y=1.99 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_260_n N_VPWR_c_1370_n 0.00754494f $X=6.02 $Y=1.99 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_262_n N_VPWR_c_1370_n 0.00528325f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_263_n N_VPWR_c_1370_n 0.00973967f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_233_n N_A_436_413#_c_1526_n 7.60354e-19 $X=2.567 $Y=1.245
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_M1015_g N_A_436_413#_c_1526_n 0.00225592f $X=2.595 $Y=0.415
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_243_n N_A_436_413#_c_1526_n 0.0196961f $X=2.42 $Y=1.19 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_246_n N_A_436_413#_c_1526_n 0.00249824f $X=2.71 $Y=1.19
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_251_n N_A_436_413#_c_1526_n 0.00178642f $X=2.535 $Y=0.93
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_252_n N_A_436_413#_c_1526_n 0.0428455f $X=2.535 $Y=0.93
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_246_n N_A_436_413#_c_1534_n 4.58473e-19 $X=2.71 $Y=1.19
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_251_n N_A_436_413#_c_1534_n 0.00120163f $X=2.535 $Y=0.93
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_252_n N_A_436_413#_c_1534_n 0.00225275f $X=2.535 $Y=0.93
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_258_n N_A_649_413#_c_1558_n 9.58523e-19 $X=3.155 $Y=1.99
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_245_n N_A_649_413#_c_1559_n 3.42555e-19 $X=5.96 $Y=1.19
+ $X2=0 $Y2=0
cc_382 N_A_27_47#_c_257_n N_A_649_413#_c_1560_n 3.72601e-19 $X=3.155 $Y=1.89
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_c_241_n N_VGND_M1024_d 0.00227127f $X=0.66 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_384 N_A_27_47#_M1003_g N_VGND_c_1629_n 0.00585385f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_M1003_g N_VGND_c_1630_n 0.0046934f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_M1020_g N_VGND_c_1636_n 0.00357877f $X=6.11 $Y=0.415 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_240_n N_VGND_c_1640_n 0.0109767f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_388 N_A_27_47#_c_241_n N_VGND_c_1640_n 0.00244154f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_M1015_g N_VGND_c_1641_n 0.00585385f $X=2.595 $Y=0.415 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_251_n N_VGND_c_1641_n 2.22902e-19 $X=2.535 $Y=0.93 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_M1003_g N_VGND_c_1643_n 0.00317372f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_240_n N_VGND_c_1643_n 0.00923148f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_241_n N_VGND_c_1643_n 0.0224548f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_394 N_A_27_47#_c_244_n N_VGND_c_1643_n 9.39106e-19 $X=0.89 $Y=1.19 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_c_250_n N_VGND_c_1643_n 6.78636e-19 $X=0.99 $Y=1.235 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_M1024_s N_VGND_c_1646_n 0.00296179f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_M1003_g N_VGND_c_1646_n 0.0120602f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_M1015_g N_VGND_c_1646_n 0.00656718f $X=2.595 $Y=0.415 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_M1020_g N_VGND_c_1646_n 0.00586124f $X=6.11 $Y=0.415 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_240_n N_VGND_c_1646_n 0.00916732f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_241_n N_VGND_c_1646_n 0.00625251f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_252_n N_VGND_c_1646_n 0.00669148f $X=2.535 $Y=0.93 $X2=0
+ $Y2=0
cc_403 N_D_c_474_n N_A_211_363#_c_530_n 0.00426071f $X=2.09 $Y=1.89 $X2=0 $Y2=0
cc_404 N_D_c_475_n N_A_211_363#_c_530_n 0.00889704f $X=2.09 $Y=1.99 $X2=0 $Y2=0
cc_405 N_D_c_473_n N_A_211_363#_c_530_n 0.0147096f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_406 N_D_c_473_n N_A_211_363#_c_524_n 8.60547e-19 $X=2.115 $Y=1.465 $X2=0
+ $Y2=0
cc_407 N_D_c_474_n N_A_211_363#_c_536_n 0.00272445f $X=2.09 $Y=1.89 $X2=0 $Y2=0
cc_408 N_D_c_475_n N_A_211_363#_c_536_n 0.00214948f $X=2.09 $Y=1.99 $X2=0 $Y2=0
cc_409 D N_A_211_363#_c_536_n 0.0230339f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_410 N_D_c_472_n N_A_211_363#_c_536_n 0.00255825f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_411 N_D_c_473_n N_A_211_363#_c_536_n 0.00149021f $X=2.115 $Y=1.465 $X2=0
+ $Y2=0
cc_412 D N_A_211_363#_c_537_n 0.00286939f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_413 N_D_c_472_n N_A_211_363#_c_529_n 0.10825f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_414 N_D_c_473_n N_A_211_363#_c_529_n 7.67912e-19 $X=2.115 $Y=1.465 $X2=0
+ $Y2=0
cc_415 N_D_c_473_n N_A_211_363#_c_543_n 5.04388e-19 $X=2.115 $Y=1.465 $X2=0
+ $Y2=0
cc_416 N_D_c_475_n N_VPWR_c_1372_n 0.00574486f $X=2.09 $Y=1.99 $X2=0 $Y2=0
cc_417 N_D_c_472_n N_VPWR_c_1372_n 0.00239948f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_418 N_D_c_473_n N_VPWR_c_1372_n 0.00185248f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_419 D N_VPWR_c_1380_n 0.00542885f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_420 N_D_c_475_n N_VPWR_c_1382_n 0.0061573f $X=2.09 $Y=1.99 $X2=0 $Y2=0
cc_421 N_D_c_475_n N_VPWR_c_1370_n 0.00837936f $X=2.09 $Y=1.99 $X2=0 $Y2=0
cc_422 D N_VPWR_c_1370_n 0.00410324f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_423 N_D_c_474_n N_A_436_413#_c_1526_n 0.00612884f $X=2.09 $Y=1.89 $X2=0 $Y2=0
cc_424 N_D_c_475_n N_A_436_413#_c_1526_n 0.0169987f $X=2.09 $Y=1.99 $X2=0 $Y2=0
cc_425 N_D_M1008_g N_A_436_413#_c_1526_n 0.0210981f $X=2.115 $Y=0.445 $X2=0
+ $Y2=0
cc_426 D N_A_436_413#_c_1526_n 0.0149603f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_427 N_D_c_472_n N_A_436_413#_c_1526_n 0.0783188f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_428 N_D_c_473_n N_A_436_413#_c_1526_n 0.0117503f $X=2.115 $Y=1.465 $X2=0
+ $Y2=0
cc_429 N_D_M1008_g N_A_436_413#_c_1534_n 0.00540291f $X=2.115 $Y=0.445 $X2=0
+ $Y2=0
cc_430 N_D_c_472_n N_VGND_M1008_s 0.00428207f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_431 N_D_c_472_n N_VGND_c_1629_n 0.0025095f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_432 N_D_M1008_g N_VGND_c_1630_n 0.00942073f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_433 N_D_c_472_n N_VGND_c_1630_n 0.0275242f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_434 N_D_M1008_g N_VGND_c_1641_n 0.00418817f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_435 N_D_M1008_g N_VGND_c_1646_n 0.00807145f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_436 N_D_c_472_n N_VGND_c_1646_n 0.00539668f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_437 N_A_211_363#_c_534_n N_A_751_289#_M1017_d 7.49776e-19 $X=6.145 $Y=1.58
+ $X2=0 $Y2=0
cc_438 N_A_211_363#_c_535_n N_A_751_289#_M1017_d 0.00159488f $X=5.775 $Y=1.58
+ $X2=0 $Y2=0
cc_439 N_A_211_363#_c_538_n N_A_751_289#_M1017_d 0.00261316f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_440 N_A_211_363#_c_538_n N_A_751_289#_c_739_n 0.00533159f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_441 N_A_211_363#_M1019_g N_A_751_289#_M1005_g 0.0112388f $X=3.135 $Y=0.415
+ $X2=0 $Y2=0
cc_442 N_A_211_363#_c_538_n N_A_751_289#_c_741_n 0.0234027f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_443 N_A_211_363#_c_523_n N_A_751_289#_c_762_n 0.00342606f $X=5.565 $Y=0.705
+ $X2=0 $Y2=0
cc_444 N_A_211_363#_c_535_n N_A_751_289#_c_738_n 0.00165359f $X=5.775 $Y=1.58
+ $X2=0 $Y2=0
cc_445 N_A_211_363#_c_538_n N_A_751_289#_c_764_n 0.00739158f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_446 N_A_211_363#_c_534_n N_A_751_289#_c_751_n 0.00255823f $X=6.145 $Y=1.58
+ $X2=0 $Y2=0
cc_447 N_A_211_363#_c_535_n N_A_751_289#_c_751_n 0.0112322f $X=5.775 $Y=1.58
+ $X2=0 $Y2=0
cc_448 N_A_211_363#_c_538_n N_A_751_289#_c_751_n 0.0226052f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_449 N_A_211_363#_c_540_n N_A_751_289#_c_751_n 0.00120279f $X=6.555 $Y=1.87
+ $X2=0 $Y2=0
cc_450 N_A_211_363#_c_541_n N_A_751_289#_c_751_n 0.00459528f $X=6.495 $Y=1.74
+ $X2=0 $Y2=0
cc_451 N_A_211_363#_c_538_n N_A_751_289#_c_770_n 0.00696959f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_452 N_A_211_363#_c_525_n N_A_751_289#_c_755_n 0.0376406f $X=5.69 $Y=0.87
+ $X2=0 $Y2=0
cc_453 N_A_211_363#_c_526_n N_A_751_289#_c_755_n 0.00342606f $X=5.69 $Y=0.87
+ $X2=0 $Y2=0
cc_454 N_A_211_363#_c_535_n N_A_751_289#_c_743_n 0.00831119f $X=5.775 $Y=1.58
+ $X2=0 $Y2=0
cc_455 N_A_211_363#_c_538_n N_RESET_B_c_848_n 0.00331104f $X=6.41 $Y=1.87 $X2=0
+ $Y2=0
cc_456 N_A_211_363#_c_525_n N_RESET_B_c_853_n 0.0114823f $X=5.69 $Y=0.87 $X2=0
+ $Y2=0
cc_457 N_A_211_363#_c_526_n N_RESET_B_c_853_n 0.00488746f $X=5.69 $Y=0.87 $X2=0
+ $Y2=0
cc_458 N_A_211_363#_c_541_n N_RESET_B_c_853_n 2.59948e-19 $X=6.495 $Y=1.74 $X2=0
+ $Y2=0
cc_459 N_A_211_363#_c_523_n N_A_534_47#_M1011_g 0.0104452f $X=5.565 $Y=0.705
+ $X2=0 $Y2=0
cc_460 N_A_211_363#_c_525_n N_A_534_47#_c_995_n 8.91412e-19 $X=5.69 $Y=0.87
+ $X2=0 $Y2=0
cc_461 N_A_211_363#_c_526_n N_A_534_47#_c_995_n 0.00332535f $X=5.69 $Y=0.87
+ $X2=0 $Y2=0
cc_462 N_A_211_363#_c_535_n N_A_534_47#_c_995_n 0.00102943f $X=5.775 $Y=1.58
+ $X2=0 $Y2=0
cc_463 N_A_211_363#_c_538_n N_A_534_47#_c_995_n 9.64167e-19 $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_464 N_A_211_363#_c_535_n N_A_534_47#_c_996_n 9.82465e-19 $X=5.775 $Y=1.58
+ $X2=0 $Y2=0
cc_465 N_A_211_363#_c_538_n N_A_534_47#_c_996_n 0.00310577f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_466 N_A_211_363#_c_530_n N_A_534_47#_c_1006_n 0.00489977f $X=2.61 $Y=1.99
+ $X2=0 $Y2=0
cc_467 N_A_211_363#_c_538_n N_A_534_47#_c_1006_n 0.00524205f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_468 N_A_211_363#_c_539_n N_A_534_47#_c_1006_n 0.00310705f $X=2.955 $Y=1.87
+ $X2=0 $Y2=0
cc_469 N_A_211_363#_c_543_n N_A_534_47#_c_1006_n 0.0210219f $X=2.94 $Y=1.77
+ $X2=0 $Y2=0
cc_470 N_A_211_363#_M1019_g N_A_534_47#_c_1007_n 0.0120245f $X=3.135 $Y=0.415
+ $X2=0 $Y2=0
cc_471 N_A_211_363#_c_527_n N_A_534_47#_c_1007_n 0.0135671f $X=3.045 $Y=0.9
+ $X2=0 $Y2=0
cc_472 N_A_211_363#_c_528_n N_A_534_47#_c_1007_n 0.00340759f $X=3.135 $Y=0.9
+ $X2=0 $Y2=0
cc_473 N_A_211_363#_c_530_n N_A_534_47#_c_997_n 0.00108731f $X=2.61 $Y=1.99
+ $X2=0 $Y2=0
cc_474 N_A_211_363#_c_524_n N_A_534_47#_c_997_n 0.0155497f $X=2.94 $Y=1.575
+ $X2=0 $Y2=0
cc_475 N_A_211_363#_c_538_n N_A_534_47#_c_997_n 0.0156914f $X=6.41 $Y=1.87 $X2=0
+ $Y2=0
cc_476 N_A_211_363#_c_539_n N_A_534_47#_c_997_n 0.00128013f $X=2.955 $Y=1.87
+ $X2=0 $Y2=0
cc_477 N_A_211_363#_c_543_n N_A_534_47#_c_997_n 0.0288769f $X=2.94 $Y=1.77 $X2=0
+ $Y2=0
cc_478 N_A_211_363#_M1019_g N_A_534_47#_c_990_n 0.00658961f $X=3.135 $Y=0.415
+ $X2=0 $Y2=0
cc_479 N_A_211_363#_c_524_n N_A_534_47#_c_990_n 0.00727785f $X=2.94 $Y=1.575
+ $X2=0 $Y2=0
cc_480 N_A_211_363#_c_527_n N_A_534_47#_c_990_n 0.0136322f $X=3.045 $Y=0.9 $X2=0
+ $Y2=0
cc_481 N_A_211_363#_c_528_n N_A_534_47#_c_990_n 0.00151989f $X=3.135 $Y=0.9
+ $X2=0 $Y2=0
cc_482 N_A_211_363#_c_524_n N_A_534_47#_c_992_n 0.0122861f $X=2.94 $Y=1.575
+ $X2=0 $Y2=0
cc_483 N_A_211_363#_c_527_n N_A_534_47#_c_992_n 7.9625e-19 $X=3.045 $Y=0.9 $X2=0
+ $Y2=0
cc_484 N_A_211_363#_c_538_n N_A_534_47#_c_992_n 0.00764582f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_485 N_A_211_363#_c_526_n N_A_534_47#_c_994_n 0.0104452f $X=5.69 $Y=0.87 $X2=0
+ $Y2=0
cc_486 N_A_211_363#_c_531_n N_A_1323_21#_c_1118_n 0.0248077f $X=6.56 $Y=1.99
+ $X2=0 $Y2=0
cc_487 N_A_211_363#_c_541_n N_A_1323_21#_c_1118_n 0.0011829f $X=6.495 $Y=1.74
+ $X2=0 $Y2=0
cc_488 N_A_211_363#_c_531_n N_A_1323_21#_c_1132_n 0.0361201f $X=6.56 $Y=1.99
+ $X2=0 $Y2=0
cc_489 N_A_211_363#_c_531_n N_A_1323_21#_c_1129_n 5.49659e-19 $X=6.56 $Y=1.99
+ $X2=0 $Y2=0
cc_490 N_A_211_363#_c_523_n N_A_1128_47#_c_1275_n 0.00359811f $X=5.565 $Y=0.705
+ $X2=0 $Y2=0
cc_491 N_A_211_363#_c_525_n N_A_1128_47#_c_1275_n 0.00280345f $X=5.69 $Y=0.87
+ $X2=0 $Y2=0
cc_492 N_A_211_363#_c_526_n N_A_1128_47#_c_1275_n 0.00230884f $X=5.69 $Y=0.87
+ $X2=0 $Y2=0
cc_493 N_A_211_363#_c_531_n N_A_1128_47#_c_1278_n 0.0185724f $X=6.56 $Y=1.99
+ $X2=0 $Y2=0
cc_494 N_A_211_363#_c_534_n N_A_1128_47#_c_1278_n 0.0011512f $X=6.145 $Y=1.58
+ $X2=0 $Y2=0
cc_495 N_A_211_363#_c_538_n N_A_1128_47#_c_1278_n 0.00257887f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_496 N_A_211_363#_c_540_n N_A_1128_47#_c_1278_n 0.0034064f $X=6.555 $Y=1.87
+ $X2=0 $Y2=0
cc_497 N_A_211_363#_c_541_n N_A_1128_47#_c_1278_n 0.032649f $X=6.495 $Y=1.74
+ $X2=0 $Y2=0
cc_498 N_A_211_363#_c_540_n N_A_1128_47#_c_1270_n 0.00122541f $X=6.555 $Y=1.87
+ $X2=0 $Y2=0
cc_499 N_A_211_363#_c_541_n N_A_1128_47#_c_1270_n 3.14787e-19 $X=6.495 $Y=1.74
+ $X2=0 $Y2=0
cc_500 N_A_211_363#_c_531_n N_A_1128_47#_c_1271_n 0.00429683f $X=6.56 $Y=1.99
+ $X2=0 $Y2=0
cc_501 N_A_211_363#_c_540_n N_A_1128_47#_c_1271_n 0.0011225f $X=6.555 $Y=1.87
+ $X2=0 $Y2=0
cc_502 N_A_211_363#_c_541_n N_A_1128_47#_c_1271_n 0.0130673f $X=6.495 $Y=1.74
+ $X2=0 $Y2=0
cc_503 N_A_211_363#_c_531_n N_A_1128_47#_c_1272_n 0.0023218f $X=6.56 $Y=1.99
+ $X2=0 $Y2=0
cc_504 N_A_211_363#_c_540_n N_A_1128_47#_c_1272_n 0.00815331f $X=6.555 $Y=1.87
+ $X2=0 $Y2=0
cc_505 N_A_211_363#_c_531_n N_A_1128_47#_c_1274_n 0.00135273f $X=6.56 $Y=1.99
+ $X2=0 $Y2=0
cc_506 N_A_211_363#_c_541_n N_A_1128_47#_c_1274_n 0.0263238f $X=6.495 $Y=1.74
+ $X2=0 $Y2=0
cc_507 N_A_211_363#_c_538_n N_VPWR_M1017_s 0.00197335f $X=6.41 $Y=1.87 $X2=0
+ $Y2=0
cc_508 N_A_211_363#_c_529_n N_VPWR_c_1371_n 0.0202126f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_509 N_A_211_363#_c_536_n N_VPWR_c_1372_n 0.00331175f $X=2.665 $Y=1.87 $X2=0
+ $Y2=0
cc_510 N_A_211_363#_c_529_n N_VPWR_c_1372_n 0.00971431f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_511 N_A_211_363#_c_538_n N_VPWR_c_1373_n 0.0013967f $X=6.41 $Y=1.87 $X2=0
+ $Y2=0
cc_512 N_A_211_363#_c_538_n N_VPWR_c_1374_n 0.00349784f $X=6.41 $Y=1.87 $X2=0
+ $Y2=0
cc_513 N_A_211_363#_c_529_n N_VPWR_c_1380_n 0.0120448f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_514 N_A_211_363#_c_530_n N_VPWR_c_1382_n 0.00536466f $X=2.61 $Y=1.99 $X2=0
+ $Y2=0
cc_515 N_A_211_363#_c_543_n N_VPWR_c_1382_n 0.00228808f $X=2.94 $Y=1.77 $X2=0
+ $Y2=0
cc_516 N_A_211_363#_c_531_n N_VPWR_c_1384_n 0.00429453f $X=6.56 $Y=1.99 $X2=0
+ $Y2=0
cc_517 N_A_211_363#_c_530_n N_VPWR_c_1370_n 0.00747183f $X=2.61 $Y=1.99 $X2=0
+ $Y2=0
cc_518 N_A_211_363#_c_531_n N_VPWR_c_1370_n 0.00604257f $X=6.56 $Y=1.99 $X2=0
+ $Y2=0
cc_519 N_A_211_363#_c_536_n N_VPWR_c_1370_n 0.0632497f $X=2.665 $Y=1.87 $X2=0
+ $Y2=0
cc_520 N_A_211_363#_c_537_n N_VPWR_c_1370_n 0.0182006f $X=1.345 $Y=1.87 $X2=0
+ $Y2=0
cc_521 N_A_211_363#_c_538_n N_VPWR_c_1370_n 0.160365f $X=6.41 $Y=1.87 $X2=0
+ $Y2=0
cc_522 N_A_211_363#_c_539_n N_VPWR_c_1370_n 0.0159027f $X=2.955 $Y=1.87 $X2=0
+ $Y2=0
cc_523 N_A_211_363#_c_540_n N_VPWR_c_1370_n 0.0155966f $X=6.555 $Y=1.87 $X2=0
+ $Y2=0
cc_524 N_A_211_363#_c_529_n N_VPWR_c_1370_n 0.0029375f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_525 N_A_211_363#_c_543_n N_VPWR_c_1370_n 0.00171007f $X=2.94 $Y=1.77 $X2=0
+ $Y2=0
cc_526 N_A_211_363#_c_530_n N_A_436_413#_c_1526_n 0.00555682f $X=2.61 $Y=1.99
+ $X2=0 $Y2=0
cc_527 N_A_211_363#_c_524_n N_A_436_413#_c_1526_n 0.00584184f $X=2.94 $Y=1.575
+ $X2=0 $Y2=0
cc_528 N_A_211_363#_c_536_n N_A_436_413#_c_1526_n 0.0231912f $X=2.665 $Y=1.87
+ $X2=0 $Y2=0
cc_529 N_A_211_363#_c_539_n N_A_436_413#_c_1526_n 0.00120648f $X=2.955 $Y=1.87
+ $X2=0 $Y2=0
cc_530 N_A_211_363#_c_543_n N_A_436_413#_c_1526_n 0.0229875f $X=2.94 $Y=1.77
+ $X2=0 $Y2=0
cc_531 N_A_211_363#_c_538_n N_A_649_413#_c_1559_n 0.0328406f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_532 N_A_211_363#_c_538_n N_A_649_413#_c_1560_n 0.00857493f $X=6.41 $Y=1.87
+ $X2=0 $Y2=0
cc_533 N_A_211_363#_c_529_n N_VGND_c_1629_n 0.00732874f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_534 N_A_211_363#_c_529_n N_VGND_c_1630_n 0.00532595f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_535 N_A_211_363#_c_523_n N_VGND_c_1636_n 0.0055129f $X=5.565 $Y=0.705 $X2=0
+ $Y2=0
cc_536 N_A_211_363#_c_525_n N_VGND_c_1636_n 0.00198565f $X=5.69 $Y=0.87 $X2=0
+ $Y2=0
cc_537 N_A_211_363#_c_526_n N_VGND_c_1636_n 3.67755e-19 $X=5.69 $Y=0.87 $X2=0
+ $Y2=0
cc_538 N_A_211_363#_M1019_g N_VGND_c_1641_n 0.00368123f $X=3.135 $Y=0.415 $X2=0
+ $Y2=0
cc_539 N_A_211_363#_M1003_d N_VGND_c_1646_n 0.00535012f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_540 N_A_211_363#_M1019_g N_VGND_c_1646_n 0.00634244f $X=3.135 $Y=0.415 $X2=0
+ $Y2=0
cc_541 N_A_211_363#_c_523_n N_VGND_c_1646_n 0.00673892f $X=5.565 $Y=0.705 $X2=0
+ $Y2=0
cc_542 N_A_211_363#_c_525_n N_VGND_c_1646_n 0.00157806f $X=5.69 $Y=0.87 $X2=0
+ $Y2=0
cc_543 N_A_211_363#_c_529_n N_VGND_c_1646_n 0.00616598f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_544 N_A_751_289#_c_739_n N_RESET_B_c_848_n 0.0307401f $X=3.855 $Y=1.99 $X2=0
+ $Y2=0
cc_545 N_A_751_289#_M1005_g N_RESET_B_c_848_n 0.017872f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_546 N_A_751_289#_c_741_n N_RESET_B_c_848_n 0.0136984f $X=5.155 $Y=1.61 $X2=0
+ $Y2=0
cc_547 N_A_751_289#_c_738_n N_RESET_B_c_848_n 4.27876e-19 $X=5.24 $Y=1.525 $X2=0
+ $Y2=0
cc_548 N_A_751_289#_c_764_n N_RESET_B_c_848_n 0.00261768f $X=5.24 $Y=1.835 $X2=0
+ $Y2=0
cc_549 N_A_751_289#_c_770_n N_RESET_B_c_848_n 8.57239e-19 $X=5.325 $Y=1.92 $X2=0
+ $Y2=0
cc_550 N_A_751_289#_c_739_n N_RESET_B_c_860_n 0.0135184f $X=3.855 $Y=1.99 $X2=0
+ $Y2=0
cc_551 N_A_751_289#_M1005_g N_RESET_B_c_851_n 9.66214e-19 $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_552 N_A_751_289#_M1005_g N_RESET_B_c_852_n 0.0140645f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_553 N_A_751_289#_c_738_n N_RESET_B_c_852_n 0.00416146f $X=5.24 $Y=1.525 $X2=0
+ $Y2=0
cc_554 N_A_751_289#_c_755_n N_RESET_B_c_852_n 0.00174392f $X=5.195 $Y=0.835
+ $X2=0 $Y2=0
cc_555 N_A_751_289#_M1011_d N_RESET_B_c_853_n 7.46919e-19 $X=5.145 $Y=0.235
+ $X2=0 $Y2=0
cc_556 N_A_751_289#_c_741_n N_RESET_B_c_853_n 2.29961e-19 $X=5.155 $Y=1.61 $X2=0
+ $Y2=0
cc_557 N_A_751_289#_c_738_n N_RESET_B_c_853_n 0.00732299f $X=5.24 $Y=1.525 $X2=0
+ $Y2=0
cc_558 N_A_751_289#_c_788_p N_RESET_B_c_853_n 0.00383699f $X=5.3 $Y=0.36 $X2=0
+ $Y2=0
cc_559 N_A_751_289#_c_755_n N_RESET_B_c_853_n 0.010258f $X=5.195 $Y=0.835 $X2=0
+ $Y2=0
cc_560 N_A_751_289#_c_738_n N_RESET_B_c_854_n 0.00131045f $X=5.24 $Y=1.525 $X2=0
+ $Y2=0
cc_561 N_A_751_289#_c_755_n N_RESET_B_c_854_n 0.001782f $X=5.195 $Y=0.835 $X2=0
+ $Y2=0
cc_562 N_A_751_289#_M1005_g N_RESET_B_c_856_n 0.0637423f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_563 N_A_751_289#_c_762_n N_RESET_B_c_856_n 9.56876e-19 $X=5.195 $Y=0.705
+ $X2=0 $Y2=0
cc_564 N_A_751_289#_c_762_n N_A_534_47#_M1011_g 0.00765085f $X=5.195 $Y=0.705
+ $X2=0 $Y2=0
cc_565 N_A_751_289#_c_738_n N_A_534_47#_M1011_g 0.0131624f $X=5.24 $Y=1.525
+ $X2=0 $Y2=0
cc_566 N_A_751_289#_c_788_p N_A_534_47#_M1011_g 0.00354914f $X=5.3 $Y=0.36 $X2=0
+ $Y2=0
cc_567 N_A_751_289#_c_755_n N_A_534_47#_M1011_g 0.00550334f $X=5.195 $Y=0.835
+ $X2=0 $Y2=0
cc_568 N_A_751_289#_c_741_n N_A_534_47#_c_995_n 2.85533e-19 $X=5.155 $Y=1.61
+ $X2=0 $Y2=0
cc_569 N_A_751_289#_c_738_n N_A_534_47#_c_995_n 0.00905557f $X=5.24 $Y=1.525
+ $X2=0 $Y2=0
cc_570 N_A_751_289#_c_751_n N_A_534_47#_c_995_n 0.00146276f $X=5.645 $Y=1.92
+ $X2=0 $Y2=0
cc_571 N_A_751_289#_c_743_n N_A_534_47#_c_995_n 0.00504486f $X=5.24 $Y=1.61
+ $X2=0 $Y2=0
cc_572 N_A_751_289#_c_764_n N_A_534_47#_c_996_n 0.00526605f $X=5.24 $Y=1.835
+ $X2=0 $Y2=0
cc_573 N_A_751_289#_c_751_n N_A_534_47#_c_996_n 0.0159952f $X=5.645 $Y=1.92
+ $X2=0 $Y2=0
cc_574 N_A_751_289#_c_754_n N_A_534_47#_c_996_n 0.00472286f $X=5.73 $Y=2.3 $X2=0
+ $Y2=0
cc_575 N_A_751_289#_c_743_n N_A_534_47#_c_996_n 0.00385062f $X=5.24 $Y=1.61
+ $X2=0 $Y2=0
cc_576 N_A_751_289#_c_739_n N_A_534_47#_c_1006_n 0.00126119f $X=3.855 $Y=1.99
+ $X2=0 $Y2=0
cc_577 N_A_751_289#_M1005_g N_A_534_47#_c_1007_n 0.0046466f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_578 N_A_751_289#_c_739_n N_A_534_47#_c_997_n 0.00525152f $X=3.855 $Y=1.99
+ $X2=0 $Y2=0
cc_579 N_A_751_289#_M1005_g N_A_534_47#_c_997_n 0.00141578f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_580 N_A_751_289#_c_741_n N_A_534_47#_c_997_n 0.00842394f $X=5.155 $Y=1.61
+ $X2=0 $Y2=0
cc_581 N_A_751_289#_M1005_g N_A_534_47#_c_990_n 0.0114995f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_582 N_A_751_289#_c_739_n N_A_534_47#_c_991_n 0.00481281f $X=3.855 $Y=1.99
+ $X2=0 $Y2=0
cc_583 N_A_751_289#_M1005_g N_A_534_47#_c_991_n 0.0109415f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_584 N_A_751_289#_c_741_n N_A_534_47#_c_991_n 0.0694522f $X=5.155 $Y=1.61
+ $X2=0 $Y2=0
cc_585 N_A_751_289#_c_741_n N_A_534_47#_c_993_n 0.0116159f $X=5.155 $Y=1.61
+ $X2=0 $Y2=0
cc_586 N_A_751_289#_c_738_n N_A_534_47#_c_993_n 0.0244982f $X=5.24 $Y=1.525
+ $X2=0 $Y2=0
cc_587 N_A_751_289#_c_741_n N_A_534_47#_c_994_n 0.00941249f $X=5.155 $Y=1.61
+ $X2=0 $Y2=0
cc_588 N_A_751_289#_c_762_n N_A_1128_47#_c_1275_n 0.00388107f $X=5.195 $Y=0.705
+ $X2=0 $Y2=0
cc_589 N_A_751_289#_c_754_n N_A_1128_47#_c_1278_n 0.0206717f $X=5.73 $Y=2.3
+ $X2=0 $Y2=0
cc_590 N_A_751_289#_c_741_n N_VPWR_M1017_s 0.00130684f $X=5.155 $Y=1.61 $X2=0
+ $Y2=0
cc_591 N_A_751_289#_c_764_n N_VPWR_M1017_s 0.00436576f $X=5.24 $Y=1.835 $X2=0
+ $Y2=0
cc_592 N_A_751_289#_c_770_n N_VPWR_M1017_s 0.00463183f $X=5.325 $Y=1.92 $X2=0
+ $Y2=0
cc_593 N_A_751_289#_c_743_n N_VPWR_M1017_s 5.86854e-19 $X=5.24 $Y=1.61 $X2=0
+ $Y2=0
cc_594 N_A_751_289#_c_739_n N_VPWR_c_1373_n 0.00458065f $X=3.855 $Y=1.99 $X2=0
+ $Y2=0
cc_595 N_A_751_289#_c_741_n N_VPWR_c_1374_n 0.00261535f $X=5.155 $Y=1.61 $X2=0
+ $Y2=0
cc_596 N_A_751_289#_c_751_n N_VPWR_c_1374_n 0.00266364f $X=5.645 $Y=1.92 $X2=0
+ $Y2=0
cc_597 N_A_751_289#_c_770_n N_VPWR_c_1374_n 0.0134465f $X=5.325 $Y=1.92 $X2=0
+ $Y2=0
cc_598 N_A_751_289#_c_754_n N_VPWR_c_1374_n 0.0178901f $X=5.73 $Y=2.3 $X2=0
+ $Y2=0
cc_599 N_A_751_289#_c_739_n N_VPWR_c_1382_n 0.00525574f $X=3.855 $Y=1.99 $X2=0
+ $Y2=0
cc_600 N_A_751_289#_c_751_n N_VPWR_c_1384_n 0.00269374f $X=5.645 $Y=1.92 $X2=0
+ $Y2=0
cc_601 N_A_751_289#_c_754_n N_VPWR_c_1384_n 0.0117479f $X=5.73 $Y=2.3 $X2=0
+ $Y2=0
cc_602 N_A_751_289#_M1017_d N_VPWR_c_1370_n 0.00349593f $X=5.565 $Y=1.645 $X2=0
+ $Y2=0
cc_603 N_A_751_289#_c_739_n N_VPWR_c_1370_n 0.00713038f $X=3.855 $Y=1.99 $X2=0
+ $Y2=0
cc_604 N_A_751_289#_c_751_n N_VPWR_c_1370_n 0.00240965f $X=5.645 $Y=1.92 $X2=0
+ $Y2=0
cc_605 N_A_751_289#_c_770_n N_VPWR_c_1370_n 4.80263e-19 $X=5.325 $Y=1.92 $X2=0
+ $Y2=0
cc_606 N_A_751_289#_c_754_n N_VPWR_c_1370_n 0.00306902f $X=5.73 $Y=2.3 $X2=0
+ $Y2=0
cc_607 N_A_751_289#_c_739_n N_A_649_413#_c_1558_n 0.00426538f $X=3.855 $Y=1.99
+ $X2=0 $Y2=0
cc_608 N_A_751_289#_c_739_n N_A_649_413#_c_1559_n 0.0170667f $X=3.855 $Y=1.99
+ $X2=0 $Y2=0
cc_609 N_A_751_289#_c_741_n N_A_649_413#_c_1559_n 0.0615757f $X=5.155 $Y=1.61
+ $X2=0 $Y2=0
cc_610 N_A_751_289#_c_770_n N_A_649_413#_c_1559_n 0.00490929f $X=5.325 $Y=1.92
+ $X2=0 $Y2=0
cc_611 N_A_751_289#_c_762_n N_VGND_c_1631_n 0.00648459f $X=5.195 $Y=0.705 $X2=0
+ $Y2=0
cc_612 N_A_751_289#_c_788_p N_VGND_c_1631_n 0.0112895f $X=5.3 $Y=0.36 $X2=0
+ $Y2=0
cc_613 N_A_751_289#_c_788_p N_VGND_c_1636_n 0.0201433f $X=5.3 $Y=0.36 $X2=0
+ $Y2=0
cc_614 N_A_751_289#_M1005_g N_VGND_c_1641_n 0.00585385f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_615 N_A_751_289#_M1011_d N_VGND_c_1646_n 0.00245937f $X=5.145 $Y=0.235 $X2=0
+ $Y2=0
cc_616 N_A_751_289#_M1005_g N_VGND_c_1646_n 0.0067129f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_617 N_A_751_289#_c_788_p N_VGND_c_1646_n 0.00653072f $X=5.3 $Y=0.36 $X2=0
+ $Y2=0
cc_618 N_RESET_B_c_852_n N_A_534_47#_M1011_g 0.0015858f $X=4.55 $Y=0.85 $X2=0
+ $Y2=0
cc_619 N_RESET_B_c_853_n N_A_534_47#_M1011_g 0.00427213f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_620 N_RESET_B_c_854_n N_A_534_47#_M1011_g 0.00177034f $X=4.745 $Y=0.85 $X2=0
+ $Y2=0
cc_621 N_RESET_B_c_855_n N_A_534_47#_M1011_g 0.00598938f $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_856_n N_A_534_47#_M1011_g 0.0101327f $X=4.395 $Y=0.765 $X2=0
+ $Y2=0
cc_623 N_RESET_B_c_851_n N_A_534_47#_c_990_n 0.00211912f $X=4.63 $Y=0.85 $X2=0
+ $Y2=0
cc_624 N_RESET_B_c_852_n N_A_534_47#_c_990_n 0.0174468f $X=4.55 $Y=0.85 $X2=0
+ $Y2=0
cc_625 N_RESET_B_c_848_n N_A_534_47#_c_991_n 0.0112487f $X=4.39 $Y=1.89 $X2=0
+ $Y2=0
cc_626 N_RESET_B_c_851_n N_A_534_47#_c_991_n 8.00435e-19 $X=4.63 $Y=0.85 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_852_n N_A_534_47#_c_991_n 0.0538781f $X=4.55 $Y=0.85 $X2=0
+ $Y2=0
cc_628 N_RESET_B_c_853_n N_A_534_47#_c_991_n 4.07958e-19 $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_629 N_RESET_B_c_854_n N_A_534_47#_c_991_n 4.16664e-19 $X=4.745 $Y=0.85 $X2=0
+ $Y2=0
cc_630 N_RESET_B_c_855_n N_A_534_47#_c_991_n 0.00314016f $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_631 N_RESET_B_c_848_n N_A_534_47#_c_993_n 8.14528e-19 $X=4.39 $Y=1.89 $X2=0
+ $Y2=0
cc_632 N_RESET_B_c_852_n N_A_534_47#_c_993_n 8.03226e-19 $X=4.55 $Y=0.85 $X2=0
+ $Y2=0
cc_633 N_RESET_B_c_853_n N_A_534_47#_c_993_n 0.00422691f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_855_n N_A_534_47#_c_993_n 5.19504e-19 $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_635 N_RESET_B_c_848_n N_A_534_47#_c_994_n 0.0184537f $X=4.39 $Y=1.89 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_853_n N_A_534_47#_c_994_n 0.00102675f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_637 N_RESET_B_c_855_n N_A_534_47#_c_994_n 0.00613378f $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_638 N_RESET_B_c_853_n N_A_1323_21#_M1009_g 0.00239769f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_639 N_RESET_B_c_857_n N_A_1323_21#_c_1118_n 0.00970863f $X=7.695 $Y=1.12
+ $X2=0 $Y2=0
cc_640 N_RESET_B_c_858_n N_A_1323_21#_c_1118_n 0.00399835f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_850_n N_A_1323_21#_c_1132_n 0.00970863f $X=7.66 $Y=1.89 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_862_n N_A_1323_21#_c_1132_n 0.00960841f $X=7.66 $Y=1.99 $X2=0
+ $Y2=0
cc_643 N_RESET_B_M1021_g N_A_1323_21#_c_1121_n 3.6807e-19 $X=7.635 $Y=0.445
+ $X2=0 $Y2=0
cc_644 N_RESET_B_c_853_n N_A_1323_21#_c_1121_n 0.0124388f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_645 RESET_B N_A_1323_21#_c_1121_n 2.6274e-19 $X=7.635 $Y=0.765 $X2=0 $Y2=0
cc_646 N_RESET_B_c_858_n N_A_1323_21#_c_1121_n 0.014229f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_647 N_RESET_B_M1021_g N_A_1323_21#_c_1156_n 0.012015f $X=7.635 $Y=0.445 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_853_n N_A_1323_21#_c_1156_n 0.00464811f $X=7.575 $Y=0.85
+ $X2=0 $Y2=0
cc_649 RESET_B N_A_1323_21#_c_1156_n 9.43613e-19 $X=7.635 $Y=0.765 $X2=0 $Y2=0
cc_650 N_RESET_B_c_857_n N_A_1323_21#_c_1156_n 3.87365e-19 $X=7.695 $Y=1.12
+ $X2=0 $Y2=0
cc_651 N_RESET_B_c_858_n N_A_1323_21#_c_1156_n 0.0200404f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_652 N_RESET_B_c_862_n N_A_1323_21#_c_1136_n 0.00534288f $X=7.66 $Y=1.99 $X2=0
+ $Y2=0
cc_653 RESET_B N_A_1323_21#_c_1123_n 0.00157555f $X=7.635 $Y=0.765 $X2=0 $Y2=0
cc_654 N_RESET_B_c_858_n N_A_1323_21#_c_1123_n 0.0186693f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_655 N_RESET_B_c_858_n N_A_1323_21#_c_1124_n 0.00395187f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_656 N_RESET_B_M1021_g N_A_1323_21#_c_1126_n 0.00672753f $X=7.635 $Y=0.445
+ $X2=0 $Y2=0
cc_657 N_RESET_B_c_858_n N_A_1323_21#_c_1126_n 0.0169692f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_658 N_RESET_B_c_853_n N_A_1323_21#_c_1127_n 0.0165023f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_659 RESET_B N_A_1323_21#_c_1127_n 3.01996e-19 $X=7.635 $Y=0.765 $X2=0 $Y2=0
cc_660 N_RESET_B_c_858_n N_A_1323_21#_c_1128_n 0.0111143f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_661 N_RESET_B_M1021_g N_A_1323_21#_c_1129_n 0.0118207f $X=7.635 $Y=0.445
+ $X2=0 $Y2=0
cc_662 N_RESET_B_c_853_n N_A_1323_21#_c_1129_n 0.00568196f $X=7.575 $Y=0.85
+ $X2=0 $Y2=0
cc_663 N_RESET_B_c_858_n N_A_1323_21#_c_1129_n 0.00204709f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_664 N_RESET_B_c_850_n N_A_1128_47#_c_1268_n 0.0295113f $X=7.66 $Y=1.89 $X2=0
+ $Y2=0
cc_665 N_RESET_B_c_862_n N_A_1128_47#_c_1268_n 0.0119493f $X=7.66 $Y=1.99 $X2=0
+ $Y2=0
cc_666 N_RESET_B_M1021_g N_A_1128_47#_M1022_g 0.0262711f $X=7.635 $Y=0.445 $X2=0
+ $Y2=0
cc_667 N_RESET_B_c_850_n N_A_1128_47#_M1022_g 0.00757221f $X=7.66 $Y=1.89 $X2=0
+ $Y2=0
cc_668 N_RESET_B_c_857_n N_A_1128_47#_M1022_g 0.015633f $X=7.695 $Y=1.12 $X2=0
+ $Y2=0
cc_669 N_RESET_B_c_858_n N_A_1128_47#_M1022_g 0.0071022f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_670 N_RESET_B_c_853_n N_A_1128_47#_c_1275_n 0.0119217f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_671 N_RESET_B_c_853_n N_A_1128_47#_c_1267_n 0.0198537f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_672 N_RESET_B_c_853_n N_A_1128_47#_c_1270_n 0.00591815f $X=7.575 $Y=0.85
+ $X2=0 $Y2=0
cc_673 N_RESET_B_c_850_n N_A_1128_47#_c_1272_n 0.00123249f $X=7.66 $Y=1.89 $X2=0
+ $Y2=0
cc_674 N_RESET_B_c_862_n N_A_1128_47#_c_1272_n 6.69096e-19 $X=7.66 $Y=1.99 $X2=0
+ $Y2=0
cc_675 N_RESET_B_c_850_n N_A_1128_47#_c_1273_n 0.0184545f $X=7.66 $Y=1.89 $X2=0
+ $Y2=0
cc_676 RESET_B N_A_1128_47#_c_1273_n 8.81753e-19 $X=7.635 $Y=0.765 $X2=0 $Y2=0
cc_677 N_RESET_B_c_857_n N_A_1128_47#_c_1273_n 4.16268e-19 $X=7.695 $Y=1.12
+ $X2=0 $Y2=0
cc_678 N_RESET_B_c_858_n N_A_1128_47#_c_1273_n 0.0314839f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_679 N_RESET_B_c_850_n N_A_1128_47#_c_1274_n 0.00113482f $X=7.66 $Y=1.89 $X2=0
+ $Y2=0
cc_680 N_RESET_B_c_853_n N_A_1128_47#_c_1274_n 0.00477698f $X=7.575 $Y=0.85
+ $X2=0 $Y2=0
cc_681 N_RESET_B_c_858_n N_A_1128_47#_c_1274_n 0.00340885f $X=7.72 $Y=0.85 $X2=0
+ $Y2=0
cc_682 N_RESET_B_c_860_n N_VPWR_c_1373_n 0.0117385f $X=4.39 $Y=1.99 $X2=0 $Y2=0
cc_683 N_RESET_B_c_860_n N_VPWR_c_1374_n 0.00502266f $X=4.39 $Y=1.99 $X2=0 $Y2=0
cc_684 N_RESET_B_c_862_n N_VPWR_c_1375_n 0.00869911f $X=7.66 $Y=1.99 $X2=0 $Y2=0
cc_685 N_RESET_B_c_860_n N_VPWR_c_1388_n 0.0046377f $X=4.39 $Y=1.99 $X2=0 $Y2=0
cc_686 N_RESET_B_c_862_n N_VPWR_c_1389_n 0.00643335f $X=7.66 $Y=1.99 $X2=0 $Y2=0
cc_687 N_RESET_B_c_862_n N_VPWR_c_1393_n 7.70004e-19 $X=7.66 $Y=1.99 $X2=0 $Y2=0
cc_688 N_RESET_B_c_860_n N_VPWR_c_1370_n 0.0062934f $X=4.39 $Y=1.99 $X2=0 $Y2=0
cc_689 N_RESET_B_c_862_n N_VPWR_c_1370_n 0.0108009f $X=7.66 $Y=1.99 $X2=0 $Y2=0
cc_690 N_RESET_B_c_848_n N_A_649_413#_c_1559_n 0.00268737f $X=4.39 $Y=1.89 $X2=0
+ $Y2=0
cc_691 N_RESET_B_c_860_n N_A_649_413#_c_1559_n 0.0117053f $X=4.39 $Y=1.99 $X2=0
+ $Y2=0
cc_692 N_RESET_B_c_860_n N_A_649_413#_c_1561_n 0.00449002f $X=4.39 $Y=1.99 $X2=0
+ $Y2=0
cc_693 N_RESET_B_c_853_n N_VGND_M1007_d 0.00351032f $X=7.575 $Y=0.85 $X2=0 $Y2=0
cc_694 N_RESET_B_c_854_n N_VGND_M1007_d 8.33031e-19 $X=4.745 $Y=0.85 $X2=0 $Y2=0
cc_695 N_RESET_B_c_851_n N_VGND_c_1631_n 0.00336536f $X=4.63 $Y=0.85 $X2=0 $Y2=0
cc_696 N_RESET_B_c_852_n N_VGND_c_1631_n 0.00639968f $X=4.55 $Y=0.85 $X2=0 $Y2=0
cc_697 N_RESET_B_c_853_n N_VGND_c_1631_n 0.00182136f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_698 N_RESET_B_c_855_n N_VGND_c_1631_n 2.19293e-19 $X=4.37 $Y=0.93 $X2=0 $Y2=0
cc_699 N_RESET_B_c_856_n N_VGND_c_1631_n 0.0112955f $X=4.395 $Y=0.765 $X2=0
+ $Y2=0
cc_700 N_RESET_B_M1021_g N_VGND_c_1632_n 0.00368875f $X=7.635 $Y=0.445 $X2=0
+ $Y2=0
cc_701 N_RESET_B_c_853_n N_VGND_c_1632_n 0.00458378f $X=7.575 $Y=0.85 $X2=0
+ $Y2=0
cc_702 N_RESET_B_M1021_g N_VGND_c_1638_n 0.00366111f $X=7.635 $Y=0.445 $X2=0
+ $Y2=0
cc_703 N_RESET_B_c_855_n N_VGND_c_1641_n 0.00100696f $X=4.37 $Y=0.93 $X2=0 $Y2=0
cc_704 N_RESET_B_c_856_n N_VGND_c_1641_n 0.00585385f $X=4.395 $Y=0.765 $X2=0
+ $Y2=0
cc_705 N_RESET_B_M1021_g N_VGND_c_1646_n 0.00683955f $X=7.635 $Y=0.445 $X2=0
+ $Y2=0
cc_706 N_RESET_B_c_851_n N_VGND_c_1646_n 0.0408566f $X=4.63 $Y=0.85 $X2=0 $Y2=0
cc_707 N_RESET_B_c_852_n N_VGND_c_1646_n 0.0119964f $X=4.55 $Y=0.85 $X2=0 $Y2=0
cc_708 N_RESET_B_c_853_n N_VGND_c_1646_n 0.134751f $X=7.575 $Y=0.85 $X2=0 $Y2=0
cc_709 RESET_B N_VGND_c_1646_n 0.0144453f $X=7.635 $Y=0.765 $X2=0 $Y2=0
cc_710 N_RESET_B_c_856_n N_VGND_c_1646_n 0.00624005f $X=4.395 $Y=0.765 $X2=0
+ $Y2=0
cc_711 N_RESET_B_c_858_n A_1542_47# 0.00172041f $X=7.72 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_712 N_A_534_47#_c_996_n N_VPWR_c_1374_n 0.0112655f $X=5.475 $Y=1.57 $X2=0
+ $Y2=0
cc_713 N_A_534_47#_c_994_n N_VPWR_c_1374_n 0.00136666f $X=4.9 $Y=1.17 $X2=0
+ $Y2=0
cc_714 N_A_534_47#_c_1006_n N_VPWR_c_1382_n 0.0397322f $X=3.195 $Y=2.3 $X2=0
+ $Y2=0
cc_715 N_A_534_47#_c_996_n N_VPWR_c_1384_n 0.00406603f $X=5.475 $Y=1.57 $X2=0
+ $Y2=0
cc_716 N_A_534_47#_M1028_d N_VPWR_c_1370_n 0.00234562f $X=2.7 $Y=2.065 $X2=0
+ $Y2=0
cc_717 N_A_534_47#_c_996_n N_VPWR_c_1370_n 0.0046037f $X=5.475 $Y=1.57 $X2=0
+ $Y2=0
cc_718 N_A_534_47#_c_1006_n N_VPWR_c_1370_n 0.0114216f $X=3.195 $Y=2.3 $X2=0
+ $Y2=0
cc_719 N_A_534_47#_c_1006_n N_A_436_413#_c_1526_n 0.0188635f $X=3.195 $Y=2.3
+ $X2=0 $Y2=0
cc_720 N_A_534_47#_c_1006_n N_A_649_413#_M1004_d 0.00438274f $X=3.195 $Y=2.3
+ $X2=-0.19 $Y2=-0.24
cc_721 N_A_534_47#_c_997_n N_A_649_413#_M1004_d 6.31229e-19 $X=3.28 $Y=2.135
+ $X2=-0.19 $Y2=-0.24
cc_722 N_A_534_47#_c_1006_n N_A_649_413#_c_1558_n 0.0195259f $X=3.195 $Y=2.3
+ $X2=0 $Y2=0
cc_723 N_A_534_47#_c_997_n N_A_649_413#_c_1558_n 0.00726911f $X=3.28 $Y=2.135
+ $X2=0 $Y2=0
cc_724 N_A_534_47#_c_996_n N_A_649_413#_c_1559_n 0.00129931f $X=5.475 $Y=1.57
+ $X2=0 $Y2=0
cc_725 N_A_534_47#_c_991_n N_A_649_413#_c_1559_n 4.0432e-19 $X=4.815 $Y=1.27
+ $X2=0 $Y2=0
cc_726 N_A_534_47#_c_997_n N_A_649_413#_c_1560_n 0.0133546f $X=3.28 $Y=2.135
+ $X2=0 $Y2=0
cc_727 N_A_534_47#_c_992_n N_A_649_413#_c_1560_n 0.0035943f $X=3.6 $Y=1.27 $X2=0
+ $Y2=0
cc_728 N_A_534_47#_c_996_n N_A_649_413#_c_1561_n 0.00258461f $X=5.475 $Y=1.57
+ $X2=0 $Y2=0
cc_729 N_A_534_47#_M1011_g N_VGND_c_1631_n 0.00658363f $X=5.07 $Y=0.555 $X2=0
+ $Y2=0
cc_730 N_A_534_47#_c_991_n N_VGND_c_1631_n 0.00221854f $X=4.815 $Y=1.27 $X2=0
+ $Y2=0
cc_731 N_A_534_47#_c_993_n N_VGND_c_1631_n 6.77929e-19 $X=4.9 $Y=1.17 $X2=0
+ $Y2=0
cc_732 N_A_534_47#_c_994_n N_VGND_c_1631_n 0.001314f $X=4.9 $Y=1.17 $X2=0 $Y2=0
cc_733 N_A_534_47#_M1011_g N_VGND_c_1636_n 0.00466263f $X=5.07 $Y=0.555 $X2=0
+ $Y2=0
cc_734 N_A_534_47#_c_1007_n N_VGND_c_1641_n 0.0410995f $X=3.43 $Y=0.39 $X2=0
+ $Y2=0
cc_735 N_A_534_47#_M1015_d N_VGND_c_1646_n 0.00362422f $X=2.67 $Y=0.235 $X2=0
+ $Y2=0
cc_736 N_A_534_47#_M1011_g N_VGND_c_1646_n 0.00661852f $X=5.07 $Y=0.555 $X2=0
+ $Y2=0
cc_737 N_A_534_47#_c_1007_n N_VGND_c_1646_n 0.0322161f $X=3.43 $Y=0.39 $X2=0
+ $Y2=0
cc_738 N_A_534_47#_c_1007_n A_642_47# 0.0142113f $X=3.43 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_739 N_A_534_47#_c_990_n A_642_47# 0.00606937f $X=3.515 $Y=1.185 $X2=-0.19
+ $Y2=-0.24
cc_740 N_A_1323_21#_c_1135_n N_A_1128_47#_c_1268_n 0.0158639f $X=8.44 $Y=2 $X2=0
+ $Y2=0
cc_741 N_A_1323_21#_c_1136_n N_A_1128_47#_c_1268_n 2.53623e-19 $X=7.98 $Y=2
+ $X2=0 $Y2=0
cc_742 N_A_1323_21#_c_1124_n N_A_1128_47#_c_1268_n 0.00703285f $X=8.525 $Y=1.915
+ $X2=0 $Y2=0
cc_743 N_A_1323_21#_c_1156_n N_A_1128_47#_M1022_g 0.0129796f $X=8.29 $Y=0.38
+ $X2=0 $Y2=0
cc_744 N_A_1323_21#_c_1123_n N_A_1128_47#_M1022_g 0.0109251f $X=8.462 $Y=1.075
+ $X2=0 $Y2=0
cc_745 N_A_1323_21#_c_1124_n N_A_1128_47#_M1022_g 0.00825738f $X=8.525 $Y=1.915
+ $X2=0 $Y2=0
cc_746 N_A_1323_21#_c_1128_n N_A_1128_47#_M1022_g 0.00599567f $X=8.29 $Y=1.075
+ $X2=0 $Y2=0
cc_747 N_A_1323_21#_M1009_g N_A_1128_47#_c_1275_n 0.00822642f $X=6.69 $Y=0.445
+ $X2=0 $Y2=0
cc_748 N_A_1323_21#_c_1126_n N_A_1128_47#_c_1275_n 3.32251e-19 $X=7.145 $Y=0.695
+ $X2=0 $Y2=0
cc_749 N_A_1323_21#_c_1132_n N_A_1128_47#_c_1278_n 0.0123388f $X=6.97 $Y=1.99
+ $X2=0 $Y2=0
cc_750 N_A_1323_21#_M1009_g N_A_1128_47#_c_1267_n 0.00759465f $X=6.69 $Y=0.445
+ $X2=0 $Y2=0
cc_751 N_A_1323_21#_c_1126_n N_A_1128_47#_c_1267_n 0.0048113f $X=7.145 $Y=0.695
+ $X2=0 $Y2=0
cc_752 N_A_1323_21#_c_1127_n N_A_1128_47#_c_1267_n 0.0198469f $X=7.145 $Y=0.865
+ $X2=0 $Y2=0
cc_753 N_A_1323_21#_c_1129_n N_A_1128_47#_c_1267_n 0.0105225f $X=6.97 $Y=0.98
+ $X2=0 $Y2=0
cc_754 N_A_1323_21#_c_1118_n N_A_1128_47#_c_1270_n 0.00134264f $X=6.97 $Y=1.89
+ $X2=0 $Y2=0
cc_755 N_A_1323_21#_c_1129_n N_A_1128_47#_c_1270_n 0.00566981f $X=6.97 $Y=0.98
+ $X2=0 $Y2=0
cc_756 N_A_1323_21#_c_1118_n N_A_1128_47#_c_1272_n 0.00450946f $X=6.97 $Y=1.89
+ $X2=0 $Y2=0
cc_757 N_A_1323_21#_c_1132_n N_A_1128_47#_c_1272_n 0.00757038f $X=6.97 $Y=1.99
+ $X2=0 $Y2=0
cc_758 N_A_1323_21#_c_1118_n N_A_1128_47#_c_1273_n 0.00463648f $X=6.97 $Y=1.89
+ $X2=0 $Y2=0
cc_759 N_A_1323_21#_c_1121_n N_A_1128_47#_c_1273_n 0.00651701f $X=7.04 $Y=0.98
+ $X2=0 $Y2=0
cc_760 N_A_1323_21#_c_1135_n N_A_1128_47#_c_1273_n 0.0200685f $X=8.44 $Y=2 $X2=0
+ $Y2=0
cc_761 N_A_1323_21#_c_1136_n N_A_1128_47#_c_1273_n 0.0138731f $X=7.98 $Y=2 $X2=0
+ $Y2=0
cc_762 N_A_1323_21#_c_1124_n N_A_1128_47#_c_1273_n 0.0141871f $X=8.525 $Y=1.915
+ $X2=0 $Y2=0
cc_763 N_A_1323_21#_c_1129_n N_A_1128_47#_c_1273_n 8.79183e-19 $X=6.97 $Y=0.98
+ $X2=0 $Y2=0
cc_764 N_A_1323_21#_c_1118_n N_A_1128_47#_c_1274_n 0.0215514f $X=6.97 $Y=1.89
+ $X2=0 $Y2=0
cc_765 N_A_1323_21#_c_1121_n N_A_1128_47#_c_1274_n 0.00750417f $X=7.04 $Y=0.98
+ $X2=0 $Y2=0
cc_766 N_A_1323_21#_c_1129_n N_A_1128_47#_c_1274_n 0.00115411f $X=6.97 $Y=0.98
+ $X2=0 $Y2=0
cc_767 N_A_1323_21#_c_1135_n N_VPWR_M1013_d 0.00227961f $X=8.44 $Y=2 $X2=0 $Y2=0
cc_768 N_A_1323_21#_c_1132_n N_VPWR_c_1375_n 0.00479765f $X=6.97 $Y=1.99 $X2=0
+ $Y2=0
cc_769 N_A_1323_21#_c_1202_p N_VPWR_c_1375_n 0.011854f $X=7.895 $Y=2.21 $X2=0
+ $Y2=0
cc_770 N_A_1323_21#_c_1135_n N_VPWR_c_1376_n 0.00141081f $X=8.44 $Y=2 $X2=0
+ $Y2=0
cc_771 N_A_1323_21#_c_1133_n N_VPWR_c_1377_n 0.01287f $X=9.13 $Y=1.41 $X2=0
+ $Y2=0
cc_772 N_A_1323_21#_c_1135_n N_VPWR_c_1377_n 0.0125643f $X=8.44 $Y=2 $X2=0 $Y2=0
cc_773 N_A_1323_21#_c_1124_n N_VPWR_c_1377_n 0.0223334f $X=8.525 $Y=1.915 $X2=0
+ $Y2=0
cc_774 N_A_1323_21#_c_1125_n N_VPWR_c_1377_n 0.00960121f $X=9.17 $Y=1.16 $X2=0
+ $Y2=0
cc_775 N_A_1323_21#_c_1134_n N_VPWR_c_1379_n 0.00702795f $X=9.6 $Y=1.41 $X2=0
+ $Y2=0
cc_776 N_A_1323_21#_c_1132_n N_VPWR_c_1384_n 0.00535679f $X=6.97 $Y=1.99 $X2=0
+ $Y2=0
cc_777 N_A_1323_21#_c_1202_p N_VPWR_c_1389_n 0.00725596f $X=7.895 $Y=2.21 $X2=0
+ $Y2=0
cc_778 N_A_1323_21#_c_1135_n N_VPWR_c_1389_n 0.00257098f $X=8.44 $Y=2 $X2=0
+ $Y2=0
cc_779 N_A_1323_21#_c_1133_n N_VPWR_c_1390_n 0.00702461f $X=9.13 $Y=1.41 $X2=0
+ $Y2=0
cc_780 N_A_1323_21#_c_1134_n N_VPWR_c_1390_n 0.00673617f $X=9.6 $Y=1.41 $X2=0
+ $Y2=0
cc_781 N_A_1323_21#_c_1202_p N_VPWR_c_1393_n 0.00857113f $X=7.895 $Y=2.21 $X2=0
+ $Y2=0
cc_782 N_A_1323_21#_c_1135_n N_VPWR_c_1393_n 0.0249983f $X=8.44 $Y=2 $X2=0 $Y2=0
cc_783 N_A_1323_21#_M1025_d N_VPWR_c_1370_n 0.00459686f $X=7.75 $Y=2.065 $X2=0
+ $Y2=0
cc_784 N_A_1323_21#_c_1132_n N_VPWR_c_1370_n 0.00875627f $X=6.97 $Y=1.99 $X2=0
+ $Y2=0
cc_785 N_A_1323_21#_c_1133_n N_VPWR_c_1370_n 0.0137919f $X=9.13 $Y=1.41 $X2=0
+ $Y2=0
cc_786 N_A_1323_21#_c_1134_n N_VPWR_c_1370_n 0.0127777f $X=9.6 $Y=1.41 $X2=0
+ $Y2=0
cc_787 N_A_1323_21#_c_1202_p N_VPWR_c_1370_n 0.00608739f $X=7.895 $Y=2.21 $X2=0
+ $Y2=0
cc_788 N_A_1323_21#_c_1135_n N_VPWR_c_1370_n 0.00842505f $X=8.44 $Y=2 $X2=0
+ $Y2=0
cc_789 N_A_1323_21#_c_1119_n N_Q_c_1600_n 0.00560572f $X=9.105 $Y=0.995 $X2=0
+ $Y2=0
cc_790 N_A_1323_21#_c_1134_n N_Q_c_1601_n 0.0157372f $X=9.6 $Y=1.41 $X2=0 $Y2=0
cc_791 N_A_1323_21#_c_1119_n Q 0.00322766f $X=9.105 $Y=0.995 $X2=0 $Y2=0
cc_792 N_A_1323_21#_c_1133_n Q 2.21352e-19 $X=9.13 $Y=1.41 $X2=0 $Y2=0
cc_793 N_A_1323_21#_c_1134_n Q 0.00208431f $X=9.6 $Y=1.41 $X2=0 $Y2=0
cc_794 N_A_1323_21#_c_1120_n Q 0.0161544f $X=9.625 $Y=0.995 $X2=0 $Y2=0
cc_795 N_A_1323_21#_c_1123_n Q 3.27806e-19 $X=8.462 $Y=1.075 $X2=0 $Y2=0
cc_796 N_A_1323_21#_c_1125_n Q 0.0242623f $X=9.17 $Y=1.16 $X2=0 $Y2=0
cc_797 N_A_1323_21#_c_1130_n Q 0.0281063f $X=9.6 $Y=1.202 $X2=0 $Y2=0
cc_798 N_A_1323_21#_c_1133_n Q 4.93703e-19 $X=9.13 $Y=1.41 $X2=0 $Y2=0
cc_799 N_A_1323_21#_c_1134_n Q 0.0168732f $X=9.6 $Y=1.41 $X2=0 $Y2=0
cc_800 N_A_1323_21#_c_1124_n Q 0.00230759f $X=8.525 $Y=1.915 $X2=0 $Y2=0
cc_801 N_A_1323_21#_c_1125_n Q 0.0069008f $X=9.17 $Y=1.16 $X2=0 $Y2=0
cc_802 N_A_1323_21#_c_1130_n Q 0.00754122f $X=9.6 $Y=1.202 $X2=0 $Y2=0
cc_803 N_A_1323_21#_c_1156_n N_VGND_M1009_d 0.0046492f $X=8.29 $Y=0.38 $X2=0
+ $Y2=0
cc_804 N_A_1323_21#_c_1237_p N_VGND_M1009_d 0.00501365f $X=7.335 $Y=0.38 $X2=0
+ $Y2=0
cc_805 N_A_1323_21#_c_1126_n N_VGND_M1009_d 0.00623681f $X=7.145 $Y=0.695 $X2=0
+ $Y2=0
cc_806 N_A_1323_21#_M1009_g N_VGND_c_1632_n 0.00539093f $X=6.69 $Y=0.445 $X2=0
+ $Y2=0
cc_807 N_A_1323_21#_c_1237_p N_VGND_c_1632_n 0.0138309f $X=7.335 $Y=0.38 $X2=0
+ $Y2=0
cc_808 N_A_1323_21#_c_1126_n N_VGND_c_1632_n 0.00432168f $X=7.145 $Y=0.695 $X2=0
+ $Y2=0
cc_809 N_A_1323_21#_c_1127_n N_VGND_c_1632_n 0.00296625f $X=7.145 $Y=0.865 $X2=0
+ $Y2=0
cc_810 N_A_1323_21#_c_1129_n N_VGND_c_1632_n 0.00449912f $X=6.97 $Y=0.98 $X2=0
+ $Y2=0
cc_811 N_A_1323_21#_c_1119_n N_VGND_c_1633_n 0.00460404f $X=9.105 $Y=0.995 $X2=0
+ $Y2=0
cc_812 N_A_1323_21#_c_1122_n N_VGND_c_1633_n 0.0138368f $X=8.462 $Y=0.465 $X2=0
+ $Y2=0
cc_813 N_A_1323_21#_c_1123_n N_VGND_c_1633_n 0.0329132f $X=8.462 $Y=1.075 $X2=0
+ $Y2=0
cc_814 N_A_1323_21#_c_1125_n N_VGND_c_1633_n 0.0138247f $X=9.17 $Y=1.16 $X2=0
+ $Y2=0
cc_815 N_A_1323_21#_c_1120_n N_VGND_c_1635_n 0.00438629f $X=9.625 $Y=0.995 $X2=0
+ $Y2=0
cc_816 N_A_1323_21#_M1009_g N_VGND_c_1636_n 0.0052466f $X=6.69 $Y=0.445 $X2=0
+ $Y2=0
cc_817 N_A_1323_21#_c_1156_n N_VGND_c_1638_n 0.0428842f $X=8.29 $Y=0.38 $X2=0
+ $Y2=0
cc_818 N_A_1323_21#_c_1237_p N_VGND_c_1638_n 0.0094263f $X=7.335 $Y=0.38 $X2=0
+ $Y2=0
cc_819 N_A_1323_21#_c_1122_n N_VGND_c_1638_n 0.0192713f $X=8.462 $Y=0.465 $X2=0
+ $Y2=0
cc_820 N_A_1323_21#_c_1127_n N_VGND_c_1638_n 0.00295587f $X=7.145 $Y=0.865 $X2=0
+ $Y2=0
cc_821 N_A_1323_21#_c_1119_n N_VGND_c_1642_n 0.00540385f $X=9.105 $Y=0.995 $X2=0
+ $Y2=0
cc_822 N_A_1323_21#_c_1120_n N_VGND_c_1642_n 0.00439206f $X=9.625 $Y=0.995 $X2=0
+ $Y2=0
cc_823 N_A_1323_21#_M1022_d N_VGND_c_1646_n 0.00212393f $X=8.24 $Y=0.235 $X2=0
+ $Y2=0
cc_824 N_A_1323_21#_M1009_g N_VGND_c_1646_n 0.00767715f $X=6.69 $Y=0.445 $X2=0
+ $Y2=0
cc_825 N_A_1323_21#_c_1119_n N_VGND_c_1646_n 0.0110239f $X=9.105 $Y=0.995 $X2=0
+ $Y2=0
cc_826 N_A_1323_21#_c_1120_n N_VGND_c_1646_n 0.00713099f $X=9.625 $Y=0.995 $X2=0
+ $Y2=0
cc_827 N_A_1323_21#_c_1156_n N_VGND_c_1646_n 0.0229709f $X=8.29 $Y=0.38 $X2=0
+ $Y2=0
cc_828 N_A_1323_21#_c_1237_p N_VGND_c_1646_n 0.00303501f $X=7.335 $Y=0.38 $X2=0
+ $Y2=0
cc_829 N_A_1323_21#_c_1122_n N_VGND_c_1646_n 0.013024f $X=8.462 $Y=0.465 $X2=0
+ $Y2=0
cc_830 N_A_1323_21#_c_1127_n N_VGND_c_1646_n 0.00230277f $X=7.145 $Y=0.865 $X2=0
+ $Y2=0
cc_831 N_A_1323_21#_c_1129_n N_VGND_c_1646_n 3.40468e-19 $X=6.97 $Y=0.98 $X2=0
+ $Y2=0
cc_832 N_A_1323_21#_c_1156_n A_1542_47# 0.00913475f $X=8.29 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_833 N_A_1128_47#_c_1268_n N_VPWR_c_1375_n 7.10488e-19 $X=8.14 $Y=1.99 $X2=0
+ $Y2=0
cc_834 N_A_1128_47#_c_1278_n N_VPWR_c_1375_n 0.0138682f $X=6.835 $Y=2.295 $X2=0
+ $Y2=0
cc_835 N_A_1128_47#_c_1273_n N_VPWR_c_1375_n 0.00900963f $X=8.105 $Y=1.66 $X2=0
+ $Y2=0
cc_836 N_A_1128_47#_c_1268_n N_VPWR_c_1377_n 0.0041455f $X=8.14 $Y=1.99 $X2=0
+ $Y2=0
cc_837 N_A_1128_47#_c_1278_n N_VPWR_c_1384_n 0.0560426f $X=6.835 $Y=2.295 $X2=0
+ $Y2=0
cc_838 N_A_1128_47#_c_1268_n N_VPWR_c_1389_n 0.00315029f $X=8.14 $Y=1.99 $X2=0
+ $Y2=0
cc_839 N_A_1128_47#_c_1268_n N_VPWR_c_1393_n 0.011239f $X=8.14 $Y=1.99 $X2=0
+ $Y2=0
cc_840 N_A_1128_47#_M1018_d N_VPWR_c_1370_n 0.00235763f $X=6.11 $Y=2.065 $X2=0
+ $Y2=0
cc_841 N_A_1128_47#_c_1268_n N_VPWR_c_1370_n 0.00380683f $X=8.14 $Y=1.99 $X2=0
+ $Y2=0
cc_842 N_A_1128_47#_c_1278_n N_VPWR_c_1370_n 0.0217736f $X=6.835 $Y=2.295 $X2=0
+ $Y2=0
cc_843 N_A_1128_47#_c_1278_n A_1330_413# 0.00337251f $X=6.835 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_844 N_A_1128_47#_c_1275_n N_VGND_c_1632_n 0.0212215f $X=6.485 $Y=0.395 $X2=0
+ $Y2=0
cc_845 N_A_1128_47#_M1022_g N_VGND_c_1633_n 0.00271655f $X=8.165 $Y=0.445 $X2=0
+ $Y2=0
cc_846 N_A_1128_47#_c_1275_n N_VGND_c_1636_n 0.055255f $X=6.485 $Y=0.395 $X2=0
+ $Y2=0
cc_847 N_A_1128_47#_M1022_g N_VGND_c_1638_n 0.00366111f $X=8.165 $Y=0.445 $X2=0
+ $Y2=0
cc_848 N_A_1128_47#_M1014_d N_VGND_c_1646_n 0.00285894f $X=5.64 $Y=0.235 $X2=0
+ $Y2=0
cc_849 N_A_1128_47#_M1022_g N_VGND_c_1646_n 0.00694048f $X=8.165 $Y=0.445 $X2=0
+ $Y2=0
cc_850 N_A_1128_47#_c_1275_n N_VGND_c_1646_n 0.0157978f $X=6.485 $Y=0.395 $X2=0
+ $Y2=0
cc_851 N_A_1128_47#_c_1275_n A_1237_47# 0.00726387f $X=6.485 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_852 N_A_1128_47#_c_1267_n A_1237_47# 0.00153033f $X=6.57 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_853 N_VPWR_c_1370_n N_A_436_413#_M1000_d 0.0027906f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_854 N_VPWR_c_1372_n N_A_436_413#_c_1526_n 0.0166788f $X=1.855 $Y=2.34 $X2=0
+ $Y2=0
cc_855 N_VPWR_c_1382_n N_A_436_413#_c_1526_n 0.0166511f $X=3.99 $Y=2.72 $X2=0
+ $Y2=0
cc_856 N_VPWR_c_1370_n N_A_436_413#_c_1526_n 0.00548998f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_857 N_VPWR_c_1370_n N_A_649_413#_M1004_d 0.00497477f $X=9.89 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_858 N_VPWR_c_1370_n N_A_649_413#_M1023_d 0.00230036f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_859 N_VPWR_c_1382_n N_A_649_413#_c_1558_n 0.00730735f $X=3.99 $Y=2.72 $X2=0
+ $Y2=0
cc_860 N_VPWR_c_1370_n N_A_649_413#_c_1558_n 0.00287341f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_861 N_VPWR_c_1373_n N_A_649_413#_c_1559_n 0.0209399f $X=4.155 $Y=2.29 $X2=0
+ $Y2=0
cc_862 N_VPWR_c_1382_n N_A_649_413#_c_1559_n 0.00434397f $X=3.99 $Y=2.72 $X2=0
+ $Y2=0
cc_863 N_VPWR_c_1388_n N_A_649_413#_c_1559_n 0.00330997f $X=5.005 $Y=2.72 $X2=0
+ $Y2=0
cc_864 N_VPWR_c_1370_n N_A_649_413#_c_1559_n 0.00597125f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_865 N_VPWR_c_1373_n N_A_649_413#_c_1561_n 0.0102921f $X=4.155 $Y=2.29 $X2=0
+ $Y2=0
cc_866 N_VPWR_c_1374_n N_A_649_413#_c_1561_n 0.010735f $X=5.24 $Y=2.34 $X2=0
+ $Y2=0
cc_867 N_VPWR_c_1388_n N_A_649_413#_c_1561_n 0.00730735f $X=5.005 $Y=2.72 $X2=0
+ $Y2=0
cc_868 N_VPWR_c_1370_n N_A_649_413#_c_1561_n 0.00287341f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_869 N_VPWR_c_1370_n A_1330_413# 0.0017642f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_870 N_VPWR_c_1370_n N_Q_M1002_s 0.00300692f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_871 N_VPWR_c_1379_n N_Q_c_1601_n 0.0401623f $X=9.835 $Y=1.96 $X2=0 $Y2=0
cc_872 N_VPWR_c_1390_n N_Q_c_1601_n 0.0169389f $X=9.75 $Y=2.72 $X2=0 $Y2=0
cc_873 N_VPWR_c_1370_n N_Q_c_1601_n 0.010932f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_874 N_VPWR_M1012_d Q 0.00398456f $X=9.69 $Y=1.485 $X2=0 $Y2=0
cc_875 N_VPWR_c_1379_n Q 0.0136682f $X=9.835 $Y=1.96 $X2=0 $Y2=0
cc_876 N_A_436_413#_c_1534_n N_VGND_c_1630_n 0.0110402f $X=2.33 $Y=0.39 $X2=0
+ $Y2=0
cc_877 N_A_436_413#_c_1534_n N_VGND_c_1641_n 0.01815f $X=2.33 $Y=0.39 $X2=0
+ $Y2=0
cc_878 N_A_436_413#_M1008_d N_VGND_c_1646_n 0.00280585f $X=2.19 $Y=0.235 $X2=0
+ $Y2=0
cc_879 N_A_436_413#_c_1534_n N_VGND_c_1646_n 0.0145599f $X=2.33 $Y=0.39 $X2=0
+ $Y2=0
cc_880 Q N_VGND_M1026_s 0.00315665f $X=9.79 $Y=0.765 $X2=0 $Y2=0
cc_881 Q N_VGND_c_1633_n 0.00703777f $X=9.79 $Y=0.765 $X2=0 $Y2=0
cc_882 Q N_VGND_c_1634_n 0.00131872f $X=9.79 $Y=0.765 $X2=0 $Y2=0
cc_883 Q N_VGND_c_1635_n 0.012101f $X=9.79 $Y=0.765 $X2=0 $Y2=0
cc_884 N_Q_c_1600_n N_VGND_c_1642_n 0.0227501f $X=9.365 $Y=0.39 $X2=0 $Y2=0
cc_885 Q N_VGND_c_1642_n 0.00250268f $X=9.79 $Y=0.765 $X2=0 $Y2=0
cc_886 N_Q_M1016_d N_VGND_c_1646_n 0.00305741f $X=9.18 $Y=0.235 $X2=0 $Y2=0
cc_887 N_Q_c_1600_n N_VGND_c_1646_n 0.0142238f $X=9.365 $Y=0.39 $X2=0 $Y2=0
cc_888 Q N_VGND_c_1646_n 0.00802519f $X=9.79 $Y=0.765 $X2=0 $Y2=0
cc_889 N_VGND_c_1646_n A_642_47# 0.0129748f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24
cc_890 N_VGND_c_1646_n A_805_47# 0.00196784f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24
cc_891 N_VGND_c_1646_n A_1237_47# 0.00285227f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24
cc_892 N_VGND_c_1646_n A_1542_47# 0.0028237f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24
