* File: sky130_fd_sc_hdll__nor2_8.pex.spice
* Created: Wed Sep  2 08:39:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR2_8%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 70 71 76
r140 71 72 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.805 $Y=1.202
+ $X2=3.83 $Y2=1.202
r141 69 71 17.6821 $w=3.68e-07 $l=1.35e-07 $layer=POLY_cond $X=3.67 $Y=1.202
+ $X2=3.805 $Y2=1.202
r142 69 70 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=3.67
+ $Y=1.16 $X2=3.67 $Y2=1.16
r143 67 69 43.8777 $w=3.68e-07 $l=3.35e-07 $layer=POLY_cond $X=3.335 $Y=1.202
+ $X2=3.67 $Y2=1.202
r144 66 67 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.31 $Y=1.202
+ $X2=3.335 $Y2=1.202
r145 65 66 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=2.865 $Y=1.202
+ $X2=3.31 $Y2=1.202
r146 64 65 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.84 $Y=1.202
+ $X2=2.865 $Y2=1.202
r147 63 64 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.84 $Y2=1.202
r148 62 63 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.37 $Y=1.202
+ $X2=2.395 $Y2=1.202
r149 61 62 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=2.37 $Y2=1.202
r150 60 61 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.9 $Y=1.202
+ $X2=1.925 $Y2=1.202
r151 59 60 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.9 $Y2=1.202
r152 58 59 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r153 57 58 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.43 $Y2=1.202
r154 56 57 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r155 55 76 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=0.6 $Y=1.175 $X2=0.69
+ $Y2=1.175
r156 54 56 47.1522 $w=3.68e-07 $l=3.6e-07 $layer=POLY_cond $X=0.6 $Y=1.202
+ $X2=0.96 $Y2=1.202
r157 54 55 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r158 52 54 11.1332 $w=3.68e-07 $l=8.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.6 $Y2=1.202
r159 51 52 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r160 49 70 162.482 $w=1.98e-07 $l=2.93e-06 $layer=LI1_cond $X=0.74 $Y=1.175
+ $X2=3.67 $Y2=1.175
r161 49 76 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=0.74 $Y=1.175
+ $X2=0.69 $Y2=1.175
r162 46 72 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=1.202
r163 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=0.56
r164 43 71 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.202
r165 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.985
r166 40 67 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.202
r167 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.985
r168 37 66 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=1.202
r169 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=0.56
r170 34 65 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.202
r171 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.985
r172 31 64 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=1.202
r173 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=0.56
r174 28 63 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.202
r175 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r176 25 62 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=1.202
r177 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=0.56
r178 22 61 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r179 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r180 19 60 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.9 $Y2=1.202
r181 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.9 $Y2=0.56
r182 16 59 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r183 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r184 13 58 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r185 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r186 10 57 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r187 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r188 7 56 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r189 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=0.56
r190 4 52 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r191 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r192 1 51 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r193 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_8%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 68 71 76
r139 71 72 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=7.565 $Y=1.202
+ $X2=7.59 $Y2=1.202
r140 70 71 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=7.095 $Y=1.202
+ $X2=7.565 $Y2=1.202
r141 69 70 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=7.07 $Y=1.202
+ $X2=7.095 $Y2=1.202
r142 67 69 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=7.055 $Y=1.202
+ $X2=7.07 $Y2=1.202
r143 67 68 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=7.055
+ $Y=1.16 $X2=7.055 $Y2=1.16
r144 65 67 56.3207 $w=3.68e-07 $l=4.3e-07 $layer=POLY_cond $X=6.625 $Y=1.202
+ $X2=7.055 $Y2=1.202
r145 64 65 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.6 $Y=1.202
+ $X2=6.625 $Y2=1.202
r146 63 64 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=6.155 $Y=1.202
+ $X2=6.6 $Y2=1.202
r147 62 63 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.13 $Y=1.202
+ $X2=6.155 $Y2=1.202
r148 61 62 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=5.685 $Y=1.202
+ $X2=6.13 $Y2=1.202
r149 60 61 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.66 $Y=1.202
+ $X2=5.685 $Y2=1.202
r150 59 60 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=5.215 $Y=1.202
+ $X2=5.66 $Y2=1.202
r151 58 59 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.19 $Y=1.202
+ $X2=5.215 $Y2=1.202
r152 57 58 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=4.745 $Y=1.202
+ $X2=5.19 $Y2=1.202
r153 56 57 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.72 $Y=1.202
+ $X2=4.745 $Y2=1.202
r154 55 76 51.5727 $w=1.98e-07 $l=9.3e-07 $layer=LI1_cond $X=4.375 $Y=1.175
+ $X2=5.305 $Y2=1.175
r155 54 56 45.1875 $w=3.68e-07 $l=3.45e-07 $layer=POLY_cond $X=4.375 $Y=1.202
+ $X2=4.72 $Y2=1.202
r156 54 55 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=4.375
+ $Y=1.16 $X2=4.375 $Y2=1.16
r157 52 54 13.0978 $w=3.68e-07 $l=1e-07 $layer=POLY_cond $X=4.275 $Y=1.202
+ $X2=4.375 $Y2=1.202
r158 51 52 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.25 $Y=1.202
+ $X2=4.275 $Y2=1.202
r159 49 68 95.6591 $w=1.98e-07 $l=1.725e-06 $layer=LI1_cond $X=5.33 $Y=1.175
+ $X2=7.055 $Y2=1.175
r160 49 76 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=5.33 $Y=1.175
+ $X2=5.305 $Y2=1.175
r161 46 72 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.59 $Y=0.995
+ $X2=7.59 $Y2=1.202
r162 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.59 $Y=0.995
+ $X2=7.59 $Y2=0.56
r163 43 71 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.565 $Y=1.41
+ $X2=7.565 $Y2=1.202
r164 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.565 $Y=1.41
+ $X2=7.565 $Y2=1.985
r165 40 70 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.095 $Y=1.41
+ $X2=7.095 $Y2=1.202
r166 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.095 $Y=1.41
+ $X2=7.095 $Y2=1.985
r167 37 69 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.07 $Y=0.995
+ $X2=7.07 $Y2=1.202
r168 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.07 $Y=0.995
+ $X2=7.07 $Y2=0.56
r169 34 65 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.625 $Y=1.41
+ $X2=6.625 $Y2=1.202
r170 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.625 $Y=1.41
+ $X2=6.625 $Y2=1.985
r171 31 64 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.6 $Y=0.995
+ $X2=6.6 $Y2=1.202
r172 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.6 $Y=0.995
+ $X2=6.6 $Y2=0.56
r173 28 63 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.155 $Y=1.41
+ $X2=6.155 $Y2=1.202
r174 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.155 $Y=1.41
+ $X2=6.155 $Y2=1.985
r175 25 62 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.13 $Y=0.995
+ $X2=6.13 $Y2=1.202
r176 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.13 $Y=0.995
+ $X2=6.13 $Y2=0.56
r177 22 61 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.685 $Y=1.41
+ $X2=5.685 $Y2=1.202
r178 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.685 $Y=1.41
+ $X2=5.685 $Y2=1.985
r179 19 60 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.66 $Y=0.995
+ $X2=5.66 $Y2=1.202
r180 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.66 $Y=0.995
+ $X2=5.66 $Y2=0.56
r181 16 59 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.202
r182 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.985
r183 13 58 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.202
r184 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r185 10 57 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.202
r186 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.985
r187 7 56 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.72 $Y=0.995
+ $X2=4.72 $Y2=1.202
r188 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.72 $Y=0.995
+ $X2=4.72 $Y2=0.56
r189 4 52 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.202
r190 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.985
r191 1 51 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.25 $Y=0.995
+ $X2=4.25 $Y2=1.202
r192 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.25 $Y=0.995
+ $X2=4.25 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_8%A_27_297# 1 2 3 4 5 6 7 8 9 28 30 32 36 38
+ 42 44 48 50 52 53 54 58 60 64 66 70 72 76 81 83 85 90 91 92
r103 74 76 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.8 $Y=2.295
+ $X2=7.8 $Y2=1.96
r104 73 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.985 $Y=2.38
+ $X2=6.86 $Y2=2.38
r105 72 74 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.675 $Y=2.38
+ $X2=7.8 $Y2=2.295
r106 72 73 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.675 $Y=2.38
+ $X2=6.985 $Y2=2.38
r107 68 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.86 $Y=2.295
+ $X2=6.86 $Y2=2.38
r108 68 70 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.86 $Y=2.295
+ $X2=6.86 $Y2=1.96
r109 67 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.045 $Y=2.38
+ $X2=5.92 $Y2=2.38
r110 66 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.735 $Y=2.38
+ $X2=6.86 $Y2=2.38
r111 66 67 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.735 $Y=2.38
+ $X2=6.045 $Y2=2.38
r112 62 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.295
+ $X2=5.92 $Y2=2.38
r113 62 64 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.92 $Y=2.295
+ $X2=5.92 $Y2=1.96
r114 61 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.105 $Y=2.38
+ $X2=4.98 $Y2=2.38
r115 60 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.795 $Y=2.38
+ $X2=5.92 $Y2=2.38
r116 60 61 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.795 $Y=2.38
+ $X2=5.105 $Y2=2.38
r117 56 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.295
+ $X2=4.98 $Y2=2.38
r118 56 58 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.98 $Y=2.295
+ $X2=4.98 $Y2=1.96
r119 55 89 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.165 $Y=2.38
+ $X2=4.04 $Y2=2.38
r120 54 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=2.38
+ $X2=4.98 $Y2=2.38
r121 54 55 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.855 $Y=2.38
+ $X2=4.165 $Y2=2.38
r122 53 89 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.295
+ $X2=4.04 $Y2=2.38
r123 52 87 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=1.56
r124 52 53 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=2.295
r125 51 85 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.225 $Y=1.56
+ $X2=3.1 $Y2=1.56
r126 50 87 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.915 $Y=1.56
+ $X2=4.04 $Y2=1.56
r127 50 51 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=3.915 $Y=1.56
+ $X2=3.225 $Y2=1.56
r128 46 85 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.1 $Y=1.665
+ $X2=3.1 $Y2=1.56
r129 46 48 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.1 $Y=1.665
+ $X2=3.1 $Y2=2.3
r130 45 83 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=1.56
+ $X2=2.16 $Y2=1.56
r131 44 85 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.975 $Y=1.56
+ $X2=3.1 $Y2=1.56
r132 44 45 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=2.975 $Y=1.56
+ $X2=2.285 $Y2=1.56
r133 40 83 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.56
r134 40 42 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=2.3
r135 39 81 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=1.56
+ $X2=1.22 $Y2=1.56
r136 38 83 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=1.56
+ $X2=2.16 $Y2=1.56
r137 38 39 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=1.56
+ $X2=1.345 $Y2=1.56
r138 34 81 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.56
r139 34 36 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=2.3
r140 33 79 4.31179 $w=2.1e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=1.56
+ $X2=0.247 $Y2=1.56
r141 32 81 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.56
+ $X2=1.22 $Y2=1.56
r142 32 33 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.56
+ $X2=0.405 $Y2=1.56
r143 28 79 2.86543 $w=3.15e-07 $l=1.05e-07 $layer=LI1_cond $X=0.247 $Y=1.665
+ $X2=0.247 $Y2=1.56
r144 28 30 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=0.247 $Y=1.665
+ $X2=0.247 $Y2=2.3
r145 9 76 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.655
+ $Y=1.485 $X2=7.8 $Y2=1.96
r146 8 70 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.715
+ $Y=1.485 $X2=6.86 $Y2=1.96
r147 7 64 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.775
+ $Y=1.485 $X2=5.92 $Y2=1.96
r148 6 58 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.835
+ $Y=1.485 $X2=4.98 $Y2=1.96
r149 5 89 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.485 $X2=4.04 $Y2=2.3
r150 5 87 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.485 $X2=4.04 $Y2=1.62
r151 4 85 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=1.62
r152 4 48 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=2.3
r153 3 83 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.62
r154 3 42 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.3
r155 2 81 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r156 2 36 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r157 1 79 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r158 1 30 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_8%VPWR 1 2 3 4 17 19 23 25 29 31 35 37 44 45
+ 48 51 54 57
r99 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r100 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r101 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r102 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r103 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r104 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r105 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r106 44 45 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r107 42 45 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=8.05 $Y2=2.72
r108 42 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r109 41 44 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=8.05 $Y2=2.72
r110 41 42 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r111 39 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.695 $Y=2.72
+ $X2=3.57 $Y2=2.72
r112 39 41 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.695 $Y=2.72
+ $X2=3.91 $Y2=2.72
r113 37 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r114 33 57 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=2.635
+ $X2=3.57 $Y2=2.72
r115 33 35 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.57 $Y=2.635
+ $X2=3.57 $Y2=2
r116 32 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.63 $Y2=2.72
r117 31 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.445 $Y=2.72
+ $X2=3.57 $Y2=2.72
r118 31 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.445 $Y=2.72
+ $X2=2.755 $Y2=2.72
r119 27 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=2.635
+ $X2=2.63 $Y2=2.72
r120 27 29 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.63 $Y=2.635
+ $X2=2.63 $Y2=2
r121 26 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.69 $Y2=2.72
r122 25 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=2.63 $Y2=2.72
r123 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=1.815 $Y2=2.72
r124 21 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=2.72
r125 21 23 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=2
r126 20 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r127 19 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=1.69 $Y2=2.72
r128 19 20 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=0.875 $Y2=2.72
r129 15 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r130 15 17 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2
r131 4 35 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=2
r132 3 29 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=2
r133 2 23 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=2
r134 1 17 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_8%Y 1 2 3 4 5 6 7 8 9 10 11 12 39 41 42 45 47
+ 51 53 57 59 63 67 69 70 71 75 79 81 83 87 91 93 95 99 101 102 103 104 105 106
+ 107 108 110 113
r223 112 113 9.45786 $w=7.33e-07 $l=5.4e-07 $layer=LI1_cond $X=7.742 $Y=0.905
+ $X2=7.742 $Y2=1.445
r224 110 112 13.3681 $w=3.76e-07 $l=5.85837e-07 $layer=LI1_cond $X=7.33 $Y=0.49
+ $X2=7.742 $Y2=0.905
r225 97 113 2.37703 $w=4.07e-07 $l=3.24731e-07 $layer=LI1_cond $X=7.33 $Y=1.615
+ $X2=7.615 $Y2=1.53
r226 97 99 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=7.33 $Y=1.615
+ $X2=7.33 $Y2=1.62
r227 96 107 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.555 $Y=0.815
+ $X2=6.365 $Y2=0.815
r228 95 110 10.305 $w=3.76e-07 $l=4.18927e-07 $layer=LI1_cond $X=7.115 $Y=0.815
+ $X2=7.33 $Y2=0.49
r229 95 96 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=7.115 $Y=0.815
+ $X2=6.555 $Y2=0.815
r230 94 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.515 $Y=1.53
+ $X2=6.39 $Y2=1.53
r231 93 113 4.61444 $w=1.7e-07 $l=4.1e-07 $layer=LI1_cond $X=7.205 $Y=1.53
+ $X2=7.615 $Y2=1.53
r232 93 94 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.205 $Y=1.53
+ $X2=6.515 $Y2=1.53
r233 89 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.615
+ $X2=6.39 $Y2=1.53
r234 89 91 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.39 $Y=1.615
+ $X2=6.39 $Y2=1.62
r235 85 107 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.365 $Y=0.725
+ $X2=6.365 $Y2=0.815
r236 85 87 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.365 $Y=0.725
+ $X2=6.365 $Y2=0.39
r237 84 105 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.615 $Y=0.815
+ $X2=5.425 $Y2=0.815
r238 83 107 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.175 $Y=0.815
+ $X2=6.365 $Y2=0.815
r239 83 84 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.175 $Y=0.815
+ $X2=5.615 $Y2=0.815
r240 82 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.575 $Y=1.53
+ $X2=5.45 $Y2=1.53
r241 81 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.265 $Y=1.53
+ $X2=6.39 $Y2=1.53
r242 81 82 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.265 $Y=1.53
+ $X2=5.575 $Y2=1.53
r243 77 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=1.615
+ $X2=5.45 $Y2=1.53
r244 77 79 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.45 $Y=1.615
+ $X2=5.45 $Y2=1.62
r245 73 105 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.425 $Y=0.725
+ $X2=5.425 $Y2=0.815
r246 73 75 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.425 $Y=0.725
+ $X2=5.425 $Y2=0.39
r247 72 104 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.675 $Y=0.815
+ $X2=4.485 $Y2=0.815
r248 71 105 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.235 $Y=0.815
+ $X2=5.425 $Y2=0.815
r249 71 72 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.235 $Y=0.815
+ $X2=4.675 $Y2=0.815
r250 69 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.325 $Y=1.53
+ $X2=5.45 $Y2=1.53
r251 69 70 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.325 $Y=1.53
+ $X2=4.635 $Y2=1.53
r252 65 70 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.51 $Y=1.615
+ $X2=4.635 $Y2=1.53
r253 65 67 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.51 $Y=1.615
+ $X2=4.51 $Y2=1.62
r254 61 104 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.485 $Y=0.725
+ $X2=4.485 $Y2=0.815
r255 61 63 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.485 $Y=0.725
+ $X2=4.485 $Y2=0.39
r256 60 103 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.735 $Y=0.815
+ $X2=3.545 $Y2=0.815
r257 59 104 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.295 $Y=0.815
+ $X2=4.485 $Y2=0.815
r258 59 60 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.295 $Y=0.815
+ $X2=3.735 $Y2=0.815
r259 55 103 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.545 $Y2=0.815
r260 55 57 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.545 $Y2=0.39
r261 54 102 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.795 $Y=0.815
+ $X2=2.605 $Y2=0.815
r262 53 103 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=3.545 $Y2=0.815
r263 53 54 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=2.795 $Y2=0.815
r264 49 102 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.605 $Y2=0.815
r265 49 51 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.605 $Y2=0.39
r266 48 101 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=0.815
+ $X2=1.665 $Y2=0.815
r267 47 102 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=2.605 $Y2=0.815
r268 47 48 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=1.855 $Y2=0.815
r269 43 101 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.815
r270 43 45 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.39
r271 41 101 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=1.665 $Y2=0.815
r272 41 42 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=0.915 $Y2=0.815
r273 37 42 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.815
r274 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r275 12 99 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=7.185
+ $Y=1.485 $X2=7.33 $Y2=1.62
r276 11 91 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.245
+ $Y=1.485 $X2=6.39 $Y2=1.62
r277 10 79 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.305
+ $Y=1.485 $X2=5.45 $Y2=1.62
r278 9 67 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.365
+ $Y=1.485 $X2=4.51 $Y2=1.62
r279 8 110 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.145
+ $Y=0.235 $X2=7.33 $Y2=0.39
r280 7 87 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.205
+ $Y=0.235 $X2=6.39 $Y2=0.39
r281 6 75 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.265
+ $Y=0.235 $X2=5.45 $Y2=0.39
r282 5 63 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.325
+ $Y=0.235 $X2=4.51 $Y2=0.39
r283 4 57 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.235 $X2=3.57 $Y2=0.39
r284 3 51 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.235 $X2=2.63 $Y2=0.39
r285 2 45 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r286 1 39 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_8%VGND 1 2 3 4 5 6 7 8 9 28 30 32 36 40 44 48
+ 52 56 60 64 67 68 70 71 73 74 76 77 79 80 82 83 84 85 86 87 113 118
r146 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r147 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r148 110 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r149 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r150 107 110 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r151 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r152 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r153 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r154 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r155 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r156 98 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r157 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r158 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r159 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r160 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r161 92 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.15 $Y2=0
r162 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r163 89 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r164 89 91 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=2.07 $Y2=0
r165 87 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r166 87 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r167 85 109 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.59 $Y2=0
r168 85 86 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.715 $Y=0 $X2=7.86
+ $Y2=0
r169 84 112 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=8.005 $Y=0 $X2=8.05
+ $Y2=0
r170 84 86 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=8.005 $Y=0 $X2=7.86
+ $Y2=0
r171 82 106 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.775 $Y=0
+ $X2=6.67 $Y2=0
r172 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.86
+ $Y2=0
r173 81 109 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.945 $Y=0
+ $X2=7.59 $Y2=0
r174 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.945 $Y=0 $X2=6.86
+ $Y2=0
r175 79 103 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0
+ $X2=5.75 $Y2=0
r176 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.92
+ $Y2=0
r177 78 106 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.005 $Y=0
+ $X2=6.67 $Y2=0
r178 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0 $X2=5.92
+ $Y2=0
r179 76 100 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=4.83 $Y2=0
r180 76 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.98
+ $Y2=0
r181 75 103 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.065 $Y=0
+ $X2=5.75 $Y2=0
r182 75 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=4.98
+ $Y2=0
r183 73 97 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.955 $Y=0 $X2=3.91
+ $Y2=0
r184 73 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0 $X2=4.04
+ $Y2=0
r185 72 100 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.125 $Y=0
+ $X2=4.83 $Y2=0
r186 72 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0 $X2=4.04
+ $Y2=0
r187 70 94 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=2.99
+ $Y2=0
r188 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.1
+ $Y2=0
r189 69 97 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=3.91 $Y2=0
r190 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.1
+ $Y2=0
r191 67 91 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r192 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.16
+ $Y2=0
r193 66 94 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.99 $Y2=0
r194 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r195 62 86 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.86 $Y=0.085
+ $X2=7.86 $Y2=0
r196 62 64 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=7.86 $Y=0.085
+ $X2=7.86 $Y2=0.39
r197 58 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.86 $Y=0.085
+ $X2=6.86 $Y2=0
r198 58 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.86 $Y=0.085
+ $X2=6.86 $Y2=0.39
r199 54 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r200 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.39
r201 50 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r202 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.39
r203 46 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r204 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.39
r205 42 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0
r206 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0.39
r207 38 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r208 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.39
r209 34 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r210 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r211 33 115 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r212 32 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r213 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=0.365 $Y2=0
r214 28 115 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r215 28 30 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r216 9 64 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.665
+ $Y=0.235 $X2=7.8 $Y2=0.39
r217 8 60 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.675
+ $Y=0.235 $X2=6.86 $Y2=0.39
r218 7 56 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.735
+ $Y=0.235 $X2=5.92 $Y2=0.39
r219 6 52 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.795
+ $Y=0.235 $X2=4.98 $Y2=0.39
r220 5 48 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.39
r221 4 44 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.39
r222 3 40 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.16 $Y2=0.39
r223 2 36 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
r224 1 30 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

