* File: sky130_fd_sc_hdll__inv_8.pex.spice
* Created: Thu Aug 27 19:09:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INV_8%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 50 51 52 53 54 80 81
r160 81 82 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.95 $Y=1.202
+ $X2=3.975 $Y2=1.202
r161 79 81 30.7799 $w=3.68e-07 $l=2.35e-07 $layer=POLY_cond $X=3.715 $Y=1.202
+ $X2=3.95 $Y2=1.202
r162 79 80 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.715
+ $Y=1.16 $X2=3.715 $Y2=1.16
r163 77 79 30.7799 $w=3.68e-07 $l=2.35e-07 $layer=POLY_cond $X=3.48 $Y=1.202
+ $X2=3.715 $Y2=1.202
r164 76 77 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.455 $Y=1.202
+ $X2=3.48 $Y2=1.202
r165 75 76 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=3.01 $Y=1.202
+ $X2=3.455 $Y2=1.202
r166 74 75 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.985 $Y=1.202
+ $X2=3.01 $Y2=1.202
r167 73 74 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=2.54 $Y=1.202
+ $X2=2.985 $Y2=1.202
r168 72 73 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.515 $Y=1.202
+ $X2=2.54 $Y2=1.202
r169 71 72 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=2.07 $Y=1.202
+ $X2=2.515 $Y2=1.202
r170 70 71 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.045 $Y=1.202
+ $X2=2.07 $Y2=1.202
r171 69 70 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=1.6 $Y=1.202
+ $X2=2.045 $Y2=1.202
r172 68 69 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.575 $Y=1.202
+ $X2=1.6 $Y2=1.202
r173 67 68 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=1.13 $Y=1.202
+ $X2=1.575 $Y2=1.202
r174 66 67 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.105 $Y=1.202
+ $X2=1.13 $Y2=1.202
r175 64 66 27.5054 $w=3.68e-07 $l=2.1e-07 $layer=POLY_cond $X=0.895 $Y=1.202
+ $X2=1.105 $Y2=1.202
r176 64 65 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=0.895
+ $Y=1.16 $X2=0.895 $Y2=1.16
r177 62 64 30.7799 $w=3.68e-07 $l=2.35e-07 $layer=POLY_cond $X=0.66 $Y=1.202
+ $X2=0.895 $Y2=1.202
r178 61 62 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.635 $Y=1.202
+ $X2=0.66 $Y2=1.202
r179 54 80 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=3.45 $Y=1.2
+ $X2=3.715 $Y2=1.2
r180 53 54 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.99 $Y=1.2 $X2=3.45
+ $Y2=1.2
r181 52 53 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=1.2 $X2=2.99
+ $Y2=1.2
r182 51 52 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.07 $Y=1.2 $X2=2.53
+ $Y2=1.2
r183 50 51 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.61 $Y=1.2 $X2=2.07
+ $Y2=1.2
r184 49 50 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=1.61
+ $Y2=1.2
r185 49 65 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.15 $Y=1.2
+ $X2=0.895 $Y2=1.2
r186 46 82 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.975 $Y=0.995
+ $X2=3.975 $Y2=1.202
r187 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.975 $Y=0.995
+ $X2=3.975 $Y2=0.56
r188 43 81 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.95 $Y=1.41
+ $X2=3.95 $Y2=1.202
r189 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.95 $Y=1.41
+ $X2=3.95 $Y2=1.985
r190 40 77 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.48 $Y=1.41
+ $X2=3.48 $Y2=1.202
r191 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.48 $Y=1.41
+ $X2=3.48 $Y2=1.985
r192 37 76 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.455 $Y=0.995
+ $X2=3.455 $Y2=1.202
r193 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.455 $Y=0.995
+ $X2=3.455 $Y2=0.56
r194 34 75 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.01 $Y=1.41
+ $X2=3.01 $Y2=1.202
r195 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.01 $Y=1.41
+ $X2=3.01 $Y2=1.985
r196 31 74 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.985 $Y=0.995
+ $X2=2.985 $Y2=1.202
r197 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.985 $Y=0.995
+ $X2=2.985 $Y2=0.56
r198 28 73 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.54 $Y=1.41
+ $X2=2.54 $Y2=1.202
r199 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.54 $Y=1.41
+ $X2=2.54 $Y2=1.985
r200 25 72 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.515 $Y=0.995
+ $X2=2.515 $Y2=1.202
r201 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.515 $Y=0.995
+ $X2=2.515 $Y2=0.56
r202 22 71 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.07 $Y=1.41
+ $X2=2.07 $Y2=1.202
r203 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.07 $Y=1.41
+ $X2=2.07 $Y2=1.985
r204 19 70 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.045 $Y=0.995
+ $X2=2.045 $Y2=1.202
r205 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.045 $Y=0.995
+ $X2=2.045 $Y2=0.56
r206 16 69 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.6 $Y=1.41 $X2=1.6
+ $Y2=1.202
r207 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.6 $Y=1.41
+ $X2=1.6 $Y2=1.985
r208 13 68 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.575 $Y=0.995
+ $X2=1.575 $Y2=1.202
r209 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.575 $Y=0.995
+ $X2=1.575 $Y2=0.56
r210 10 67 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.13 $Y=1.41
+ $X2=1.13 $Y2=1.202
r211 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.13 $Y=1.41
+ $X2=1.13 $Y2=1.985
r212 7 66 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.105 $Y=0.995
+ $X2=1.105 $Y2=1.202
r213 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.105 $Y=0.995
+ $X2=1.105 $Y2=0.56
r214 4 62 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.66 $Y=1.41
+ $X2=0.66 $Y2=1.202
r215 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.66 $Y=1.41
+ $X2=0.66 $Y2=1.985
r216 1 61 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=1.202
r217 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_8%VPWR 1 2 3 4 5 16 18 22 26 30 32 34 37 38 40
+ 41 43 44 45 57 66
c72 5 0 1.55756e-19 $X=4.04 $Y=1.485
c73 1 0 1.5644e-19 $X=0.3 $Y=1.485
r74 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r75 60 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r76 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r77 57 65 4.3205 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=4.1 $Y=2.72 $X2=4.35
+ $Y2=2.72
r78 57 59 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.1 $Y=2.72 $X2=3.91
+ $Y2=2.72
r79 56 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r80 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r81 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r82 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r83 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r84 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r85 47 62 3.91904 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=2.72
+ $X2=0.255 $Y2=2.72
r86 47 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.51 $Y=2.72 $X2=1.15
+ $Y2=2.72
r87 45 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r88 45 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r89 43 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.16 $Y=2.72
+ $X2=2.99 $Y2=2.72
r90 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=2.72
+ $X2=3.245 $Y2=2.72
r91 42 59 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=3.91 $Y2=2.72
r92 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=3.245 $Y2=2.72
r93 40 52 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=2.72 $X2=2.07
+ $Y2=2.72
r94 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=2.72
+ $X2=2.305 $Y2=2.72
r95 39 55 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.39 $Y=2.72 $X2=2.99
+ $Y2=2.72
r96 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=2.72
+ $X2=2.305 $Y2=2.72
r97 37 49 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.28 $Y=2.72
+ $X2=1.15 $Y2=2.72
r98 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=2.72
+ $X2=1.365 $Y2=2.72
r99 36 52 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=2.07 $Y2=2.72
r100 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=1.365 $Y2=2.72
r101 32 65 3.19717 $w=3e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.25 $Y=2.635
+ $X2=4.35 $Y2=2.72
r102 32 34 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=4.25 $Y=2.635
+ $X2=4.25 $Y2=2
r103 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=2.635
+ $X2=3.245 $Y2=2.72
r104 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.245 $Y=2.635
+ $X2=3.245 $Y2=2
r105 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=2.635
+ $X2=2.305 $Y2=2.72
r106 24 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.305 $Y=2.635
+ $X2=2.305 $Y2=2
r107 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=2.635
+ $X2=1.365 $Y2=2.72
r108 20 22 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.365 $Y=2.635
+ $X2=1.365 $Y2=2
r109 16 62 3.25818 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.382 $Y=2.635
+ $X2=0.255 $Y2=2.72
r110 16 18 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.382 $Y=2.635
+ $X2=0.382 $Y2=2
r111 5 34 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.04
+ $Y=1.485 $X2=4.185 $Y2=2
r112 4 30 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.1
+ $Y=1.485 $X2=3.245 $Y2=2
r113 3 26 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.16
+ $Y=1.485 $X2=2.305 $Y2=2
r114 2 22 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=1.485 $X2=1.365 $Y2=2
r115 1 18 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.3
+ $Y=1.485 $X2=0.425 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_8%Y 1 2 3 4 5 6 7 8 25 26 27 28 31 35 37 39 43
+ 47 49 51 55 59 61 63 67 71 73 75 79 81 82 84 85 87 88 90 93 94
c185 94 0 1.55756e-19 $X=4.38 $Y=1.19
c186 93 0 1.5644e-19 $X=0.23 $Y=1.19
r187 92 94 10.9842 $w=3.18e-07 $l=3.05e-07 $layer=LI1_cond $X=4.345 $Y=1.495
+ $X2=4.345 $Y2=1.19
r188 91 94 10.2639 $w=3.18e-07 $l=2.85e-07 $layer=LI1_cond $X=4.345 $Y=0.905
+ $X2=4.345 $Y2=1.19
r189 78 93 10.1883 $w=3.43e-07 $l=3.05e-07 $layer=LI1_cond $X=0.257 $Y=1.495
+ $X2=0.257 $Y2=1.19
r190 77 93 9.52018 $w=3.43e-07 $l=2.85e-07 $layer=LI1_cond $X=0.257 $Y=0.905
+ $X2=0.257 $Y2=1.19
r191 76 90 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.88 $Y=1.58
+ $X2=3.69 $Y2=1.58
r192 75 92 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=4.185 $Y=1.58
+ $X2=4.345 $Y2=1.495
r193 75 76 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.185 $Y=1.58
+ $X2=3.88 $Y2=1.58
r194 74 88 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.88 $Y=0.81
+ $X2=3.69 $Y2=0.81
r195 73 91 7.40893 $w=1.9e-07 $l=2.0199e-07 $layer=LI1_cond $X=4.185 $Y=0.81
+ $X2=4.345 $Y2=0.905
r196 73 74 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=4.185 $Y=0.81
+ $X2=3.88 $Y2=0.81
r197 69 90 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=1.665
+ $X2=3.69 $Y2=1.58
r198 69 71 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.69 $Y=1.665
+ $X2=3.69 $Y2=2.34
r199 65 88 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.69 $Y=0.715
+ $X2=3.69 $Y2=0.81
r200 65 67 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.69 $Y=0.715
+ $X2=3.69 $Y2=0.38
r201 64 87 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.94 $Y=1.58
+ $X2=2.75 $Y2=1.58
r202 63 90 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.5 $Y=1.58 $X2=3.69
+ $Y2=1.58
r203 63 64 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.5 $Y=1.58
+ $X2=2.94 $Y2=1.58
r204 62 85 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=2.94 $Y=0.81
+ $X2=2.75 $Y2=0.81
r205 61 88 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.5 $Y=0.81 $X2=3.69
+ $Y2=0.81
r206 61 62 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=3.5 $Y=0.81 $X2=2.94
+ $Y2=0.81
r207 57 87 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=1.665
+ $X2=2.75 $Y2=1.58
r208 57 59 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.75 $Y=1.665
+ $X2=2.75 $Y2=2.34
r209 53 85 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.75 $Y=0.715
+ $X2=2.75 $Y2=0.81
r210 53 55 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.75 $Y=0.715
+ $X2=2.75 $Y2=0.38
r211 52 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2 $Y=1.58 $X2=1.81
+ $Y2=1.58
r212 51 87 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.56 $Y=1.58
+ $X2=2.75 $Y2=1.58
r213 51 52 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.56 $Y=1.58 $X2=2
+ $Y2=1.58
r214 50 82 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=2 $Y=0.81 $X2=1.81
+ $Y2=0.81
r215 49 85 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=2.56 $Y=0.81
+ $X2=2.75 $Y2=0.81
r216 49 50 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=2.56 $Y=0.81 $X2=2
+ $Y2=0.81
r217 45 84 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=1.665
+ $X2=1.81 $Y2=1.58
r218 45 47 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.81 $Y=1.665
+ $X2=1.81 $Y2=2.34
r219 41 82 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.81 $Y=0.715
+ $X2=1.81 $Y2=0.81
r220 41 43 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.81 $Y=0.715
+ $X2=1.81 $Y2=0.38
r221 40 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.06 $Y=1.58
+ $X2=0.87 $Y2=1.58
r222 39 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=1.58
+ $X2=1.81 $Y2=1.58
r223 39 40 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.62 $Y=1.58
+ $X2=1.06 $Y2=1.58
r224 38 79 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=1.06 $Y=0.81
+ $X2=0.87 $Y2=0.81
r225 37 82 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.81
+ $X2=1.81 $Y2=0.81
r226 37 38 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=1.62 $Y=0.81
+ $X2=1.06 $Y2=0.81
r227 33 81 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=1.665
+ $X2=0.87 $Y2=1.58
r228 33 35 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.87 $Y=1.665
+ $X2=0.87 $Y2=2.34
r229 29 79 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=0.87 $Y=0.715
+ $X2=0.87 $Y2=0.81
r230 29 31 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.87 $Y=0.715
+ $X2=0.87 $Y2=0.38
r231 28 78 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.43 $Y=1.58
+ $X2=0.257 $Y2=1.495
r232 27 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.68 $Y=1.58
+ $X2=0.87 $Y2=1.58
r233 27 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.68 $Y=1.58
+ $X2=0.43 $Y2=1.58
r234 26 77 7.58838 $w=1.9e-07 $l=2.15323e-07 $layer=LI1_cond $X=0.43 $Y=0.81
+ $X2=0.257 $Y2=0.905
r235 25 79 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=0.68 $Y=0.81
+ $X2=0.87 $Y2=0.81
r236 25 26 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=0.68 $Y=0.81
+ $X2=0.43 $Y2=0.81
r237 8 90 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=1.485 $X2=3.715 $Y2=1.66
r238 8 71 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=1.485 $X2=3.715 $Y2=2.34
r239 7 87 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.485 $X2=2.775 $Y2=1.66
r240 7 59 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.485 $X2=2.775 $Y2=2.34
r241 6 84 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.69
+ $Y=1.485 $X2=1.835 $Y2=1.66
r242 6 47 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.69
+ $Y=1.485 $X2=1.835 $Y2=2.34
r243 5 81 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.75
+ $Y=1.485 $X2=0.895 $Y2=1.66
r244 5 35 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.75
+ $Y=1.485 $X2=0.895 $Y2=2.34
r245 4 67 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.53
+ $Y=0.235 $X2=3.715 $Y2=0.38
r246 3 55 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.59
+ $Y=0.235 $X2=2.775 $Y2=0.38
r247 2 43 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.65
+ $Y=0.235 $X2=1.835 $Y2=0.38
r248 1 31 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=0.71
+ $Y=0.235 $X2=0.895 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_8%VGND 1 2 3 4 5 16 18 22 26 30 32 34 37 38 40
+ 41 43 44 45 57 66
r82 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r83 60 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r84 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r85 57 65 4.36388 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=4.1 $Y=0 $X2=4.35
+ $Y2=0
r86 57 59 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.1 $Y=0 $X2=3.91
+ $Y2=0
r87 56 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r88 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r89 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r90 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r91 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r92 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r93 47 62 3.91904 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.255
+ $Y2=0
r94 47 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=1.15
+ $Y2=0
r95 45 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r96 45 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r97 43 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.16 $Y=0 $X2=2.99
+ $Y2=0
r98 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=0 $X2=3.245
+ $Y2=0
r99 42 59 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.91
+ $Y2=0
r100 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.245
+ $Y2=0
r101 40 52 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.07
+ $Y2=0
r102 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.305
+ $Y2=0
r103 39 55 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.99
+ $Y2=0
r104 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.305
+ $Y2=0
r105 37 49 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.15
+ $Y2=0
r106 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.365
+ $Y2=0
r107 36 52 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=2.07
+ $Y2=0
r108 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.365
+ $Y2=0
r109 32 65 3.19436 $w=3.05e-07 $l=1.33918e-07 $layer=LI1_cond $X=4.252 $Y=0.085
+ $X2=4.35 $Y2=0
r110 32 34 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=4.252 $Y=0.085
+ $X2=4.252 $Y2=0.38
r111 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=0.085
+ $X2=3.245 $Y2=0
r112 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.245 $Y=0.085
+ $X2=3.245 $Y2=0.38
r113 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0
r114 24 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0.38
r115 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=0.085
+ $X2=1.365 $Y2=0
r116 20 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.365 $Y=0.085
+ $X2=1.365 $Y2=0.38
r117 16 62 3.25818 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.382 $Y=0.085
+ $X2=0.255 $Y2=0
r118 16 18 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.382 $Y=0.085
+ $X2=0.382 $Y2=0.38
r119 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.05
+ $Y=0.235 $X2=4.185 $Y2=0.38
r120 4 30 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.235 $X2=3.245 $Y2=0.38
r121 3 26 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.235 $X2=2.305 $Y2=0.38
r122 2 22 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.18
+ $Y=0.235 $X2=1.365 $Y2=0.38
r123 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.3
+ $Y=0.235 $X2=0.425 $Y2=0.38
.ends

