* NGSPICE file created from sky130_fd_sc_hdll__nand4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
M1000 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=1.0157e+12p ps=8.13e+06u
M1001 VGND A_N a_40_93# VNB nshort w=420000u l=150000u
+  ad=2.6875e+11p pd=2.18e+06u as=1.323e+11p ps=1.47e+06u
M1002 VPWR A_N a_40_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 VPWR a_40_93# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_431_47# B a_334_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=2.1775e+11p ps=1.97e+06u
M1005 Y a_40_93# a_431_47# VNB nshort w=650000u l=150000u
+  ad=2.925e+11p pd=2.2e+06u as=0p ps=0u
M1006 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_334_47# C a_251_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u
M1008 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_251_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

