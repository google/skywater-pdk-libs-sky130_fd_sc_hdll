* NGSPICE file created from sky130_fd_sc_hdll__a22oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=5.8e+11p ps=5.16e+06u
M1001 Y B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=1.755e+11p ps=1.84e+06u
M1002 a_117_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_411_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1004 VPWR A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1005 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_411_47# VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1007 a_119_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

