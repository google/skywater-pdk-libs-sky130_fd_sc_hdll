* File: sky130_fd_sc_hdll__inv_1.pex.spice
* Created: Wed Sep  2 08:32:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INV_1%A 1 3 4 6 7 11 15
r20 11 15 11.2843 $w=2.38e-07 $l=2.35e-07 $layer=LI1_cond $X=0.485 $Y=1.195
+ $X2=0.25 $Y2=1.195
r21 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=1.16 $X2=0.485 $Y2=1.16
r22 7 15 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=0.245 $Y=1.195
+ $X2=0.25 $Y2=1.195
r23 4 10 40.0415 $w=4.22e-07 $l=2.33345e-07 $layer=POLY_cond $X=0.725 $Y=0.995
+ $X2=0.56 $Y2=1.16
r24 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.725 $Y=0.995
+ $X2=0.725 $Y2=0.56
r25 1 10 44.7429 $w=4.22e-07 $l=3.1225e-07 $layer=POLY_cond $X=0.7 $Y=1.41
+ $X2=0.56 $Y2=1.16
r26 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.7 $Y=1.41 $X2=0.7
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_1%VPWR 1 6 11 12 13 20 21
r14 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r15 13 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r16 13 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r17 11 16 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.34 $Y=2.72
+ $X2=0.23 $Y2=2.72
r18 11 12 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.34 $Y=2.72
+ $X2=0.445 $Y2=2.72
r19 10 20 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.55 $Y=2.72 $X2=1.15
+ $Y2=2.72
r20 10 12 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.55 $Y=2.72
+ $X2=0.445 $Y2=2.72
r21 6 9 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=0.445 $Y=1.66
+ $X2=0.445 $Y2=2.34
r22 4 12 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.445 $Y=2.635
+ $X2=0.445 $Y2=2.72
r23 4 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.445 $Y=2.635
+ $X2=0.445 $Y2=2.34
r24 1 9 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.34
+ $Y=1.485 $X2=0.465 $Y2=2.34
r25 1 6 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.34
+ $Y=1.485 $X2=0.465 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_1%Y 1 2 9 13 16 17 26
r19 26 27 3.30959 $w=5.13e-07 $l=4.5e-08 $layer=LI1_cond $X=1.027 $Y=1.53
+ $X2=1.027 $Y2=1.485
r20 17 30 2.55473 $w=5.13e-07 $l=1.1e-07 $layer=LI1_cond $X=1.027 $Y=1.55
+ $X2=1.027 $Y2=1.66
r21 17 26 0.464496 $w=5.13e-07 $l=2e-08 $layer=LI1_cond $X=1.027 $Y=1.55
+ $X2=1.027 $Y2=1.53
r22 17 27 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=1.14 $Y=1.465
+ $X2=1.14 $Y2=1.485
r23 16 17 10.9283 $w=2.88e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=1.19
+ $X2=1.14 $Y2=1.465
r24 15 16 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.14 $Y=0.885
+ $X2=1.14 $Y2=1.19
r25 13 15 13.5285 $w=5.13e-07 $l=4.85e-07 $layer=LI1_cond $X=1.027 $Y=0.4
+ $X2=1.027 $Y2=0.885
r26 7 30 1.90444 $w=5.13e-07 $l=8.2e-08 $layer=LI1_cond $X=1.027 $Y=1.742
+ $X2=1.027 $Y2=1.66
r27 7 9 13.8884 $w=5.13e-07 $l=5.98e-07 $layer=LI1_cond $X=1.027 $Y=1.742
+ $X2=1.027 $Y2=2.34
r28 2 30 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.79
+ $Y=1.485 $X2=0.935 $Y2=1.66
r29 2 9 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.79
+ $Y=1.485 $X2=0.935 $Y2=2.34
r30 1 13 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.8
+ $Y=0.235 $X2=0.935 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_1%VGND 1 6 9 10 11 18 19
r14 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r15 11 19 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r16 11 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r17 9 14 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.23
+ $Y2=0
r18 9 10 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.435
+ $Y2=0
r19 8 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=1.15
+ $Y2=0
r20 8 10 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.435
+ $Y2=0
r21 4 10 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.435 $Y=0.085
+ $X2=0.435 $Y2=0
r22 4 6 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.435 $Y=0.085
+ $X2=0.435 $Y2=0.4
r23 1 6 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.34
+ $Y=0.235 $X2=0.465 $Y2=0.4
.ends

