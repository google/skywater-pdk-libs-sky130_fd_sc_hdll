* File: sky130_fd_sc_hdll__a2bb2oi_2.pxi.spice
* Created: Thu Aug 27 18:55:09 2020
* 
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%B1 N_B1_c_81_n N_B1_M1005_g N_B1_c_82_n
+ N_B1_M1010_g N_B1_c_83_n N_B1_M1009_g N_B1_c_84_n N_B1_M1011_g N_B1_c_89_n
+ N_B1_c_85_n B1 B1 PM_SKY130_FD_SC_HDLL__A2BB2OI_2%B1
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%B2 N_B2_c_155_n N_B2_M1003_g N_B2_c_159_n
+ N_B2_M1000_g N_B2_c_160_n N_B2_M1016_g N_B2_c_156_n N_B2_M1019_g B2
+ N_B2_c_157_n N_B2_c_158_n B2 PM_SKY130_FD_SC_HDLL__A2BB2OI_2%B2
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_455_21# N_A_455_21#_M1004_d
+ N_A_455_21#_M1006_s N_A_455_21#_M1001_s N_A_455_21#_c_199_n
+ N_A_455_21#_M1014_g N_A_455_21#_c_206_n N_A_455_21#_M1002_g
+ N_A_455_21#_c_200_n N_A_455_21#_M1015_g N_A_455_21#_c_207_n
+ N_A_455_21#_M1007_g N_A_455_21#_c_201_n N_A_455_21#_c_208_n
+ N_A_455_21#_c_217_p N_A_455_21#_c_202_n N_A_455_21#_c_223_p
+ N_A_455_21#_c_271_p N_A_455_21#_c_203_n N_A_455_21#_c_204_n
+ N_A_455_21#_c_205_n PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_455_21#
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A1_N N_A1_N_c_300_n N_A1_N_M1004_g
+ N_A1_N_c_304_n N_A1_N_M1012_g N_A1_N_c_305_n N_A1_N_M1018_g N_A1_N_c_301_n
+ N_A1_N_M1013_g A1_N N_A1_N_c_303_n A1_N PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A1_N
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A2_N N_A2_N_c_345_n N_A2_N_M1006_g
+ N_A2_N_c_349_n N_A2_N_M1001_g N_A2_N_c_350_n N_A2_N_M1008_g N_A2_N_c_346_n
+ N_A2_N_M1017_g A2_N N_A2_N_c_348_n A2_N PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A2_N
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_27_297# N_A_27_297#_M1005_s
+ N_A_27_297#_M1000_d N_A_27_297#_M1009_s N_A_27_297#_M1007_d
+ N_A_27_297#_c_410_p N_A_27_297#_c_387_n N_A_27_297#_c_382_n
+ N_A_27_297#_c_406_p N_A_27_297#_c_392_n N_A_27_297#_c_383_n
+ N_A_27_297#_c_409_p N_A_27_297#_c_401_n N_A_27_297#_c_395_n
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%VPWR N_VPWR_M1005_d N_VPWR_M1016_s
+ N_VPWR_M1012_s N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n N_VPWR_c_429_n
+ N_VPWR_c_430_n N_VPWR_c_431_n VPWR N_VPWR_c_432_n N_VPWR_c_433_n
+ N_VPWR_c_425_n N_VPWR_c_435_n N_VPWR_c_436_n
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%Y N_Y_M1003_d N_Y_M1014_s N_Y_M1002_s
+ N_Y_c_503_n N_Y_c_511_n N_Y_c_504_n N_Y_c_505_n Y Y
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_2%Y
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_695_297# N_A_695_297#_M1012_d
+ N_A_695_297#_M1018_d N_A_695_297#_M1008_d N_A_695_297#_c_552_n
+ N_A_695_297#_c_553_n N_A_695_297#_c_554_n N_A_695_297#_c_576_n
+ N_A_695_297#_c_578_n N_A_695_297#_c_548_n N_A_695_297#_c_549_n
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_695_297#
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%VGND N_VGND_M1010_s N_VGND_M1011_s
+ N_VGND_M1015_d N_VGND_M1013_s N_VGND_M1017_d N_VGND_c_583_n N_VGND_c_584_n
+ N_VGND_c_585_n N_VGND_c_586_n N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n
+ N_VGND_c_590_n N_VGND_c_591_n VGND N_VGND_c_592_n N_VGND_c_593_n
+ N_VGND_c_594_n N_VGND_c_595_n N_VGND_c_596_n N_VGND_c_597_n
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_2%VGND
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_119_47# N_A_119_47#_M1010_d
+ N_A_119_47#_M1019_s N_A_119_47#_c_669_n N_A_119_47#_c_668_n
+ N_A_119_47#_c_673_n PM_SKY130_FD_SC_HDLL__A2BB2OI_2%A_119_47#
cc_1 VNB N_B1_c_81_n 0.0326155f $X=-0.325 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_B1_c_82_n 0.0218895f $X=-0.325 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_B1_c_83_n 0.0219112f $X=-0.325 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_4 VNB N_B1_c_84_n 0.0166622f $X=-0.325 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_B1_c_85_n 0.00408992f $X=-0.325 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_6 VNB B1 0.014715f $X=-0.325 $Y=-0.24 $X2=0.31 $Y2=1.105
cc_7 VNB N_B2_c_155_n 0.0170715f $X=-0.325 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_B2_c_156_n 0.0173947f $X=-0.325 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_9 VNB N_B2_c_157_n 0.00161932f $X=-0.325 $Y=-0.24 $X2=1.905 $Y2=1.53
cc_10 VNB N_B2_c_158_n 0.0364654f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_455_21#_c_199_n 0.0164563f $X=-0.325 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_12 VNB N_A_455_21#_c_200_n 0.0193466f $X=-0.325 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_13 VNB N_A_455_21#_c_201_n 0.00498466f $X=-0.325 $Y=-0.24 $X2=0.31 $Y2=1.445
cc_14 VNB N_A_455_21#_c_202_n 0.00630004f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_455_21#_c_203_n 0.00593529f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_455_21#_c_204_n 0.00262404f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_455_21#_c_205_n 0.0597903f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A1_N_c_300_n 0.0216159f $X=-0.325 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_19 VNB N_A1_N_c_301_n 0.0169382f $X=-0.325 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_20 VNB A1_N 0.0092683f $X=-0.325 $Y=-0.24 $X2=1.715 $Y2=1.53
cc_21 VNB N_A1_N_c_303_n 0.0381985f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A2_N_c_345_n 0.0169338f $X=-0.325 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_23 VNB N_A2_N_c_346_n 0.0223809f $X=-0.325 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_24 VNB A2_N 0.0113855f $X=-0.325 $Y=-0.24 $X2=1.715 $Y2=1.53
cc_25 VNB N_A2_N_c_348_n 0.0442958f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_425_n 0.250759f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_503_n 0.0106741f $X=-0.325 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_28 VNB N_Y_c_504_n 0.00259728f $X=-0.325 $Y=-0.24 $X2=1.905 $Y2=1.53
cc_29 VNB N_Y_c_505_n 8.10088e-19 $X=-0.325 $Y=-0.24 $X2=0.31 $Y2=1.105
cc_30 VNB Y 8.7147e-19 $X=-0.325 $Y=-0.24 $X2=0.31 $Y2=1.445
cc_31 VNB N_VGND_c_583_n 0.0110494f $X=-0.325 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_32 VNB N_VGND_c_584_n 0.00651836f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_585_n 0.00467156f $X=-0.325 $Y=-0.24 $X2=0.31 $Y2=1.445
cc_34 VNB N_VGND_c_586_n 0.00467156f $X=-0.325 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_35 VNB N_VGND_c_587_n 0.00800025f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_588_n 0.0192911f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_589_n 0.00323964f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_590_n 0.0201171f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_591_n 0.00326991f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_592_n 0.0407218f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_593_n 0.0153494f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_594_n 0.306718f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_595_n 0.00323964f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_596_n 0.0200006f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_597_n 0.0208884f $X=-0.325 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_119_47#_c_668_n 0.00320511f $X=-0.325 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_47 VPB N_B1_c_81_n 0.0301878f $X=-0.325 $Y=1.305 $X2=0.495 $Y2=1.41
cc_48 VPB N_B1_c_83_n 0.0247986f $X=-0.325 $Y=1.305 $X2=1.905 $Y2=1.41
cc_49 VPB N_B1_c_89_n 0.00884837f $X=-0.325 $Y=1.305 $X2=1.715 $Y2=1.53
cc_50 VPB N_B1_c_85_n 0.00300004f $X=-0.325 $Y=1.305 $X2=1.88 $Y2=1.16
cc_51 VPB B1 0.0149906f $X=-0.325 $Y=1.305 $X2=0.31 $Y2=1.105
cc_52 VPB N_B2_c_159_n 0.0159975f $X=-0.325 $Y=1.305 $X2=0.52 $Y2=0.995
cc_53 VPB N_B2_c_160_n 0.0159964f $X=-0.325 $Y=1.305 $X2=1.905 $Y2=1.41
cc_54 VPB N_B2_c_158_n 0.0193497f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_455_21#_c_206_n 0.0161002f $X=-0.325 $Y=1.305 $X2=1.715 $Y2=1.53
cc_56 VPB N_A_455_21#_c_207_n 0.0189026f $X=-0.325 $Y=1.305 $X2=1.905 $Y2=1.53
cc_57 VPB N_A_455_21#_c_208_n 0.0195882f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_455_21#_c_203_n 0.00766108f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_455_21#_c_205_n 0.0303659f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A1_N_c_304_n 0.0201091f $X=-0.325 $Y=1.305 $X2=0.52 $Y2=0.995
cc_61 VPB N_A1_N_c_305_n 0.0160057f $X=-0.325 $Y=1.305 $X2=1.905 $Y2=1.41
cc_62 VPB N_A1_N_c_303_n 0.0206567f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A2_N_c_349_n 0.0160057f $X=-0.325 $Y=1.305 $X2=0.52 $Y2=0.995
cc_64 VPB N_A2_N_c_350_n 0.0202816f $X=-0.325 $Y=1.305 $X2=1.905 $Y2=1.41
cc_65 VPB N_A2_N_c_348_n 0.0235665f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_297#_c_382_n 0.00692367f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_297#_c_383_n 0.00148837f $X=-0.325 $Y=1.305 $X2=0.375 $Y2=1.16
cc_68 VPB N_VPWR_c_426_n 0.00516582f $X=-0.325 $Y=1.305 $X2=1.93 $Y2=0.56
cc_69 VPB N_VPWR_c_427_n 0.0195604f $X=-0.325 $Y=1.305 $X2=0.64 $Y2=1.53
cc_70 VPB N_VPWR_c_428_n 0.00516582f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_429_n 0.00516582f $X=-0.325 $Y=1.305 $X2=0.31 $Y2=1.445
cc_72 VPB N_VPWR_c_430_n 0.0537613f $X=-0.325 $Y=1.305 $X2=0.435 $Y2=1.16
cc_73 VPB N_VPWR_c_431_n 0.00478242f $X=-0.325 $Y=1.305 $X2=0.41 $Y2=1.16
cc_74 VPB N_VPWR_c_432_n 0.0190625f $X=-0.325 $Y=1.305 $X2=0.375 $Y2=1.16
cc_75 VPB N_VPWR_c_433_n 0.0466991f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_425_n 0.0677482f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_435_n 0.00478242f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_436_n 0.00478242f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_695_297#_c_548_n 0.00594067f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_695_297#_c_549_n 0.00164584f $X=-0.325 $Y=1.305 $X2=0 $Y2=0
cc_81 N_B1_c_82_n N_B2_c_155_n 0.0165288f $X=0.52 $Y=0.995 $X2=-0.325 $Y2=-0.24
cc_82 N_B1_c_81_n N_B2_c_159_n 0.037155f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B1_c_89_n N_B2_c_159_n 0.0113958f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_84 B1 N_B2_c_159_n 9.98963e-19 $X=0.31 $Y=1.105 $X2=0 $Y2=0
cc_85 N_B1_c_83_n N_B2_c_160_n 0.0371417f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B1_c_89_n N_B2_c_160_n 0.0122112f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_87 N_B1_c_85_n N_B2_c_160_n 0.00101445f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_88 N_B1_c_84_n N_B2_c_156_n 0.0223996f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B1_c_81_n N_B2_c_157_n 7.33201e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B1_c_83_n N_B2_c_157_n 2.06373e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B1_c_89_n N_B2_c_157_n 0.0416942f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_92 N_B1_c_85_n N_B2_c_157_n 0.0117433f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_93 B1 N_B2_c_157_n 0.0151943f $X=0.31 $Y=1.105 $X2=0 $Y2=0
cc_94 N_B1_c_81_n N_B2_c_158_n 0.0165288f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B1_c_83_n N_B2_c_158_n 0.0264727f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B1_c_89_n N_B2_c_158_n 0.00803891f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_97 N_B1_c_85_n N_B2_c_158_n 0.00478003f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_98 B1 N_B2_c_158_n 0.00413013f $X=0.31 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B1_c_84_n N_A_455_21#_c_199_n 0.0261773f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B1_c_83_n N_A_455_21#_c_206_n 0.0212009f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B1_c_85_n N_A_455_21#_c_206_n 0.00170023f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B1_c_83_n N_A_455_21#_c_205_n 0.0262229f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B1_c_85_n N_A_455_21#_c_205_n 0.00284749f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_104 B1 N_A_27_297#_M1005_s 0.00284151f $X=0.31 $Y=1.105 $X2=-0.325 $Y2=-0.24
cc_105 N_B1_c_89_n N_A_27_297#_M1000_d 0.00187091f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_106 N_B1_c_85_n N_A_27_297#_M1009_s 0.00197697f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_107 N_B1_c_81_n N_A_27_297#_c_387_n 0.0112216f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_108 N_B1_c_89_n N_A_27_297#_c_387_n 0.02495f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_109 B1 N_A_27_297#_c_387_n 0.0134161f $X=0.31 $Y=1.105 $X2=0 $Y2=0
cc_110 N_B1_c_81_n N_A_27_297#_c_382_n 3.96914e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_111 B1 N_A_27_297#_c_382_n 0.0188817f $X=0.31 $Y=1.105 $X2=0 $Y2=0
cc_112 N_B1_c_83_n N_A_27_297#_c_392_n 0.0115302f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B1_c_89_n N_A_27_297#_c_392_n 0.0218268f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_114 N_B1_c_85_n N_A_27_297#_c_392_n 0.020493f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_115 N_B1_c_89_n N_A_27_297#_c_395_n 0.0143191f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_116 N_B1_c_89_n N_VPWR_M1005_d 0.00187547f $X=1.715 $Y=1.53 $X2=-0.325
+ $Y2=-0.24
cc_117 N_B1_c_89_n N_VPWR_M1016_s 0.00172342f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_118 N_B1_c_85_n N_VPWR_M1016_s 7.76441e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B1_c_81_n N_VPWR_c_426_n 0.00300743f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B1_c_83_n N_VPWR_c_428_n 0.00300743f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B1_c_83_n N_VPWR_c_430_n 0.00702461f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_122 N_B1_c_81_n N_VPWR_c_432_n 0.00702461f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B1_c_81_n N_VPWR_c_425_n 0.00787122f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B1_c_83_n N_VPWR_c_425_n 0.006985f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B1_c_83_n N_Y_c_503_n 0.00437722f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_126 N_B1_c_84_n N_Y_c_503_n 0.0126966f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B1_c_89_n N_Y_c_503_n 0.00852213f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_128 N_B1_c_85_n N_Y_c_503_n 0.0294729f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_129 N_B1_c_84_n N_Y_c_511_n 8.5962e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B1_c_83_n Y 0.00163786f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_131 N_B1_c_85_n Y 0.0250172f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_132 N_B1_c_81_n N_VGND_c_584_n 0.00176179f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_133 N_B1_c_82_n N_VGND_c_584_n 0.00614111f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_134 B1 N_VGND_c_584_n 0.0145468f $X=0.31 $Y=1.105 $X2=0 $Y2=0
cc_135 N_B1_c_84_n N_VGND_c_585_n 0.00268723f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B1_c_82_n N_VGND_c_592_n 0.00463936f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B1_c_84_n N_VGND_c_592_n 0.00437852f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_138 N_B1_c_82_n N_VGND_c_594_n 0.00876414f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B1_c_84_n N_VGND_c_594_n 0.00605933f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B1_c_82_n N_A_119_47#_c_669_n 0.00382935f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B1_c_82_n N_A_119_47#_c_668_n 0.00725663f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B1_c_89_n N_A_119_47#_c_668_n 0.00646027f $X=1.715 $Y=1.53 $X2=0 $Y2=0
cc_143 B1 N_A_119_47#_c_668_n 0.0101175f $X=0.31 $Y=1.105 $X2=0 $Y2=0
cc_144 N_B2_c_159_n N_A_27_297#_c_387_n 0.011229f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B2_c_160_n N_A_27_297#_c_392_n 0.011229f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B2_c_159_n N_VPWR_c_426_n 0.00300743f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B2_c_159_n N_VPWR_c_427_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B2_c_160_n N_VPWR_c_427_n 0.00702461f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B2_c_160_n N_VPWR_c_428_n 0.00300743f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B2_c_159_n N_VPWR_c_425_n 0.00695979f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B2_c_160_n N_VPWR_c_425_n 0.00695979f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B2_c_156_n N_Y_c_503_n 0.0106996f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B2_c_155_n N_Y_c_504_n 0.00387597f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B2_c_157_n N_Y_c_504_n 0.0338933f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B2_c_158_n N_Y_c_504_n 0.0047334f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_156 N_B2_c_155_n N_VGND_c_592_n 0.00357877f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_157 N_B2_c_156_n N_VGND_c_592_n 0.00357877f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_158 N_B2_c_155_n N_VGND_c_594_n 0.005504f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_159 N_B2_c_156_n N_VGND_c_594_n 0.00562222f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B2_c_155_n N_A_119_47#_c_673_n 0.0112873f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B2_c_156_n N_A_119_47#_c_673_n 0.0101195f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B2_c_157_n N_A_119_47#_c_673_n 0.00310861f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_455_21#_c_201_n N_A1_N_c_300_n 0.0108074f $X=3.855 $Y=0.815
+ $X2=-0.325 $Y2=-0.24
cc_164 N_A_455_21#_c_217_p N_A1_N_c_300_n 0.0110728f $X=4.07 $Y=0.39 $X2=-0.325
+ $Y2=-0.24
cc_165 N_A_455_21#_c_203_n N_A1_N_c_300_n 0.0025955f $X=3.08 $Y=1.16 $X2=-0.325
+ $Y2=-0.24
cc_166 N_A_455_21#_c_204_n N_A1_N_c_300_n 0.00119564f $X=4.045 $Y=0.815
+ $X2=-0.325 $Y2=-0.24
cc_167 N_A_455_21#_c_208_n N_A1_N_c_304_n 0.0137819f $X=4.885 $Y=1.53 $X2=0
+ $Y2=0
cc_168 N_A_455_21#_c_208_n N_A1_N_c_305_n 0.011867f $X=4.885 $Y=1.53 $X2=0 $Y2=0
cc_169 N_A_455_21#_c_202_n N_A1_N_c_301_n 0.0106151f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_170 N_A_455_21#_c_223_p N_A1_N_c_301_n 5.32212e-19 $X=5.01 $Y=0.39 $X2=0
+ $Y2=0
cc_171 N_A_455_21#_c_201_n A1_N 0.0281469f $X=3.855 $Y=0.815 $X2=0 $Y2=0
cc_172 N_A_455_21#_c_208_n A1_N 0.0719255f $X=4.885 $Y=1.53 $X2=0 $Y2=0
cc_173 N_A_455_21#_c_202_n A1_N 0.0167344f $X=4.795 $Y=0.815 $X2=0 $Y2=0
cc_174 N_A_455_21#_c_203_n A1_N 0.0161058f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_455_21#_c_204_n A1_N 0.0307352f $X=4.045 $Y=0.815 $X2=0 $Y2=0
cc_176 N_A_455_21#_c_205_n A1_N 8.32501e-19 $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_177 N_A_455_21#_c_208_n N_A1_N_c_303_n 0.00798993f $X=4.885 $Y=1.53 $X2=0
+ $Y2=0
cc_178 N_A_455_21#_c_203_n N_A1_N_c_303_n 0.00330529f $X=3.08 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_A_455_21#_c_204_n N_A1_N_c_303_n 0.00486271f $X=4.045 $Y=0.815 $X2=0
+ $Y2=0
cc_180 N_A_455_21#_c_205_n N_A1_N_c_303_n 0.00689536f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_181 N_A_455_21#_c_202_n N_A2_N_c_345_n 0.0103143f $X=4.795 $Y=0.815
+ $X2=-0.325 $Y2=-0.24
cc_182 N_A_455_21#_c_223_p N_A2_N_c_345_n 0.00644736f $X=5.01 $Y=0.39 $X2=-0.325
+ $Y2=-0.24
cc_183 N_A_455_21#_c_208_n N_A2_N_c_349_n 0.0160252f $X=4.885 $Y=1.53 $X2=0
+ $Y2=0
cc_184 N_A_455_21#_c_208_n N_A2_N_c_350_n 6.32657e-19 $X=4.885 $Y=1.53 $X2=0
+ $Y2=0
cc_185 N_A_455_21#_c_202_n N_A2_N_c_346_n 2.15189e-19 $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_186 N_A_455_21#_c_208_n A2_N 0.0317474f $X=4.885 $Y=1.53 $X2=0 $Y2=0
cc_187 N_A_455_21#_c_202_n A2_N 0.0358714f $X=4.795 $Y=0.815 $X2=0 $Y2=0
cc_188 N_A_455_21#_c_208_n N_A2_N_c_348_n 0.00737024f $X=4.885 $Y=1.53 $X2=0
+ $Y2=0
cc_189 N_A_455_21#_c_202_n N_A2_N_c_348_n 0.00486271f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_190 N_A_455_21#_c_203_n N_A_27_297#_M1007_d 0.00307358f $X=3.08 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_A_455_21#_c_206_n N_A_27_297#_c_383_n 0.0137768f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_455_21#_c_207_n N_A_27_297#_c_383_n 0.0137768f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_193 N_A_455_21#_c_203_n N_A_27_297#_c_401_n 0.0121898f $X=3.08 $Y=1.16 $X2=0
+ $Y2=0
cc_194 N_A_455_21#_c_205_n N_A_27_297#_c_401_n 0.00180987f $X=2.845 $Y=1.202
+ $X2=0 $Y2=0
cc_195 N_A_455_21#_c_208_n N_VPWR_M1012_s 0.00187547f $X=4.885 $Y=1.53 $X2=0
+ $Y2=0
cc_196 N_A_455_21#_c_206_n N_VPWR_c_430_n 0.00429453f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_197 N_A_455_21#_c_207_n N_VPWR_c_430_n 0.00429453f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_198 N_A_455_21#_M1001_s N_VPWR_c_425_n 0.00232895f $X=4.865 $Y=1.485 $X2=0
+ $Y2=0
cc_199 N_A_455_21#_c_206_n N_VPWR_c_425_n 0.00609021f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_200 N_A_455_21#_c_207_n N_VPWR_c_425_n 0.00734734f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_201 N_A_455_21#_c_199_n N_Y_c_503_n 0.0122977f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_455_21#_c_199_n N_Y_c_511_n 0.00653191f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_455_21#_c_200_n N_Y_c_511_n 0.011462f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_455_21#_c_199_n N_Y_c_505_n 0.00224457f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_455_21#_c_200_n N_Y_c_505_n 0.00302768f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_455_21#_c_203_n N_Y_c_505_n 0.00923935f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_455_21#_c_199_n Y 0.00257069f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_455_21#_c_206_n Y 0.0109332f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_455_21#_c_200_n Y 0.00235369f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_455_21#_c_207_n Y 0.0158268f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_455_21#_c_203_n Y 0.0382509f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_455_21#_c_205_n Y 0.0353491f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_213 N_A_455_21#_c_208_n N_A_695_297#_M1012_d 0.00290685f $X=4.885 $Y=1.53
+ $X2=-0.325 $Y2=-0.24
cc_214 N_A_455_21#_c_208_n N_A_695_297#_M1018_d 0.00187091f $X=4.885 $Y=1.53
+ $X2=0 $Y2=0
cc_215 N_A_455_21#_c_208_n N_A_695_297#_c_552_n 0.0372789f $X=4.885 $Y=1.53
+ $X2=0 $Y2=0
cc_216 N_A_455_21#_c_208_n N_A_695_297#_c_553_n 0.0143191f $X=4.885 $Y=1.53
+ $X2=0 $Y2=0
cc_217 N_A_455_21#_M1001_s N_A_695_297#_c_554_n 0.00352392f $X=4.865 $Y=1.485
+ $X2=0 $Y2=0
cc_218 N_A_455_21#_c_271_p N_A_695_297#_c_554_n 0.0134104f $X=5.01 $Y=1.62 $X2=0
+ $Y2=0
cc_219 N_A_455_21#_c_208_n N_A_695_297#_c_548_n 0.00209545f $X=4.885 $Y=1.53
+ $X2=0 $Y2=0
cc_220 N_A_455_21#_c_208_n N_A_695_297#_c_549_n 0.0173294f $X=4.885 $Y=1.53
+ $X2=0 $Y2=0
cc_221 N_A_455_21#_c_201_n N_VGND_M1015_d 0.00591147f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_222 N_A_455_21#_c_203_n N_VGND_M1015_d 0.00458064f $X=3.08 $Y=1.16 $X2=0
+ $Y2=0
cc_223 N_A_455_21#_c_202_n N_VGND_M1013_s 0.00162089f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_224 N_A_455_21#_c_199_n N_VGND_c_585_n 0.00268723f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_455_21#_c_202_n N_VGND_c_586_n 0.0122559f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_226 N_A_455_21#_c_202_n N_VGND_c_587_n 0.00133683f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_227 N_A_455_21#_c_201_n N_VGND_c_588_n 0.00198695f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_228 N_A_455_21#_c_217_p N_VGND_c_588_n 0.0231806f $X=4.07 $Y=0.39 $X2=0 $Y2=0
cc_229 N_A_455_21#_c_202_n N_VGND_c_588_n 0.00254521f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_230 N_A_455_21#_c_202_n N_VGND_c_590_n 0.00198695f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_231 N_A_455_21#_c_223_p N_VGND_c_590_n 0.0231806f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_232 N_A_455_21#_M1004_d N_VGND_c_594_n 0.00304143f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_233 N_A_455_21#_M1006_s N_VGND_c_594_n 0.00364931f $X=4.825 $Y=0.235 $X2=0
+ $Y2=0
cc_234 N_A_455_21#_c_199_n N_VGND_c_594_n 0.00587047f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_455_21#_c_200_n N_VGND_c_594_n 0.0110773f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_455_21#_c_201_n N_VGND_c_594_n 0.00537187f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_237 N_A_455_21#_c_217_p N_VGND_c_594_n 0.0143352f $X=4.07 $Y=0.39 $X2=0 $Y2=0
cc_238 N_A_455_21#_c_202_n N_VGND_c_594_n 0.0094839f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_239 N_A_455_21#_c_223_p N_VGND_c_594_n 0.0143352f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_240 N_A_455_21#_c_203_n N_VGND_c_594_n 7.36513e-19 $X=3.08 $Y=1.16 $X2=0
+ $Y2=0
cc_241 N_A_455_21#_c_199_n N_VGND_c_596_n 0.00423334f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A_455_21#_c_200_n N_VGND_c_596_n 0.00541359f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_455_21#_c_200_n N_VGND_c_597_n 0.00617046f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_455_21#_c_201_n N_VGND_c_597_n 0.030682f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_245 N_A_455_21#_c_203_n N_VGND_c_597_n 0.0193543f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A_455_21#_c_205_n N_VGND_c_597_n 0.00137626f $X=2.845 $Y=1.202 $X2=0
+ $Y2=0
cc_247 N_A1_N_c_301_n N_A2_N_c_345_n 0.0244072f $X=4.33 $Y=0.995 $X2=-0.325
+ $Y2=-0.24
cc_248 N_A1_N_c_305_n N_A2_N_c_349_n 0.0222872f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_249 A1_N A2_N 0.0132504f $X=4.06 $Y=1.105 $X2=0 $Y2=0
cc_250 N_A1_N_c_303_n A2_N 2.09584e-19 $X=4.305 $Y=1.202 $X2=0 $Y2=0
cc_251 A1_N N_A2_N_c_348_n 0.00164236f $X=4.06 $Y=1.105 $X2=0 $Y2=0
cc_252 N_A1_N_c_303_n N_A2_N_c_348_n 0.0244072f $X=4.305 $Y=1.202 $X2=0 $Y2=0
cc_253 N_A1_N_c_304_n N_VPWR_c_429_n 0.00300743f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A1_N_c_305_n N_VPWR_c_429_n 0.00300743f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A1_N_c_304_n N_VPWR_c_430_n 0.0053025f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A1_N_c_305_n N_VPWR_c_433_n 0.0053025f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A1_N_c_304_n N_VPWR_c_425_n 0.00818727f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A1_N_c_305_n N_VPWR_c_425_n 0.00693014f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A1_N_c_304_n N_A_695_297#_c_552_n 0.0123176f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_260 N_A1_N_c_305_n N_A_695_297#_c_552_n 0.0123176f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_261 N_A1_N_c_301_n N_VGND_c_586_n 0.00268723f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A1_N_c_300_n N_VGND_c_588_n 0.00423334f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A1_N_c_301_n N_VGND_c_588_n 0.00437852f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A1_N_c_300_n N_VGND_c_594_n 0.00728222f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A1_N_c_301_n N_VGND_c_594_n 0.00615622f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A1_N_c_300_n N_VGND_c_597_n 0.00481673f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A2_N_c_349_n N_VPWR_c_433_n 0.00429453f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A2_N_c_350_n N_VPWR_c_433_n 0.00429453f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A2_N_c_349_n N_VPWR_c_425_n 0.00609021f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A2_N_c_350_n N_VPWR_c_425_n 0.00713556f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A2_N_c_349_n N_A_695_297#_c_554_n 0.0143578f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_272 N_A2_N_c_350_n N_A_695_297#_c_554_n 0.0143578f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_273 N_A2_N_c_350_n N_A_695_297#_c_548_n 7.41963e-19 $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_274 A2_N N_A_695_297#_c_548_n 0.00647905f $X=5.08 $Y=1.105 $X2=0 $Y2=0
cc_275 N_A2_N_c_345_n N_VGND_c_586_n 0.00268723f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A2_N_c_346_n N_VGND_c_587_n 0.00483862f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_277 A2_N N_VGND_c_587_n 0.00333084f $X=5.08 $Y=1.105 $X2=0 $Y2=0
cc_278 N_A2_N_c_345_n N_VGND_c_590_n 0.00423334f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A2_N_c_346_n N_VGND_c_590_n 0.00585385f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A2_N_c_345_n N_VGND_c_594_n 0.00598581f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A2_N_c_346_n N_VGND_c_594_n 0.0118977f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A_27_297#_c_387_n N_VPWR_M1005_d 0.0037528f $X=1.075 $Y=1.87 $X2=-0.325
+ $Y2=1.305
cc_283 N_A_27_297#_c_392_n N_VPWR_M1016_s 0.00371343f $X=2.015 $Y=1.87 $X2=0
+ $Y2=0
cc_284 N_A_27_297#_c_387_n N_VPWR_c_426_n 0.0132478f $X=1.075 $Y=1.87 $X2=0
+ $Y2=0
cc_285 N_A_27_297#_c_406_p N_VPWR_c_427_n 0.0149311f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_286 N_A_27_297#_c_392_n N_VPWR_c_428_n 0.0131725f $X=2.015 $Y=1.87 $X2=0
+ $Y2=0
cc_287 N_A_27_297#_c_383_n N_VPWR_c_430_n 0.0549564f $X=2.955 $Y=2.38 $X2=0
+ $Y2=0
cc_288 N_A_27_297#_c_409_p N_VPWR_c_430_n 0.015002f $X=2.265 $Y=2.38 $X2=0 $Y2=0
cc_289 N_A_27_297#_c_410_p N_VPWR_c_432_n 0.0161853f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_290 N_A_27_297#_M1005_s N_VPWR_c_425_n 0.00226492f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_291 N_A_27_297#_M1000_d N_VPWR_c_425_n 0.00250817f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_292 N_A_27_297#_M1009_s N_VPWR_c_425_n 0.00241844f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_293 N_A_27_297#_M1007_d N_VPWR_c_425_n 0.00217519f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_294 N_A_27_297#_c_410_p N_VPWR_c_425_n 0.00955092f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_295 N_A_27_297#_c_387_n N_VPWR_c_425_n 0.0141814f $X=1.075 $Y=1.87 $X2=0
+ $Y2=0
cc_296 N_A_27_297#_c_406_p N_VPWR_c_425_n 0.00955092f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_297 N_A_27_297#_c_392_n N_VPWR_c_425_n 0.0141797f $X=2.015 $Y=1.87 $X2=0
+ $Y2=0
cc_298 N_A_27_297#_c_383_n N_VPWR_c_425_n 0.0335386f $X=2.955 $Y=2.38 $X2=0
+ $Y2=0
cc_299 N_A_27_297#_c_409_p N_VPWR_c_425_n 0.00962794f $X=2.265 $Y=2.38 $X2=0
+ $Y2=0
cc_300 N_A_27_297#_c_383_n N_Y_M1002_s 0.00352392f $X=2.955 $Y=2.38 $X2=0 $Y2=0
cc_301 N_A_27_297#_c_383_n Y 0.0160463f $X=2.955 $Y=2.38 $X2=0 $Y2=0
cc_302 N_A_27_297#_c_383_n N_A_695_297#_c_549_n 0.0100846f $X=2.955 $Y=2.38
+ $X2=0 $Y2=0
cc_303 N_A_27_297#_c_401_n N_A_695_297#_c_549_n 0.0280952f $X=3.08 $Y=1.96 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_425_n N_Y_M1002_s 0.00232895f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_305 N_VPWR_c_425_n N_A_695_297#_M1012_d 0.00226208f $X=5.75 $Y=2.72
+ $X2=-0.325 $Y2=-0.24
cc_306 N_VPWR_c_425_n N_A_695_297#_M1018_d 0.00241559f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_425_n N_A_695_297#_M1008_d 0.00303346f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_308 N_VPWR_M1012_s N_A_695_297#_c_552_n 0.00348321f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_429_n N_A_695_297#_c_552_n 0.0139299f $X=4.07 $Y=2.3 $X2=0 $Y2=0
cc_310 N_VPWR_c_430_n N_A_695_297#_c_552_n 0.00254499f $X=3.945 $Y=2.72 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_433_n N_A_695_297#_c_552_n 0.00254499f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_425_n N_A_695_297#_c_552_n 0.0103134f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_433_n N_A_695_297#_c_554_n 0.0386815f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_425_n N_A_695_297#_c_554_n 0.0239144f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_433_n N_A_695_297#_c_576_n 0.015002f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_316 N_VPWR_c_425_n N_A_695_297#_c_576_n 0.00962794f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_433_n N_A_695_297#_c_578_n 0.0162563f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_425_n N_A_695_297#_c_578_n 0.00961749f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_430_n N_A_695_297#_c_549_n 0.0161853f $X=3.945 $Y=2.72 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_425_n N_A_695_297#_c_549_n 0.00955092f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_321 N_Y_c_503_n N_VGND_M1011_s 0.00162089f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_322 N_Y_c_503_n N_VGND_c_585_n 0.0122559f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_323 N_Y_c_503_n N_VGND_c_592_n 0.00255089f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_324 N_Y_M1003_d N_VGND_c_594_n 0.00297142f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_325 N_Y_M1014_s N_VGND_c_594_n 0.0025535f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_326 N_Y_c_503_n N_VGND_c_594_n 0.0105605f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_327 N_Y_c_511_n N_VGND_c_594_n 0.0141452f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_328 N_Y_c_503_n N_VGND_c_596_n 0.00198695f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_329 N_Y_c_511_n N_VGND_c_596_n 0.0224137f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_330 N_Y_c_511_n N_VGND_c_597_n 0.0204642f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_331 N_Y_c_503_n N_A_119_47#_M1019_s 0.00253211f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_332 N_Y_c_504_n N_A_119_47#_c_668_n 0.0105775f $X=1.365 $Y=0.775 $X2=0 $Y2=0
cc_333 N_Y_M1003_d N_A_119_47#_c_673_n 0.00507817f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_334 N_Y_c_503_n N_A_119_47#_c_673_n 0.017531f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_335 N_Y_c_504_n N_A_119_47#_c_673_n 0.0205972f $X=1.365 $Y=0.775 $X2=0 $Y2=0
cc_336 N_A_695_297#_c_548_n N_VGND_c_587_n 0.00532467f $X=5.48 $Y=1.62 $X2=0
+ $Y2=0
cc_337 N_VGND_c_594_n N_A_119_47#_M1010_d 0.00215206f $X=5.75 $Y=0 $X2=-0.325
+ $Y2=-0.24
cc_338 N_VGND_c_594_n N_A_119_47#_M1019_s 0.00264825f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_c_584_n N_A_119_47#_c_669_n 0.0172916f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_340 N_VGND_c_592_n N_A_119_47#_c_669_n 0.0185904f $X=2.055 $Y=0 $X2=0 $Y2=0
cc_341 N_VGND_c_594_n N_A_119_47#_c_669_n 0.0110971f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_342 N_VGND_c_584_n N_A_119_47#_c_668_n 0.0307592f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_343 N_VGND_c_592_n N_A_119_47#_c_673_n 0.0576174f $X=2.055 $Y=0 $X2=0 $Y2=0
cc_344 N_VGND_c_594_n N_A_119_47#_c_673_n 0.0366908f $X=5.75 $Y=0 $X2=0 $Y2=0
