* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__einvn_4 A TE_B VGND VNB VPB VPWR Z
X0 Z A a_222_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_27_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_222_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X3 VGND a_27_47# a_235_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Z A a_235_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR TE_B a_222_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X6 Z A a_235_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_222_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_222_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X9 a_235_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND a_27_47# a_235_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_235_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_27_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_235_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Z A a_222_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VPWR TE_B a_222_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X16 a_222_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_235_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
