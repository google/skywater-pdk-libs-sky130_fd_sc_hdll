* File: sky130_fd_sc_hdll__nor2b_4.pex.spice
* Created: Thu Aug 27 19:16:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR2B_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 44
r78 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r79 37 39 20.0833 $w=3.72e-07 $l=1.55e-07 $layer=POLY_cond $X=1.77 $Y=1.202
+ $X2=1.925 $Y2=1.202
r80 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.77
+ $Y=1.16 $X2=1.77 $Y2=1.16
r81 35 37 40.8145 $w=3.72e-07 $l=3.15e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.77 $Y2=1.202
r82 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r83 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.43 $Y2=1.202
r84 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r85 31 44 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=0.6 $Y=1.175
+ $X2=0.695 $Y2=1.175
r86 30 32 46.6452 $w=3.72e-07 $l=3.6e-07 $layer=POLY_cond $X=0.6 $Y=1.202
+ $X2=0.96 $Y2=1.202
r87 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6 $Y=1.16
+ $X2=0.6 $Y2=1.16
r88 28 30 11.0134 $w=3.72e-07 $l=8.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.6 $Y2=1.202
r89 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r90 25 38 56.8409 $w=1.98e-07 $l=1.025e-06 $layer=LI1_cond $X=0.745 $Y=1.175
+ $X2=1.77 $Y2=1.175
r91 25 44 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.175
+ $X2=0.695 $Y2=1.175
r92 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r93 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r94 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r95 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r96 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r97 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r98 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r99 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r100 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r101 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r102 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r103 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=0.56
r104 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r105 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r106 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r107 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_4%A_459_21# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 38 41 45 49 50
c105 38 0 1.49142e-19 $X=4.38 $Y=1.16
c106 22 0 1.86355e-20 $X=3.335 $Y=1.41
c107 16 0 1.05834e-19 $X=2.865 $Y=1.41
c108 10 0 1.09002e-19 $X=2.395 $Y=1.41
r109 60 61 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.78 $Y=1.202
+ $X2=3.805 $Y2=1.202
r110 59 60 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=3.335 $Y=1.202
+ $X2=3.78 $Y2=1.202
r111 58 59 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.31 $Y=1.202
+ $X2=3.335 $Y2=1.202
r112 55 56 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.84 $Y=1.202
+ $X2=2.865 $Y2=1.202
r113 54 55 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.84 $Y2=1.202
r114 53 54 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.37 $Y=1.202
+ $X2=2.395 $Y2=1.202
r115 50 61 13.6879 $w=3.72e-07 $l=1.19164e-07 $layer=POLY_cond $X=3.905 $Y=1.16
+ $X2=3.805 $Y2=1.202
r116 45 47 21.7684 $w=3.58e-07 $l=6.8e-07 $layer=LI1_cond $X=4.575 $Y=1.66
+ $X2=4.575 $Y2=2.34
r117 43 49 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=1.245
+ $X2=4.575 $Y2=1.16
r118 43 45 13.2851 $w=3.58e-07 $l=4.15e-07 $layer=LI1_cond $X=4.575 $Y=1.245
+ $X2=4.575 $Y2=1.66
r119 39 49 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=1.075
+ $X2=4.575 $Y2=1.16
r120 39 41 21.9284 $w=3.58e-07 $l=6.85e-07 $layer=LI1_cond $X=4.575 $Y=1.075
+ $X2=4.575 $Y2=0.39
r121 38 50 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=4.38 $Y=1.16
+ $X2=3.905 $Y2=1.16
r122 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.38
+ $Y=1.16 $X2=4.38 $Y2=1.16
r123 34 58 6.47849 $w=3.72e-07 $l=5e-08 $layer=POLY_cond $X=3.26 $Y=1.202
+ $X2=3.31 $Y2=1.202
r124 34 56 51.1801 $w=3.72e-07 $l=3.95e-07 $layer=POLY_cond $X=3.26 $Y=1.202
+ $X2=2.865 $Y2=1.202
r125 33 37 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=3.26 $Y=1.16
+ $X2=4.38 $Y2=1.16
r126 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.26
+ $Y=1.16 $X2=3.26 $Y2=1.16
r127 31 49 4.14084 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=4.395 $Y=1.16
+ $X2=4.575 $Y2=1.16
r128 31 37 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.395 $Y=1.16
+ $X2=4.38 $Y2=1.16
r129 28 61 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.202
r130 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.985
r131 25 60 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.78 $Y=0.995
+ $X2=3.78 $Y2=1.202
r132 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.78 $Y=0.995
+ $X2=3.78 $Y2=0.56
r133 22 59 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.202
r134 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.985
r135 19 58 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=1.202
r136 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=0.56
r137 16 56 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.202
r138 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.985
r139 13 55 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=1.202
r140 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=0.56
r141 10 54 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.202
r142 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r143 7 53 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=1.202
r144 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=0.56
r145 2 47 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=1.485 $X2=4.59 $Y2=2.34
r146 2 45 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=1.485 $X2=4.59 $Y2=1.66
r147 1 41 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=4.445
+ $Y=0.235 $X2=4.59 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_4%B_N 1 3 4 6 7 10 17
c25 7 0 1.49142e-19 $X=5.2 $Y=1.105
r26 13 17 6.58539 $w=2.43e-07 $l=1.4e-07 $layer=LI1_cond $X=5.09 $Y=1.197
+ $X2=5.23 $Y2=1.197
r27 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.09
+ $Y=1.16 $X2=5.09 $Y2=1.16
r28 10 12 35.0907 $w=3.64e-07 $l=2.65e-07 $layer=POLY_cond $X=4.825 $Y=1.202
+ $X2=5.09 $Y2=1.202
r29 9 10 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=4.8 $Y=1.202
+ $X2=4.825 $Y2=1.202
r30 7 17 2.58712 $w=2.43e-07 $l=5.5e-08 $layer=LI1_cond $X=5.285 $Y=1.197
+ $X2=5.23 $Y2=1.197
r31 4 10 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.825 $Y=1.41
+ $X2=4.825 $Y2=1.202
r32 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.825 $Y=1.41
+ $X2=4.825 $Y2=1.985
r33 1 9 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.8 $Y=0.995 $X2=4.8
+ $Y2=1.202
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=0.995 $X2=4.8
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 28 29
+ 30 32 34 36 41 47
c88 28 0 7.78669e-20 $X=2.135 $Y=1.665
r89 47 49 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.075 $Y=2.02
+ $X2=3.075 $Y2=2.38
r90 34 52 2.49659 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.025 $Y=2.295
+ $X2=4.025 $Y2=2.38
r91 34 36 18.295 $w=3.98e-07 $l=6.35e-07 $layer=LI1_cond $X=4.025 $Y=2.295
+ $X2=4.025 $Y2=1.66
r92 33 49 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.265 $Y=2.38
+ $X2=3.075 $Y2=2.38
r93 32 52 5.87433 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.825 $Y=2.38 $X2=4.025
+ $Y2=2.38
r94 32 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.825 $Y=2.38
+ $X2=3.265 $Y2=2.38
r95 31 45 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.325 $Y=2.38
+ $X2=2.135 $Y2=2.38
r96 30 49 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.885 $Y=2.38
+ $X2=3.075 $Y2=2.38
r97 30 31 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.885 $Y=2.38
+ $X2=2.325 $Y2=2.38
r98 29 45 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=2.295
+ $X2=2.135 $Y2=2.38
r99 28 43 2.69784 $w=3.8e-07 $l=1.05e-07 $layer=LI1_cond $X=2.135 $Y=1.665
+ $X2=2.135 $Y2=1.56
r100 28 29 19.1063 $w=3.78e-07 $l=6.3e-07 $layer=LI1_cond $X=2.135 $Y=1.665
+ $X2=2.135 $Y2=2.295
r101 27 41 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=1.56
+ $X2=1.22 $Y2=1.56
r102 26 43 4.88181 $w=2.1e-07 $l=1.9e-07 $layer=LI1_cond $X=1.945 $Y=1.56
+ $X2=2.135 $Y2=1.56
r103 26 27 33.8009 $w=2.08e-07 $l=6.4e-07 $layer=LI1_cond $X=1.945 $Y=1.56
+ $X2=1.305 $Y2=1.56
r104 22 41 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.56
r105 22 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=2.3
r106 21 39 3.99943 $w=2.1e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=1.56
+ $X2=0.225 $Y2=1.56
r107 20 41 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=1.56
+ $X2=1.22 $Y2=1.56
r108 20 21 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=1.56
+ $X2=0.365 $Y2=1.56
r109 16 39 2.99957 $w=2.8e-07 $l=1.05e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=1.56
r110 16 18 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=2.3
r111 5 52 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.485 $X2=4.04 $Y2=2.34
r112 5 36 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.485 $X2=4.04 $Y2=1.66
r113 4 47 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=2.02
r114 3 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.34
r115 3 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.62
r116 2 41 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r117 2 24 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r118 1 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r119 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_4%VPWR 1 2 3 12 16 18 20 24 26 31 36 45 48
+ 52
r71 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r72 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r73 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r74 43 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r75 42 43 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r76 40 43 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=4.83 $Y2=2.72
r77 40 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r78 39 42 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=4.83 $Y2=2.72
r79 39 40 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r80 37 48 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.625 $Y2=2.72
r81 37 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=2.07 $Y2=2.72
r82 36 51 5.36004 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=4.975 $Y=2.72
+ $X2=5.247 $Y2=2.72
r83 36 42 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.975 $Y=2.72
+ $X2=4.83 $Y2=2.72
r84 35 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r85 35 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r87 32 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=0.725 $Y2=2.72
r88 32 34 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r89 31 48 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.625 $Y2=2.72
r90 31 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.15 $Y2=2.72
r91 26 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.725 $Y2=2.72
r92 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r93 24 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 20 23 19.3497 $w=4.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.177 $Y=1.66
+ $X2=5.177 $Y2=2.34
r96 18 51 3.05444 $w=4.05e-07 $l=1.14782e-07 $layer=LI1_cond $X=5.177 $Y=2.635
+ $X2=5.247 $Y2=2.72
r97 18 23 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=5.177 $Y=2.635
+ $X2=5.177 $Y2=2.34
r98 14 48 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.635
+ $X2=1.625 $Y2=2.72
r99 14 16 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=1.625 $Y=2.635
+ $X2=1.625 $Y2=2
r100 10 45 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=2.72
r101 10 12 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=2
r102 3 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.915
+ $Y=1.485 $X2=5.06 $Y2=2.34
r103 3 20 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.915
+ $Y=1.485 $X2=5.06 $Y2=1.66
r104 2 16 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=2
r105 1 12 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_4%Y 1 2 3 4 5 6 21 23 24 27 29 33 36 39 41
+ 45 47 49 51 52 55 56 59 63
c114 36 0 1.55605e-19 $X=2.71 $Y=1.415
r115 59 63 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.295 $Y=1.58
+ $X2=3.3 $Y2=1.58
r116 56 63 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.485 $Y=1.58
+ $X2=3.3 $Y2=1.58
r117 56 58 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=1.58
+ $X2=3.57 $Y2=1.58
r118 53 59 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.875 $Y=1.58
+ $X2=3.295 $Y2=1.58
r119 53 55 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=1.58
+ $X2=2.71 $Y2=1.58
r120 47 58 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.57 $Y=1.745
+ $X2=3.57 $Y2=1.58
r121 47 49 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.57 $Y=1.745
+ $X2=3.57 $Y2=1.96
r122 43 45 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.545 $Y2=0.39
r123 42 52 5.32988 $w=1.8e-07 $l=2.3e-07 $layer=LI1_cond $X=2.875 $Y=0.815
+ $X2=2.645 $Y2=0.815
r124 41 43 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=3.545 $Y2=0.725
r125 41 42 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=2.875 $Y2=0.815
r126 37 55 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=2.63 $Y=1.745
+ $X2=2.71 $Y2=1.58
r127 37 39 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.63 $Y=1.745
+ $X2=2.63 $Y2=1.96
r128 36 55 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=1.415
+ $X2=2.71 $Y2=1.58
r129 35 52 1.26734 $w=3.3e-07 $l=1.1811e-07 $layer=LI1_cond $X=2.71 $Y=0.905
+ $X2=2.645 $Y2=0.815
r130 35 36 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.71 $Y=0.905
+ $X2=2.71 $Y2=1.415
r131 31 52 1.26734 $w=3.8e-07 $l=1.08167e-07 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.645 $Y2=0.815
r132 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.605 $Y2=0.39
r133 30 51 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=0.815
+ $X2=1.665 $Y2=0.815
r134 29 52 5.32988 $w=1.8e-07 $l=2.3e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=2.645 $Y2=0.815
r135 29 30 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=1.855 $Y2=0.815
r136 25 51 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.815
r137 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.39
r138 23 51 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=1.665 $Y2=0.815
r139 23 24 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=0.915 $Y2=0.815
r140 19 24 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.815
r141 19 21 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r142 6 58 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=1.62
r143 6 49 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=1.96
r144 5 55 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=1.62
r145 5 39 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=1.96
r146 4 45 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.235 $X2=3.57 $Y2=0.39
r147 3 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.235 $X2=2.63 $Y2=0.39
r148 2 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r149 1 21 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2B_4%VGND 1 2 3 4 5 6 19 21 23 27 31 35 39 41
+ 43 46 47 49 50 52 53 54 66 74 78
r90 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r91 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r92 69 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r93 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r94 66 77 4.17994 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=4.975 $Y=0 $X2=5.247
+ $Y2=0
r95 66 68 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.975 $Y=0 $X2=4.83
+ $Y2=0
r96 65 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r97 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r98 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r99 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r100 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r101 59 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r102 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r103 56 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r104 56 58 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=2.07 $Y2=0
r105 54 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r106 54 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r107 52 64 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.955 $Y=0 $X2=3.91
+ $Y2=0
r108 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0 $X2=4.04
+ $Y2=0
r109 51 68 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.125 $Y=0
+ $X2=4.83 $Y2=0
r110 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0 $X2=4.04
+ $Y2=0
r111 49 61 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=2.99
+ $Y2=0
r112 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.1
+ $Y2=0
r113 48 64 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=3.91 $Y2=0
r114 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.1
+ $Y2=0
r115 46 58 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r116 46 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.16
+ $Y2=0
r117 45 61 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.99 $Y2=0
r118 45 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r119 41 77 3.2579 $w=2.9e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.12 $Y=0.085
+ $X2=5.247 $Y2=0
r120 41 43 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=5.12 $Y=0.085
+ $X2=5.12 $Y2=0.39
r121 37 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r122 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.39
r123 33 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0
r124 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0.39
r125 29 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r126 29 31 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.39
r127 25 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r128 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r129 24 71 4.33083 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r130 23 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r131 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=0.365 $Y2=0
r132 19 71 3.02922 $w=2.8e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.182 $Y2=0
r133 19 21 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.39
r134 6 43 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.875
+ $Y=0.235 $X2=5.06 $Y2=0.39
r135 5 39 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.855
+ $Y=0.235 $X2=4.04 $Y2=0.39
r136 4 35 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.39
r137 3 31 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r138 2 27 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
r139 1 21 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

