* File: sky130_fd_sc_hdll__xor2_4.pex.spice
* Created: Wed Sep  2 08:54:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XOR2_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 50 51 52 53 54 57 60 64 78 88
c228 52 0 1.27704e-19 $X=3.1 $Y=1.53
c229 50 0 1.71198e-19 $X=2.99 $Y=1.445
r230 88 89 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.08 $Y=1.202
+ $X2=8.105 $Y2=1.202
r231 85 86 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.585 $Y=1.202
+ $X2=7.61 $Y2=1.202
r232 84 85 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=7.14 $Y=1.202
+ $X2=7.585 $Y2=1.202
r233 83 84 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.115 $Y=1.202
+ $X2=7.14 $Y2=1.202
r234 80 81 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.645 $Y=1.202
+ $X2=6.67 $Y2=1.202
r235 78 79 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.92 $Y=1.202
+ $X2=1.945 $Y2=1.202
r236 76 78 20.0833 $w=3.72e-07 $l=1.55e-07 $layer=POLY_cond $X=1.765 $Y=1.202
+ $X2=1.92 $Y2=1.202
r237 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.765
+ $Y=1.16 $X2=1.765 $Y2=1.16
r238 74 76 40.8145 $w=3.72e-07 $l=3.15e-07 $layer=POLY_cond $X=1.45 $Y=1.202
+ $X2=1.765 $Y2=1.202
r239 73 74 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.425 $Y=1.202
+ $X2=1.45 $Y2=1.202
r240 72 73 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.98 $Y=1.202
+ $X2=1.425 $Y2=1.202
r241 71 72 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.955 $Y=1.202
+ $X2=0.98 $Y2=1.202
r242 69 71 46.6452 $w=3.72e-07 $l=3.6e-07 $layer=POLY_cond $X=0.595 $Y=1.202
+ $X2=0.955 $Y2=1.202
r243 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r244 67 69 11.0134 $w=3.72e-07 $l=8.5e-08 $layer=POLY_cond $X=0.51 $Y=1.202
+ $X2=0.595 $Y2=1.202
r245 66 67 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.485 $Y=1.202
+ $X2=0.51 $Y2=1.202
r246 64 77 34.1045 $w=1.98e-07 $l=6.15e-07 $layer=LI1_cond $X=1.15 $Y=1.175
+ $X2=1.765 $Y2=1.175
r247 64 70 30.7773 $w=1.98e-07 $l=5.55e-07 $layer=LI1_cond $X=1.15 $Y=1.175
+ $X2=0.595 $Y2=1.175
r248 63 83 44.7016 $w=3.72e-07 $l=3.45e-07 $layer=POLY_cond $X=6.77 $Y=1.202
+ $X2=7.115 $Y2=1.202
r249 63 81 12.957 $w=3.72e-07 $l=1e-07 $layer=POLY_cond $X=6.77 $Y=1.202
+ $X2=6.67 $Y2=1.202
r250 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.77
+ $Y=1.16 $X2=6.77 $Y2=1.16
r251 60 77 61.8318 $w=1.98e-07 $l=1.115e-06 $layer=LI1_cond $X=2.88 $Y=1.175
+ $X2=1.765 $Y2=1.175
r252 58 88 18.1398 $w=3.72e-07 $l=1.4e-07 $layer=POLY_cond $X=7.94 $Y=1.202
+ $X2=8.08 $Y2=1.202
r253 58 86 42.7581 $w=3.72e-07 $l=3.3e-07 $layer=POLY_cond $X=7.94 $Y=1.202
+ $X2=7.61 $Y2=1.202
r254 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.94
+ $Y=1.16 $X2=7.94 $Y2=1.16
r255 55 62 3.58108 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=6.815 $Y=1.175
+ $X2=6.705 $Y2=1.175
r256 55 57 62.3864 $w=1.98e-07 $l=1.125e-06 $layer=LI1_cond $X=6.815 $Y=1.175
+ $X2=7.94 $Y2=1.175
r257 53 62 3.25553 $w=2.2e-07 $l=1e-07 $layer=LI1_cond $X=6.705 $Y=1.275
+ $X2=6.705 $Y2=1.175
r258 53 54 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=6.705 $Y=1.275
+ $X2=6.705 $Y2=1.445
r259 51 54 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.595 $Y=1.53
+ $X2=6.705 $Y2=1.445
r260 51 52 228.016 $w=1.68e-07 $l=3.495e-06 $layer=LI1_cond $X=6.595 $Y=1.53
+ $X2=3.1 $Y2=1.53
r261 50 52 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.99 $Y=1.445
+ $X2=3.1 $Y2=1.53
r262 49 60 6.83662 $w=2e-07 $l=1.51987e-07 $layer=LI1_cond $X=2.99 $Y=1.275
+ $X2=2.88 $Y2=1.175
r263 49 50 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=2.99 $Y=1.275
+ $X2=2.99 $Y2=1.445
r264 46 89 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.105 $Y=0.995
+ $X2=8.105 $Y2=1.202
r265 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.105 $Y=0.995
+ $X2=8.105 $Y2=0.56
r266 43 88 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.08 $Y=1.41
+ $X2=8.08 $Y2=1.202
r267 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.08 $Y=1.41
+ $X2=8.08 $Y2=1.985
r268 40 86 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.61 $Y=1.41
+ $X2=7.61 $Y2=1.202
r269 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.61 $Y=1.41
+ $X2=7.61 $Y2=1.985
r270 37 85 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.585 $Y=0.995
+ $X2=7.585 $Y2=1.202
r271 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.585 $Y=0.995
+ $X2=7.585 $Y2=0.56
r272 34 84 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.14 $Y=1.41
+ $X2=7.14 $Y2=1.202
r273 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.14 $Y=1.41
+ $X2=7.14 $Y2=1.985
r274 31 83 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.115 $Y=0.995
+ $X2=7.115 $Y2=1.202
r275 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.115 $Y=0.995
+ $X2=7.115 $Y2=0.56
r276 28 81 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.67 $Y=1.41
+ $X2=6.67 $Y2=1.202
r277 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.67 $Y=1.41
+ $X2=6.67 $Y2=1.985
r278 25 80 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.645 $Y=0.995
+ $X2=6.645 $Y2=1.202
r279 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.645 $Y=0.995
+ $X2=6.645 $Y2=0.56
r280 22 79 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.945 $Y=0.995
+ $X2=1.945 $Y2=1.202
r281 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.945 $Y=0.995
+ $X2=1.945 $Y2=0.56
r282 19 78 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.92 $Y=1.41
+ $X2=1.92 $Y2=1.202
r283 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.92 $Y=1.41
+ $X2=1.92 $Y2=1.985
r284 16 74 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.45 $Y=1.41
+ $X2=1.45 $Y2=1.202
r285 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.45 $Y=1.41
+ $X2=1.45 $Y2=1.985
r286 13 73 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.425 $Y=0.995
+ $X2=1.425 $Y2=1.202
r287 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.425 $Y=0.995
+ $X2=1.425 $Y2=0.56
r288 10 72 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.202
r289 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.985
r290 7 71 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=1.202
r291 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r292 4 67 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.202
r293 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.985
r294 1 66 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.202
r295 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 27 29 30 32 33 35 36 38 39 41 42 44 45 47 48 50 55 74 77 83
c152 33 0 1.11496e-19 $X=5.235 $Y=0.995
c153 10 0 1.51917e-19 $X=2.86 $Y=1.41
c154 4 0 1.71198e-19 $X=2.39 $Y=1.41
r155 77 78 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.2 $Y=1.202
+ $X2=6.225 $Y2=1.202
r156 76 77 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=5.73 $Y=1.202
+ $X2=6.2 $Y2=1.202
r157 75 76 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.705 $Y=1.202
+ $X2=5.73 $Y2=1.202
r158 74 83 51.5727 $w=1.98e-07 $l=9.3e-07 $layer=LI1_cond $X=5.285 $Y=1.175
+ $X2=4.355 $Y2=1.175
r159 73 75 54.4194 $w=3.72e-07 $l=4.2e-07 $layer=POLY_cond $X=5.285 $Y=1.202
+ $X2=5.705 $Y2=1.202
r160 73 74 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=5.285
+ $Y=1.16 $X2=5.285 $Y2=1.16
r161 71 73 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.26 $Y=1.202
+ $X2=5.285 $Y2=1.202
r162 70 71 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.235 $Y=1.202
+ $X2=5.26 $Y2=1.202
r163 69 70 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.79 $Y=1.202
+ $X2=5.235 $Y2=1.202
r164 68 69 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.765 $Y=1.202
+ $X2=4.79 $Y2=1.202
r165 66 67 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.775 $Y=1.202
+ $X2=3.8 $Y2=1.202
r166 64 66 44.0538 $w=3.72e-07 $l=3.4e-07 $layer=POLY_cond $X=3.435 $Y=1.202
+ $X2=3.775 $Y2=1.202
r167 64 65 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.435
+ $Y=1.16 $X2=3.435 $Y2=1.16
r168 62 64 13.6048 $w=3.72e-07 $l=1.05e-07 $layer=POLY_cond $X=3.33 $Y=1.202
+ $X2=3.435 $Y2=1.202
r169 61 62 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.305 $Y=1.202
+ $X2=3.33 $Y2=1.202
r170 60 61 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.86 $Y=1.202
+ $X2=3.305 $Y2=1.202
r171 59 60 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.835 $Y=1.202
+ $X2=2.86 $Y2=1.202
r172 58 59 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.39 $Y=1.202
+ $X2=2.835 $Y2=1.202
r173 57 58 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.365 $Y=1.202
+ $X2=2.39 $Y2=1.202
r174 55 83 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=4.35 $Y=1.175
+ $X2=4.355 $Y2=1.175
r175 55 65 50.7409 $w=1.98e-07 $l=9.15e-07 $layer=LI1_cond $X=4.35 $Y=1.175
+ $X2=3.435 $Y2=1.175
r176 48 78 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.225 $Y=0.995
+ $X2=6.225 $Y2=1.202
r177 48 50 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.225 $Y=0.995
+ $X2=6.225 $Y2=0.56
r178 45 77 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.2 $Y=1.41
+ $X2=6.2 $Y2=1.202
r179 45 47 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.2 $Y=1.41
+ $X2=6.2 $Y2=1.985
r180 42 76 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.73 $Y2=1.202
r181 42 44 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.73 $Y2=1.985
r182 39 75 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.705 $Y=0.995
+ $X2=5.705 $Y2=1.202
r183 39 41 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.705 $Y=0.995
+ $X2=5.705 $Y2=0.56
r184 36 71 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.26 $Y=1.41
+ $X2=5.26 $Y2=1.202
r185 36 38 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.26 $Y=1.41
+ $X2=5.26 $Y2=1.985
r186 33 70 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.235 $Y2=1.202
r187 33 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.235 $Y2=0.56
r188 30 69 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.79 $Y=1.41
+ $X2=4.79 $Y2=1.202
r189 30 32 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.79 $Y=1.41
+ $X2=4.79 $Y2=1.985
r190 27 68 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.765 $Y=0.995
+ $X2=4.765 $Y2=1.202
r191 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.765 $Y=0.995
+ $X2=4.765 $Y2=0.56
r192 26 67 13.6879 $w=3.72e-07 $l=1.19164e-07 $layer=POLY_cond $X=3.9 $Y=1.16
+ $X2=3.8 $Y2=1.202
r193 25 68 10.4487 $w=3.72e-07 $l=9.3675e-08 $layer=POLY_cond $X=4.69 $Y=1.16
+ $X2=4.765 $Y2=1.202
r194 25 26 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=4.69 $Y=1.16 $X2=3.9
+ $Y2=1.16
r195 22 67 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.8 $Y=1.41
+ $X2=3.8 $Y2=1.202
r196 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.8 $Y=1.41
+ $X2=3.8 $Y2=1.985
r197 19 66 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.775 $Y=0.995
+ $X2=3.775 $Y2=1.202
r198 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.775 $Y=0.995
+ $X2=3.775 $Y2=0.56
r199 16 62 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.33 $Y=1.41
+ $X2=3.33 $Y2=1.202
r200 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.33 $Y=1.41
+ $X2=3.33 $Y2=1.985
r201 13 61 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.305 $Y=0.995
+ $X2=3.305 $Y2=1.202
r202 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.305 $Y=0.995
+ $X2=3.305 $Y2=0.56
r203 10 60 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.86 $Y=1.41
+ $X2=2.86 $Y2=1.202
r204 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.86 $Y=1.41
+ $X2=2.86 $Y2=1.985
r205 7 59 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.835 $Y=0.995
+ $X2=2.835 $Y2=1.202
r206 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.835 $Y=0.995
+ $X2=2.835 $Y2=0.56
r207 4 58 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.39 $Y=1.41
+ $X2=2.39 $Y2=1.202
r208 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.39 $Y=1.41
+ $X2=2.39 $Y2=1.985
r209 1 57 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.365 $Y=0.995
+ $X2=2.365 $Y2=1.202
r210 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.365 $Y=0.995
+ $X2=2.365 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_4%A_112_47# 1 2 3 4 5 6 19 21 22 24 25 27 28
+ 30 31 33 34 36 37 39 40 42 44 45 46 49 51 55 57 61 65 67 71 76 77 82 85 86 87
+ 88 89 90 91 95 100 101 107 108 118
c279 101 0 2.79621e-19 $X=2.415 $Y=1.53
c280 31 0 3.03462e-20 $X=9.995 $Y=0.995
c281 25 0 9.87024e-20 $X=9.525 $Y=0.995
r282 118 119 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=10.49 $Y=1.202
+ $X2=10.515 $Y2=1.202
r283 117 118 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=10.02 $Y=1.202
+ $X2=10.49 $Y2=1.202
r284 116 117 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.995 $Y=1.202
+ $X2=10.02 $Y2=1.202
r285 113 114 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.525 $Y=1.202
+ $X2=9.55 $Y2=1.202
r286 110 111 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.055 $Y=1.202
+ $X2=9.08 $Y2=1.202
r287 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.39 $Y=1.53
+ $X2=8.39 $Y2=1.53
r288 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.27 $Y=1.53
+ $X2=2.27 $Y2=1.53
r289 101 103 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.415 $Y=1.53
+ $X2=2.27 $Y2=1.53
r290 100 107 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.245 $Y=1.53
+ $X2=8.39 $Y2=1.53
r291 100 101 7.21533 $w=1.4e-07 $l=5.83e-06 $layer=MET1_cond $X=8.245 $Y=1.53
+ $X2=2.415 $Y2=1.53
r292 95 98 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.565 $Y=1.87
+ $X2=3.565 $Y2=1.96
r293 90 93 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.625 $Y=1.87
+ $X2=2.625 $Y2=1.96
r294 90 91 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=1.87
+ $X2=2.625 $Y2=1.785
r295 89 104 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.5 $Y=1.53
+ $X2=2.27 $Y2=1.53
r296 85 104 131.46 $w=1.68e-07 $l=2.015e-06 $layer=LI1_cond $X=0.255 $Y=1.53
+ $X2=2.27 $Y2=1.53
r297 83 116 6.47849 $w=3.72e-07 $l=5e-08 $layer=POLY_cond $X=9.945 $Y=1.202
+ $X2=9.995 $Y2=1.202
r298 83 114 51.1801 $w=3.72e-07 $l=3.95e-07 $layer=POLY_cond $X=9.945 $Y=1.202
+ $X2=9.55 $Y2=1.202
r299 82 83 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.945
+ $Y=1.16 $X2=9.945 $Y2=1.16
r300 80 113 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=9.145 $Y=1.202
+ $X2=9.525 $Y2=1.202
r301 80 111 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=9.145 $Y=1.202
+ $X2=9.08 $Y2=1.202
r302 79 82 44.3636 $w=1.98e-07 $l=8e-07 $layer=LI1_cond $X=9.145 $Y=1.175
+ $X2=9.945 $Y2=1.175
r303 79 80 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.145
+ $Y=1.16 $X2=9.145 $Y2=1.16
r304 77 79 35.2136 $w=1.98e-07 $l=6.35e-07 $layer=LI1_cond $X=8.51 $Y=1.175
+ $X2=9.145 $Y2=1.175
r305 76 108 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.425 $Y=1.445
+ $X2=8.425 $Y2=1.53
r306 75 77 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=8.425 $Y=1.275
+ $X2=8.51 $Y2=1.175
r307 75 76 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.425 $Y=1.275
+ $X2=8.425 $Y2=1.445
r308 69 71 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.54 $Y=0.725
+ $X2=3.54 $Y2=0.39
r309 68 88 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.79 $Y=0.815
+ $X2=2.6 $Y2=0.815
r310 67 69 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=3.35 $Y=0.815
+ $X2=3.54 $Y2=0.725
r311 67 68 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.35 $Y=0.815
+ $X2=2.79 $Y2=0.815
r312 66 90 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.75 $Y=1.87
+ $X2=2.625 $Y2=1.87
r313 65 95 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.44 $Y=1.87
+ $X2=3.565 $Y2=1.87
r314 65 66 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.44 $Y=1.87
+ $X2=2.75 $Y2=1.87
r315 63 89 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.585 $Y=1.615
+ $X2=2.5 $Y2=1.53
r316 63 91 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.585 $Y=1.615
+ $X2=2.585 $Y2=1.785
r317 59 88 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=2.6 $Y=0.725 $X2=2.6
+ $Y2=0.815
r318 59 61 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.6 $Y=0.725
+ $X2=2.6 $Y2=0.39
r319 58 87 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.85 $Y=0.815
+ $X2=1.66 $Y2=0.815
r320 57 88 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.41 $Y=0.815
+ $X2=2.6 $Y2=0.815
r321 57 58 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.41 $Y=0.815
+ $X2=1.85 $Y2=0.815
r322 53 87 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.66 $Y=0.725 $X2=1.66
+ $Y2=0.815
r323 53 55 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.66 $Y=0.725
+ $X2=1.66 $Y2=0.39
r324 52 86 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=0.815
+ $X2=0.72 $Y2=0.815
r325 51 87 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.47 $Y=0.815
+ $X2=1.66 $Y2=0.815
r326 51 52 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.47 $Y=0.815
+ $X2=0.91 $Y2=0.815
r327 47 86 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=0.725 $X2=0.72
+ $Y2=0.815
r328 47 49 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=0.725
+ $X2=0.72 $Y2=0.39
r329 45 86 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=0.53 $Y=0.82
+ $X2=0.72 $Y2=0.815
r330 45 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.53 $Y=0.82
+ $X2=0.255 $Y2=0.82
r331 44 85 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.445
+ $X2=0.255 $Y2=1.53
r332 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=0.905
+ $X2=0.255 $Y2=0.82
r333 43 44 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.17 $Y=0.905
+ $X2=0.17 $Y2=1.445
r334 40 119 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.515 $Y=0.995
+ $X2=10.515 $Y2=1.202
r335 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.515 $Y=0.995
+ $X2=10.515 $Y2=0.56
r336 37 118 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.49 $Y=1.41
+ $X2=10.49 $Y2=1.202
r337 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.49 $Y=1.41
+ $X2=10.49 $Y2=1.985
r338 34 117 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.02 $Y=1.41
+ $X2=10.02 $Y2=1.202
r339 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.02 $Y=1.41
+ $X2=10.02 $Y2=1.985
r340 31 116 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.995 $Y=0.995
+ $X2=9.995 $Y2=1.202
r341 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.995 $Y=0.995
+ $X2=9.995 $Y2=0.56
r342 28 114 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.55 $Y=1.41
+ $X2=9.55 $Y2=1.202
r343 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.55 $Y=1.41
+ $X2=9.55 $Y2=1.985
r344 25 113 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.525 $Y=0.995
+ $X2=9.525 $Y2=1.202
r345 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.525 $Y=0.995
+ $X2=9.525 $Y2=0.56
r346 22 111 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.08 $Y=1.41
+ $X2=9.08 $Y2=1.202
r347 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.08 $Y=1.41
+ $X2=9.08 $Y2=1.985
r348 19 110 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.055 $Y=0.995
+ $X2=9.055 $Y2=1.202
r349 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.055 $Y=0.995
+ $X2=9.055 $Y2=0.56
r350 6 98 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.485 $X2=3.565 $Y2=1.96
r351 5 93 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.485 $X2=2.625 $Y2=1.96
r352 4 71 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.38
+ $Y=0.235 $X2=3.565 $Y2=0.39
r353 3 61 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.44
+ $Y=0.235 $X2=2.625 $Y2=0.39
r354 2 55 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.235 $X2=1.685 $Y2=0.39
r355 1 49 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.235 $X2=0.745 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_4%A_27_297# 1 2 3 4 5 18 22 24 26 27 28 32 35
+ 37 41
r64 41 43 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.095 $Y=2.3 $X2=3.095
+ $Y2=2.38
r65 30 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.035 $Y=2.295
+ $X2=4.035 $Y2=1.96
r66 29 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.22 $Y=2.38
+ $X2=3.095 $Y2=2.38
r67 28 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.91 $Y=2.38
+ $X2=4.035 $Y2=2.295
r68 28 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.91 $Y=2.38 $X2=3.22
+ $Y2=2.38
r69 26 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.97 $Y=2.38
+ $X2=3.095 $Y2=2.38
r70 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.97 $Y=2.38 $X2=2.28
+ $Y2=2.38
r71 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.155 $Y=2.295
+ $X2=2.28 $Y2=2.38
r72 24 39 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=2.155 $Y=2.005
+ $X2=2.155 $Y2=1.895
r73 24 25 13.3683 $w=2.48e-07 $l=2.9e-07 $layer=LI1_cond $X=2.155 $Y=2.005
+ $X2=2.155 $Y2=2.295
r74 23 37 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.34 $Y=1.895
+ $X2=1.215 $Y2=1.895
r75 22 39 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.03 $Y=1.895
+ $X2=2.155 $Y2=1.895
r76 22 23 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=2.03 $Y=1.895
+ $X2=1.34 $Y2=1.895
r77 19 35 4.18571 $w=2.2e-07 $l=1.58e-07 $layer=LI1_cond $X=0.4 $Y=1.895
+ $X2=0.242 $Y2=1.895
r78 18 37 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.09 $Y=1.895
+ $X2=1.215 $Y2=1.895
r79 18 19 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=1.09 $Y=1.895
+ $X2=0.4 $Y2=1.895
r80 5 32 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.89
+ $Y=1.485 $X2=4.035 $Y2=1.96
r81 4 41 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.95
+ $Y=1.485 $X2=3.095 $Y2=2.3
r82 3 39 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.01
+ $Y=1.485 $X2=2.155 $Y2=1.96
r83 2 37 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.485 $X2=1.215 $Y2=1.96
r84 1 35 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_4%VPWR 1 2 3 4 5 6 23 25 29 33 37 41 45 48 49
+ 51 52 54 55 57 58 59 81 82 85 88
r156 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r157 86 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r158 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r159 81 82 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r160 79 82 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=10.81 $Y2=2.72
r161 78 81 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=10.81 $Y2=2.72
r162 78 79 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r163 76 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r164 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r165 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r166 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r167 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r168 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r169 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r170 66 67 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r171 64 67 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=4.83 $Y2=2.72
r172 64 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r173 63 66 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=4.83 $Y2=2.72
r174 63 64 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r175 61 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=2.72
+ $X2=1.685 $Y2=2.72
r176 61 63 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.81 $Y=2.72
+ $X2=2.07 $Y2=2.72
r177 59 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r178 57 75 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.72 $Y=2.72
+ $X2=7.59 $Y2=2.72
r179 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.72 $Y=2.72
+ $X2=7.845 $Y2=2.72
r180 56 78 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.97 $Y=2.72 $X2=8.05
+ $Y2=2.72
r181 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.97 $Y=2.72
+ $X2=7.845 $Y2=2.72
r182 54 72 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.78 $Y=2.72
+ $X2=6.67 $Y2=2.72
r183 54 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.78 $Y=2.72
+ $X2=6.905 $Y2=2.72
r184 53 75 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.03 $Y=2.72
+ $X2=7.59 $Y2=2.72
r185 53 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.03 $Y=2.72
+ $X2=6.905 $Y2=2.72
r186 51 69 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.84 $Y=2.72 $X2=5.75
+ $Y2=2.72
r187 51 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.84 $Y=2.72
+ $X2=5.965 $Y2=2.72
r188 50 72 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.09 $Y=2.72
+ $X2=6.67 $Y2=2.72
r189 50 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.09 $Y=2.72
+ $X2=5.965 $Y2=2.72
r190 48 66 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.9 $Y=2.72 $X2=4.83
+ $Y2=2.72
r191 48 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.9 $Y=2.72
+ $X2=5.025 $Y2=2.72
r192 47 69 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.15 $Y=2.72 $X2=5.75
+ $Y2=2.72
r193 47 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.15 $Y=2.72
+ $X2=5.025 $Y2=2.72
r194 43 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=2.635
+ $X2=7.845 $Y2=2.72
r195 43 45 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.845 $Y=2.635
+ $X2=7.845 $Y2=2.34
r196 39 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=2.635
+ $X2=6.905 $Y2=2.72
r197 39 41 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=6.905 $Y=2.635
+ $X2=6.905 $Y2=2.34
r198 35 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=2.635
+ $X2=5.965 $Y2=2.72
r199 35 37 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.965 $Y=2.635
+ $X2=5.965 $Y2=2.34
r200 31 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=2.635
+ $X2=5.025 $Y2=2.72
r201 31 33 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.025 $Y=2.635
+ $X2=5.025 $Y2=2.34
r202 27 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=2.635
+ $X2=1.685 $Y2=2.72
r203 27 29 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.685 $Y=2.635
+ $X2=1.685 $Y2=2.34
r204 26 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=0.745 $Y2=2.72
r205 25 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.56 $Y=2.72
+ $X2=1.685 $Y2=2.72
r206 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.56 $Y=2.72
+ $X2=0.87 $Y2=2.72
r207 21 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.72
r208 21 23 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.34
r209 6 45 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.7
+ $Y=1.485 $X2=7.845 $Y2=2.34
r210 5 41 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.76
+ $Y=1.485 $X2=6.905 $Y2=2.34
r211 4 37 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.485 $X2=5.965 $Y2=2.34
r212 3 33 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.485 $X2=5.025 $Y2=2.34
r213 2 29 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.485 $X2=1.685 $Y2=2.34
r214 1 23 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.485 $X2=0.745 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_4%A_886_297# 1 2 3 4 5 6 7 24 28 32 36 40 42
+ 43 44 45 48 50 54 57 59 61 63 66
r110 52 54 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=10.255 $Y=2.295
+ $X2=10.255 $Y2=1.96
r111 51 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.44 $Y=2.38
+ $X2=9.315 $Y2=2.38
r112 50 52 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.13 $Y=2.38
+ $X2=10.255 $Y2=2.295
r113 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.13 $Y=2.38
+ $X2=9.44 $Y2=2.38
r114 46 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.315 $Y=2.295
+ $X2=9.315 $Y2=2.38
r115 46 48 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=9.315 $Y=2.295
+ $X2=9.315 $Y2=2
r116 44 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.19 $Y=2.38
+ $X2=9.315 $Y2=2.38
r117 44 45 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=9.19 $Y=2.38
+ $X2=8.44 $Y2=2.38
r118 43 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.315 $Y=2.295
+ $X2=8.44 $Y2=2.38
r119 42 65 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=8.315 $Y=2.005
+ $X2=8.315 $Y2=1.895
r120 42 43 13.3683 $w=2.48e-07 $l=2.9e-07 $layer=LI1_cond $X=8.315 $Y=2.005
+ $X2=8.315 $Y2=2.295
r121 41 63 6.93182 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=7.5 $Y=1.895
+ $X2=7.375 $Y2=1.895
r122 40 65 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=8.19 $Y=1.895
+ $X2=8.315 $Y2=1.895
r123 40 41 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=8.19 $Y=1.895
+ $X2=7.5 $Y2=1.895
r124 34 63 5.368 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=7.375 $Y=1.785
+ $X2=7.375 $Y2=1.895
r125 34 36 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=1.785
+ $X2=7.375 $Y2=1.62
r126 33 61 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=6.56 $Y=1.895
+ $X2=6.435 $Y2=1.895
r127 32 63 6.93182 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=7.25 $Y=1.895
+ $X2=7.375 $Y2=1.895
r128 32 33 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=7.25 $Y=1.895
+ $X2=6.56 $Y2=1.895
r129 29 59 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.62 $Y=1.895
+ $X2=5.495 $Y2=1.895
r130 28 61 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=6.31 $Y=1.895
+ $X2=6.435 $Y2=1.895
r131 28 29 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=6.31 $Y=1.895
+ $X2=5.62 $Y2=1.895
r132 25 57 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=4.68 $Y=1.895
+ $X2=4.555 $Y2=1.895
r133 24 59 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.37 $Y=1.895
+ $X2=5.495 $Y2=1.895
r134 24 25 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=5.37 $Y=1.895
+ $X2=4.68 $Y2=1.895
r135 7 54 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.11
+ $Y=1.485 $X2=10.255 $Y2=1.96
r136 6 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.17
+ $Y=1.485 $X2=9.315 $Y2=2
r137 5 65 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.17
+ $Y=1.485 $X2=8.315 $Y2=1.96
r138 4 63 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.23
+ $Y=1.485 $X2=7.375 $Y2=1.96
r139 4 36 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.485 $X2=7.375 $Y2=1.62
r140 3 61 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.29
+ $Y=1.485 $X2=6.435 $Y2=1.96
r141 2 59 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.35
+ $Y=1.485 $X2=5.495 $Y2=1.96
r142 1 57 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.485 $X2=4.555 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_4%X 1 2 3 4 5 6 7 26 28 30 34 36 40 44 46 49
+ 52 53 55 56 59 60 68 70 72 77 79
c159 70 0 9.87024e-20 $X=8.85 $Y=0.81
c160 68 0 1.11496e-19 $X=5.935 $Y=0.81
c161 53 0 3.03462e-20 $X=9.29 $Y=0.815
r162 70 72 0.113092 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.85 $Y=0.81
+ $X2=8.705 $Y2=0.81
r163 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.85 $Y=0.81
+ $X2=8.85 $Y2=0.81
r164 68 72 3.22694 $w=1.45e-07 $l=2.77e-06 $layer=MET1_cond $X=5.935 $Y=0.852
+ $X2=8.705 $Y2=0.852
r165 66 79 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=5.79 $Y=0.79
+ $X2=5.965 $Y2=0.79
r166 66 77 5.71274 $w=2.88e-07 $l=1.4e-07 $layer=LI1_cond $X=5.79 $Y=0.79
+ $X2=5.65 $Y2=0.79
r167 65 68 0.113092 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.79 $Y=0.81
+ $X2=5.935 $Y2=0.81
r168 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.79 $Y=0.81
+ $X2=5.79 $Y2=0.81
r169 60 84 12.2358 $w=4.03e-07 $l=4.3e-07 $layer=LI1_cond $X=10.752 $Y=1.87
+ $X2=10.752 $Y2=2.3
r170 57 60 6.97157 $w=4.03e-07 $l=2.45e-07 $layer=LI1_cond $X=10.752 $Y=1.625
+ $X2=10.752 $Y2=1.87
r171 57 59 2.79199 $w=3.62e-07 $l=9e-08 $layer=LI1_cond $X=10.752 $Y=1.625
+ $X2=10.752 $Y2=1.535
r172 52 71 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=9.1 $Y=0.815
+ $X2=8.85 $Y2=0.815
r173 52 53 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=9.1 $Y=0.815
+ $X2=9.29 $Y2=0.815
r174 49 59 2.79199 $w=3.62e-07 $l=1.09407e-07 $layer=LI1_cond $X=10.795 $Y=1.445
+ $X2=10.752 $Y2=1.535
r175 48 49 19.4475 $w=3.18e-07 $l=5.4e-07 $layer=LI1_cond $X=10.795 $Y=0.905
+ $X2=10.795 $Y2=1.445
r176 47 56 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.42 $Y=0.82
+ $X2=10.23 $Y2=0.82
r177 46 48 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=10.635 $Y=0.82
+ $X2=10.795 $Y2=0.905
r178 46 47 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.635 $Y=0.82
+ $X2=10.42 $Y2=0.82
r179 42 56 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.23 $Y=0.735
+ $X2=10.23 $Y2=0.82
r180 42 44 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=10.23 $Y=0.735
+ $X2=10.23 $Y2=0.39
r181 41 55 6.19399 $w=2e-07 $l=1.34629e-07 $layer=LI1_cond $X=9.91 $Y=1.535
+ $X2=9.785 $Y2=1.555
r182 40 59 3.94943 $w=1.8e-07 $l=2.02e-07 $layer=LI1_cond $X=10.55 $Y=1.535
+ $X2=10.752 $Y2=1.535
r183 40 41 39.4343 $w=1.78e-07 $l=6.4e-07 $layer=LI1_cond $X=10.55 $Y=1.535
+ $X2=9.91 $Y2=1.535
r184 37 53 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=9.48 $Y=0.82
+ $X2=9.29 $Y2=0.815
r185 36 56 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.04 $Y=0.82
+ $X2=10.23 $Y2=0.82
r186 36 37 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=10.04 $Y=0.82
+ $X2=9.48 $Y2=0.82
r187 32 53 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=9.29 $Y=0.725 $X2=9.29
+ $Y2=0.815
r188 32 34 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.29 $Y=0.725
+ $X2=9.29 $Y2=0.39
r189 31 51 3.97178 $w=2.2e-07 $l=1.45e-07 $layer=LI1_cond $X=8.97 $Y=1.555
+ $X2=8.825 $Y2=1.555
r190 30 55 6.19399 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=9.66 $Y=1.555
+ $X2=9.785 $Y2=1.555
r191 30 31 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=9.66 $Y=1.555
+ $X2=8.97 $Y2=1.555
r192 26 51 3.01307 $w=2.9e-07 $l=1.1e-07 $layer=LI1_cond $X=8.825 $Y=1.665
+ $X2=8.825 $Y2=1.555
r193 26 28 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=8.825 $Y=1.665
+ $X2=8.825 $Y2=1.96
r194 24 77 27.703 $w=2.58e-07 $l=6.25e-07 $layer=LI1_cond $X=5.025 $Y=0.775
+ $X2=5.65 $Y2=0.775
r195 7 84 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=10.58
+ $Y=1.485 $X2=10.725 $Y2=2.3
r196 7 59 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.58
+ $Y=1.485 $X2=10.725 $Y2=1.62
r197 6 55 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.64
+ $Y=1.485 $X2=9.785 $Y2=1.62
r198 5 51 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.485 $X2=8.845 $Y2=1.61
r199 5 28 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.485 $X2=8.845 $Y2=1.96
r200 4 44 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=10.07
+ $Y=0.235 $X2=10.255 $Y2=0.39
r201 3 34 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=9.13
+ $Y=0.235 $X2=9.315 $Y2=0.39
r202 2 79 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=5.78
+ $Y=0.235 $X2=5.965 $Y2=0.73
r203 1 24 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.235 $X2=5.025 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_4%VGND 1 2 3 4 5 6 7 8 9 10 31 33 35 39 41 45
+ 49 53 57 61 65 69 71 73 76 77 79 80 82 83 85 86 88 89 91 92 93 117 125 128 132
r191 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r192 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r193 126 129 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r194 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r195 120 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r196 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r197 117 131 3.40825 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.64 $Y=0 $X2=10.84
+ $Y2=0
r198 117 119 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.64 $Y=0
+ $X2=10.35 $Y2=0
r199 116 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r200 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r201 113 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=9.43 $Y2=0
r202 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r203 110 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r204 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r205 107 110 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r206 106 107 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r207 104 107 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=6.67 $Y2=0
r208 103 106 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=4.37 $Y=0
+ $X2=6.67 $Y2=0
r209 103 104 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r210 101 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.37 $Y2=0
r211 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r212 98 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r213 98 129 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.07 $Y2=0
r214 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r215 95 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.155
+ $Y2=0
r216 95 97 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.99
+ $Y2=0
r217 93 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r218 93 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r219 91 115 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.7 $Y=0 $X2=9.43
+ $Y2=0
r220 91 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.7 $Y=0 $X2=9.785
+ $Y2=0
r221 90 119 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=9.87 $Y=0
+ $X2=10.35 $Y2=0
r222 90 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.87 $Y=0 $X2=9.785
+ $Y2=0
r223 88 112 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.76 $Y=0 $X2=8.51
+ $Y2=0
r224 88 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=0 $X2=8.845
+ $Y2=0
r225 87 115 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=8.93 $Y=0 $X2=9.43
+ $Y2=0
r226 87 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.93 $Y=0 $X2=8.845
+ $Y2=0
r227 85 109 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.59
+ $Y2=0
r228 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.845
+ $Y2=0
r229 84 112 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.93 $Y=0 $X2=8.51
+ $Y2=0
r230 84 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0 $X2=7.845
+ $Y2=0
r231 82 106 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.67
+ $Y2=0
r232 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.905
+ $Y2=0
r233 81 109 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.99 $Y=0 $X2=7.59
+ $Y2=0
r234 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=0 $X2=6.905
+ $Y2=0
r235 79 100 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.95 $Y=0 $X2=3.91
+ $Y2=0
r236 79 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.95 $Y=0 $X2=4.085
+ $Y2=0
r237 78 103 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.22 $Y=0 $X2=4.37
+ $Y2=0
r238 78 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.22 $Y=0 $X2=4.085
+ $Y2=0
r239 76 97 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.01 $Y=0 $X2=2.99
+ $Y2=0
r240 76 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=0 $X2=3.095
+ $Y2=0
r241 75 100 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.91
+ $Y2=0
r242 75 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.095
+ $Y2=0
r243 71 131 3.40825 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=10.725 $Y=0.085
+ $X2=10.84 $Y2=0
r244 71 73 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.725 $Y=0.085
+ $X2=10.725 $Y2=0.39
r245 67 92 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.785 $Y=0.085
+ $X2=9.785 $Y2=0
r246 67 69 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.785 $Y=0.085
+ $X2=9.785 $Y2=0.39
r247 63 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.845 $Y=0.085
+ $X2=8.845 $Y2=0
r248 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.845 $Y=0.085
+ $X2=8.845 $Y2=0.39
r249 59 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=0.085
+ $X2=7.845 $Y2=0
r250 59 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.845 $Y=0.085
+ $X2=7.845 $Y2=0.39
r251 55 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0
r252 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0.39
r253 51 80 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0
r254 51 53 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0.39
r255 47 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0
r256 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0.39
r257 43 128 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.155 $Y2=0
r258 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.155 $Y2=0.39
r259 42 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.215
+ $Y2=0
r260 41 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.155
+ $Y2=0
r261 41 42 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.3
+ $Y2=0
r262 37 125 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=0.085
+ $X2=1.215 $Y2=0
r263 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.215 $Y=0.085
+ $X2=1.215 $Y2=0.39
r264 36 122 4.29305 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.18
+ $Y2=0
r265 35 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0 $X2=1.215
+ $Y2=0
r266 35 36 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=0.36
+ $Y2=0
r267 31 122 3.02899 $w=2.75e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.222 $Y=0.085
+ $X2=0.18 $Y2=0
r268 31 33 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.222 $Y=0.085
+ $X2=0.222 $Y2=0.39
r269 10 73 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=10.59
+ $Y=0.235 $X2=10.725 $Y2=0.39
r270 9 69 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.6
+ $Y=0.235 $X2=9.785 $Y2=0.39
r271 8 65 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=8.72
+ $Y=0.235 $X2=8.845 $Y2=0.39
r272 7 61 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.66
+ $Y=0.235 $X2=7.845 $Y2=0.39
r273 6 57 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.72
+ $Y=0.235 $X2=6.905 $Y2=0.39
r274 5 53 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.85
+ $Y=0.235 $X2=4.035 $Y2=0.39
r275 4 49 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.91
+ $Y=0.235 $X2=3.095 $Y2=0.39
r276 3 45 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.235 $X2=2.155 $Y2=0.39
r277 2 39 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.215 $Y2=0.39
r278 1 33 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.275 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_4%A_886_47# 1 2 3 4 5 16 22 23 24 28 30 34 40
r92 32 34 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.29 $Y=0.725
+ $X2=8.29 $Y2=0.39
r93 31 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.54 $Y=0.815
+ $X2=7.35 $Y2=0.815
r94 30 32 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=8.1 $Y=0.815
+ $X2=8.29 $Y2=0.725
r95 30 31 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=8.1 $Y=0.815
+ $X2=7.54 $Y2=0.815
r96 26 40 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.35 $Y=0.725 $X2=7.35
+ $Y2=0.815
r97 26 28 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.35 $Y=0.725
+ $X2=7.35 $Y2=0.39
r98 25 39 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=6.6 $Y=0.815
+ $X2=6.475 $Y2=0.815
r99 24 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.16 $Y=0.815
+ $X2=7.35 $Y2=0.815
r100 24 25 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=7.16 $Y=0.815
+ $X2=6.6 $Y2=0.815
r101 23 39 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=6.475 $Y=0.725
+ $X2=6.475 $Y2=0.815
r102 22 37 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=6.475 $Y=0.475
+ $X2=6.475 $Y2=0.365
r103 22 23 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=6.475 $Y=0.475
+ $X2=6.475 $Y2=0.725
r104 18 21 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=4.555 $Y=0.365
+ $X2=5.495 $Y2=0.365
r105 16 37 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=6.35 $Y=0.365
+ $X2=6.475 $Y2=0.365
r106 16 21 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=6.35 $Y=0.365
+ $X2=5.495 $Y2=0.365
r107 5 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.18
+ $Y=0.235 $X2=8.315 $Y2=0.39
r108 4 28 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.19
+ $Y=0.235 $X2=7.375 $Y2=0.39
r109 3 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=6.3
+ $Y=0.235 $X2=6.435 $Y2=0.73
r110 3 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.3
+ $Y=0.235 $X2=6.435 $Y2=0.39
r111 2 21 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.31
+ $Y=0.235 $X2=5.495 $Y2=0.39
r112 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.235 $X2=4.555 $Y2=0.39
.ends

