* File: sky130_fd_sc_hdll__or2b_1.pex.spice
* Created: Thu Aug 27 19:23:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR2B_1%B_N 1 3 6 8 13 16
r28 13 14 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r29 11 13 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r30 8 16 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.2 $X2=0.23
+ $Y2=1.2
r31 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r32 4 14 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r33 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.475
r34 1 13 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r35 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_1%A_27_53# 1 2 9 11 13 16 18 19 22 26 29
r50 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r51 24 32 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.16
+ $X2=0.77 $Y2=1.325
r52 24 29 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.77 $Y=1.16
+ $X2=0.77 $Y2=0.82
r53 24 26 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.895 $Y=1.16
+ $X2=1.27 $Y2=1.16
r54 22 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=1.62
+ $X2=0.73 $Y2=1.325
r55 18 29 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.77 $Y2=0.82
r56 18 19 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.42 $Y2=0.82
r57 14 19 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.42 $Y2=0.82
r58 14 16 10.7809 $w=3.08e-07 $l=2.9e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.265 $Y2=0.445
r59 11 27 44.7829 $w=4.14e-07 $l=3.10242e-07 $layer=POLY_cond $X=1.505 $Y=1.41
+ $X2=1.37 $Y2=1.16
r60 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.505 $Y=1.41
+ $X2=1.505 $Y2=1.695
r61 7 27 39.8702 $w=4.14e-07 $l=2.09105e-07 $layer=POLY_cond $X=1.47 $Y=0.995
+ $X2=1.37 $Y2=1.16
r62 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.47 $Y=0.995 $X2=1.47
+ $Y2=0.475
r63 2 22 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.62
r64 1 16 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_1%A 1 3 6 9 12 14 20 24
r47 18 24 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.06 $Y=2.25
+ $X2=1.155 $Y2=2.25
r48 17 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=2.28
+ $X2=1.225 $Y2=2.28
r49 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=2.28 $X2=1.06 $Y2=2.28
r50 14 24 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.205 $Y=2.25
+ $X2=1.155 $Y2=2.25
r51 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.94 $Y=0.475
+ $X2=1.94 $Y2=1.135
r52 4 12 101.939 $w=2e-07 $l=3.05e-07 $layer=POLY_cond $X=1.915 $Y=2.035
+ $X2=1.915 $Y2=2.34
r53 4 6 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.915 $Y=2.035
+ $X2=1.915 $Y2=1.695
r54 3 11 109.045 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=1.915 $Y=1.41
+ $X2=1.915 $Y2=1.135
r55 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.915 $Y=1.41
+ $X2=1.915 $Y2=1.695
r56 1 12 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.815 $Y=2.34 $X2=1.915
+ $Y2=2.34
r57 1 20 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.815 $Y=2.34
+ $X2=1.225 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_1%A_229_297# 1 2 7 9 10 12 13 17 19 20 24 25
+ 31 33
c59 24 0 1.07404e-19 $X=2.3 $Y=1.495
r60 31 34 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=1.16
+ $X2=2.33 $Y2=1.325
r61 31 33 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=1.16
+ $X2=2.33 $Y2=0.995
r62 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.16 $X2=2.36 $Y2=1.16
r63 25 28 2.88111 $w=4.18e-07 $l=1.05e-07 $layer=LI1_cond $X=1.25 $Y=1.58
+ $X2=1.25 $Y2=1.685
r64 24 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.3 $Y=1.495 $X2=2.3
+ $Y2=1.325
r65 21 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.3 $Y=0.825 $X2=2.3
+ $Y2=0.995
r66 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=0.74
+ $X2=2.3 $Y2=0.825
r67 19 20 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.215 $Y=0.74
+ $X2=1.765 $Y2=0.74
r68 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.68 $Y=0.655
+ $X2=1.765 $Y2=0.74
r69 15 17 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.68 $Y=0.655
+ $X2=1.68 $Y2=0.47
r70 14 25 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.46 $Y=1.58 $X2=1.25
+ $Y2=1.58
r71 13 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=1.58
+ $X2=2.3 $Y2=1.495
r72 13 14 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.215 $Y=1.58
+ $X2=1.46 $Y2=1.58
r73 10 32 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.48 $Y=0.995
+ $X2=2.39 $Y2=1.16
r74 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.48 $Y=0.995
+ $X2=2.48 $Y2=0.56
r75 7 32 47.6478 $w=3.03e-07 $l=2.80624e-07 $layer=POLY_cond $X=2.455 $Y=1.41
+ $X2=2.39 $Y2=1.16
r76 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.455 $Y=1.41
+ $X2=2.455 $Y2=1.985
r77 2 28 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.485 $X2=1.27 $Y2=1.685
r78 1 17 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.545
+ $Y=0.265 $X2=1.68 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_1%VPWR 1 2 7 9 13 15 17 22 25 30
c32 2 0 1.07404e-19 $X=2.005 $Y=1.485
r33 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r34 25 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r35 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 22 30 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.345 $Y=2.72
+ $X2=2.205 $Y2=2.72
r37 22 24 13.2765 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.345 $Y=2.72
+ $X2=2.53 $Y2=2.72
r38 21 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r39 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 18 27 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r41 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 17 30 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=2.205 $Y2=2.72
r43 17 20 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 15 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r46 11 30 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=2.635
+ $X2=2.205 $Y2=2.72
r47 11 13 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.205 $Y=2.635
+ $X2=2.205 $Y2=2
r48 7 27 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r49 7 9 44.064 $w=2.53e-07 $l=9.75e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=1.66
r50 2 13 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=2.005
+ $Y=1.485 $X2=2.215 $Y2=2
r51 1 9 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_1%X 1 2 10 13 14 15 18
r18 15 18 0.616535 $w=4.83e-07 $l=2.5e-08 $layer=LI1_cond $X=2.847 $Y=1.87
+ $X2=2.847 $Y2=1.845
r19 13 18 2.66343 $w=4.83e-07 $l=1.08e-07 $layer=LI1_cond $X=2.847 $Y=1.737
+ $X2=2.847 $Y2=1.845
r20 13 14 6.51042 $w=4.83e-07 $l=2.42e-07 $layer=LI1_cond $X=2.847 $Y=1.737
+ $X2=2.847 $Y2=1.495
r21 12 14 22.0012 $w=3.83e-07 $l=7.35e-07 $layer=LI1_cond $X=2.897 $Y=0.76
+ $X2=2.897 $Y2=1.495
r22 10 12 4.7348 $w=4.83e-07 $l=1.7e-07 $layer=LI1_cond $X=2.847 $Y=0.59
+ $X2=2.847 $Y2=0.76
r23 2 18 300 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_PDIFF $count=2 $X=2.545
+ $Y=1.485 $X2=2.69 $Y2=1.845
r24 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.235 $X2=2.69 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_1%VGND 1 2 9 11 16 19 21 29 32
r39 32 35 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.15
+ $Y2=0.4
r40 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r41 28 29 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=0.24
+ $X2=1.375 $Y2=0.24
r42 25 28 1.10407 $w=6.48e-07 $l=6e-08 $layer=LI1_cond $X=1.15 $Y=0.24 $X2=1.21
+ $Y2=0.24
r43 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r44 22 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r45 21 25 8.46455 $w=6.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.24
+ $X2=1.15 $Y2=0.24
r46 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 19 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r48 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r49 16 32 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.15
+ $Y2=0
r50 16 18 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.53
+ $Y2=0
r51 15 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r52 15 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r53 14 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.375
+ $Y2=0
r54 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r55 11 32 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.15
+ $Y2=0
r56 11 14 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.61
+ $Y2=0
r57 9 22 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.69
+ $Y2=0
r58 2 35 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.265 $X2=2.2 $Y2=0.4
r59 1 28 91 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.265 $X2=1.21 $Y2=0.4
.ends

