* File: sky130_fd_sc_hdll__isobufsrc_1.spice
* Created: Wed Sep  2 08:33:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__isobufsrc_1.pex.spice"
.subckt sky130_fd_sc_hdll__isobufsrc_1  VNB VPB A SLEEP VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_74_47#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0869439 AS=0.1092 PD=0.812523 PS=1.36 NRD=32.136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_SLEEP_M1002_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.134556 PD=0.97 PS=1.25748 NRD=2.76 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A_74_47#_M1000_g N_X_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=4.608 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_74_47#_M1005_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0972507 AS=0.1134 PD=0.834085 PS=1.38 NRD=82.7991 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1001 A_283_297# N_SLEEP_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.231549 PD=1.23 PS=1.98592 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90000.4
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1003 N_X_M1003_d N_A_74_47#_M1003_g A_283_297# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.115 PD=2.54 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
pX7_noxref noxref_10 X X PROBETYPE=1
*
.include "sky130_fd_sc_hdll__isobufsrc_1.pxi.spice"
*
.ends
*
*
