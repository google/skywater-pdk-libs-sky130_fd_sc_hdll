* File: sky130_fd_sc_hdll__a22o_4.pxi.spice
* Created: Wed Sep  2 08:18:44 2020
* 
x_PM_SKY130_FD_SC_HDLL__A22O_4%A_96_21# N_A_96_21#_M1009_s N_A_96_21#_M1011_s
+ N_A_96_21#_M1012_d N_A_96_21#_M1006_d N_A_96_21#_c_106_n N_A_96_21#_M1007_g
+ N_A_96_21#_c_123_n N_A_96_21#_M1001_g N_A_96_21#_c_107_n N_A_96_21#_M1008_g
+ N_A_96_21#_c_124_n N_A_96_21#_M1005_g N_A_96_21#_c_108_n N_A_96_21#_M1013_g
+ N_A_96_21#_c_125_n N_A_96_21#_M1018_g N_A_96_21#_c_126_n N_A_96_21#_M1022_g
+ N_A_96_21#_c_109_n N_A_96_21#_M1015_g N_A_96_21#_c_110_n N_A_96_21#_c_111_n
+ N_A_96_21#_c_112_n N_A_96_21#_c_113_n N_A_96_21#_c_128_n N_A_96_21#_c_129_n
+ N_A_96_21#_c_144_p N_A_96_21#_c_114_n N_A_96_21#_c_115_n N_A_96_21#_c_116_n
+ N_A_96_21#_c_117_n N_A_96_21#_c_118_n N_A_96_21#_c_145_p N_A_96_21#_c_119_n
+ N_A_96_21#_c_120_n N_A_96_21#_c_147_p N_A_96_21#_c_121_n N_A_96_21#_c_122_n
+ PM_SKY130_FD_SC_HDLL__A22O_4%A_96_21#
x_PM_SKY130_FD_SC_HDLL__A22O_4%B2 N_B2_c_275_n N_B2_M1012_g N_B2_c_276_n
+ N_B2_M1014_g N_B2_c_277_n N_B2_M1019_g N_B2_c_278_n N_B2_M1023_g N_B2_c_283_n
+ N_B2_c_279_n B2 B2 PM_SKY130_FD_SC_HDLL__A22O_4%B2
x_PM_SKY130_FD_SC_HDLL__A22O_4%B1 N_B1_c_355_n N_B1_M1009_g N_B1_c_359_n
+ N_B1_M1003_g N_B1_c_360_n N_B1_M1006_g N_B1_c_356_n N_B1_M1016_g B1
+ N_B1_c_358_n B1 PM_SKY130_FD_SC_HDLL__A22O_4%B1
x_PM_SKY130_FD_SC_HDLL__A22O_4%A2 N_A2_c_400_n N_A2_M1002_g N_A2_c_401_n
+ N_A2_M1000_g N_A2_c_402_n N_A2_M1010_g N_A2_c_403_n N_A2_M1004_g N_A2_c_410_n
+ N_A2_c_404_n N_A2_c_405_n N_A2_c_406_n A2 A2 PM_SKY130_FD_SC_HDLL__A22O_4%A2
x_PM_SKY130_FD_SC_HDLL__A22O_4%A1 N_A1_c_475_n N_A1_M1011_g N_A1_c_478_n
+ N_A1_M1017_g N_A1_c_479_n N_A1_M1021_g N_A1_c_476_n N_A1_M1020_g A1
+ N_A1_c_477_n A1 PM_SKY130_FD_SC_HDLL__A22O_4%A1
x_PM_SKY130_FD_SC_HDLL__A22O_4%VPWR N_VPWR_M1001_s N_VPWR_M1005_s N_VPWR_M1022_s
+ N_VPWR_M1002_d N_VPWR_M1021_d N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n
+ N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n
+ N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n
+ N_VPWR_c_533_n VPWR N_VPWR_c_534_n N_VPWR_c_519_n
+ PM_SKY130_FD_SC_HDLL__A22O_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A22O_4%X N_X_M1007_d N_X_M1013_d N_X_M1001_d N_X_M1018_d
+ N_X_c_616_n N_X_c_617_n N_X_c_621_n N_X_c_622_n N_X_c_631_n N_X_c_663_n
+ N_X_c_623_n N_X_c_618_n N_X_c_646_n N_X_c_667_n N_X_c_619_n N_X_c_624_n X
+ PM_SKY130_FD_SC_HDLL__A22O_4%X
x_PM_SKY130_FD_SC_HDLL__A22O_4%A_524_297# N_A_524_297#_M1012_s
+ N_A_524_297#_M1003_s N_A_524_297#_M1023_s N_A_524_297#_M1017_s
+ N_A_524_297#_M1010_s N_A_524_297#_c_692_n N_A_524_297#_c_696_n
+ N_A_524_297#_c_711_n N_A_524_297#_c_706_n N_A_524_297#_c_736_n
+ N_A_524_297#_c_715_n N_A_524_297#_c_689_n N_A_524_297#_c_741_n
+ N_A_524_297#_c_699_n N_A_524_297#_c_700_n N_A_524_297#_c_721_n
+ PM_SKY130_FD_SC_HDLL__A22O_4%A_524_297#
x_PM_SKY130_FD_SC_HDLL__A22O_4%VGND N_VGND_M1007_s N_VGND_M1008_s N_VGND_M1015_s
+ N_VGND_M1019_d N_VGND_M1004_s N_VGND_c_748_n N_VGND_c_749_n N_VGND_c_750_n
+ N_VGND_c_751_n N_VGND_c_752_n N_VGND_c_753_n N_VGND_c_754_n N_VGND_c_755_n
+ N_VGND_c_756_n VGND N_VGND_c_757_n N_VGND_c_758_n N_VGND_c_759_n
+ N_VGND_c_760_n N_VGND_c_761_n PM_SKY130_FD_SC_HDLL__A22O_4%VGND
x_PM_SKY130_FD_SC_HDLL__A22O_4%A_616_47# N_A_616_47#_M1014_s N_A_616_47#_M1016_d
+ N_A_616_47#_c_846_n PM_SKY130_FD_SC_HDLL__A22O_4%A_616_47#
x_PM_SKY130_FD_SC_HDLL__A22O_4%A_1008_47# N_A_1008_47#_M1000_d
+ N_A_1008_47#_M1020_d N_A_1008_47#_c_862_n N_A_1008_47#_c_878_n
+ N_A_1008_47#_c_860_n PM_SKY130_FD_SC_HDLL__A22O_4%A_1008_47#
cc_1 VNB N_A_96_21#_c_106_n 0.0196598f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_2 VNB N_A_96_21#_c_107_n 0.0167602f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.995
cc_3 VNB N_A_96_21#_c_108_n 0.0171978f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.995
cc_4 VNB N_A_96_21#_c_109_n 0.0200816f $X=-0.19 $Y=-0.24 $X2=2.015 $Y2=0.995
cc_5 VNB N_A_96_21#_c_110_n 6.30857e-19 $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=1.175
cc_6 VNB N_A_96_21#_c_111_n 6.59699e-19 $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=1.785
cc_7 VNB N_A_96_21#_c_112_n 0.00481211f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=1.075
cc_8 VNB N_A_96_21#_c_113_n 2.92694e-19 $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=0.82
cc_9 VNB N_A_96_21#_c_114_n 0.00144225f $X=-0.19 $Y=-0.24 $X2=3.775 $Y2=0.775
cc_10 VNB N_A_96_21#_c_115_n 4.62713e-19 $X=-0.19 $Y=-0.24 $X2=3.55 $Y2=0.775
cc_11 VNB N_A_96_21#_c_116_n 5.08984e-19 $X=-0.19 $Y=-0.24 $X2=5.515 $Y2=0.775
cc_12 VNB N_A_96_21#_c_117_n 0.00230068f $X=-0.19 $Y=-0.24 $X2=5.645 $Y2=0.73
cc_13 VNB N_A_96_21#_c_118_n 0.00424408f $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=1.175
cc_14 VNB N_A_96_21#_c_119_n 0.0122998f $X=-0.19 $Y=-0.24 $X2=3.42 $Y2=0.775
cc_15 VNB N_A_96_21#_c_120_n 8.62268e-19 $X=-0.19 $Y=-0.24 $X2=3.905 $Y2=0.775
cc_16 VNB N_A_96_21#_c_121_n 0.0143485f $X=-0.19 $Y=-0.24 $X2=5.385 $Y2=0.775
cc_17 VNB N_A_96_21#_c_122_n 0.0801793f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=1.202
cc_18 VNB N_B2_c_275_n 0.0270651f $X=-0.19 $Y=-0.24 $X2=3.5 $Y2=0.235
cc_19 VNB N_B2_c_276_n 0.0199816f $X=-0.19 $Y=-0.24 $X2=4.01 $Y2=1.485
cc_20 VNB N_B2_c_277_n 0.0177013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B2_c_278_n 0.0222042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_B2_c_279_n 0.00350385f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.41
cc_23 VNB B2 0.00591381f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_24 VNB N_B1_c_355_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=3.5 $Y2=0.235
cc_25 VNB N_B1_c_356_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB B1 0.00141641f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_27 VNB N_B1_c_358_n 0.0356367f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_28 VNB N_A2_c_400_n 0.0222042f $X=-0.19 $Y=-0.24 $X2=3.5 $Y2=0.235
cc_29 VNB N_A2_c_401_n 0.0177013f $X=-0.19 $Y=-0.24 $X2=4.01 $Y2=1.485
cc_30 VNB N_A2_c_402_n 0.0316299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A2_c_403_n 0.0224184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A2_c_404_n 2.72331e-19 $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.41
cc_33 VNB N_A2_c_405_n 0.00360692f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.985
cc_34 VNB N_A2_c_406_n 0.00201311f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=1.985
cc_35 VNB A2 0.0211959f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=1.985
cc_36 VNB N_A1_c_475_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=3.5 $Y2=0.235
cc_37 VNB N_A1_c_476_n 0.0176182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A1_c_477_n 0.0369743f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_39 VNB N_VPWR_c_519_n 0.288713f $X=-0.19 $Y=-0.24 $X2=3.215 $Y2=1.96
cc_40 VNB N_X_c_616_n 0.0014432f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_41 VNB N_X_c_617_n 0.00986769f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_42 VNB N_X_c_618_n 0.0052859f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.985
cc_43 VNB N_X_c_619_n 0.0025225f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=1.16
cc_44 VNB X 0.0213373f $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=1.275
cc_45 VNB N_VGND_c_748_n 0.00471611f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.985
cc_46 VNB N_VGND_c_749_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=1.41
cc_47 VNB N_VGND_c_750_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.56
cc_48 VNB N_VGND_c_751_n 0.0128075f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.41
cc_49 VNB N_VGND_c_752_n 0.00674326f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.985
cc_50 VNB N_VGND_c_753_n 0.0194857f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=1.985
cc_51 VNB N_VGND_c_754_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=2.015 $Y2=0.995
cc_52 VNB N_VGND_c_755_n 0.0413233f $X=-0.19 $Y=-0.24 $X2=2.015 $Y2=0.56
cc_53 VNB N_VGND_c_756_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=1.175
cc_54 VNB N_VGND_c_757_n 0.0130399f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.16
cc_55 VNB N_VGND_c_758_n 0.0419197f $X=-0.19 $Y=-0.24 $X2=3.775 $Y2=0.775
cc_56 VNB N_VGND_c_759_n 0.0201171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_760_n 0.0208826f $X=-0.19 $Y=-0.24 $X2=4.155 $Y2=1.87
cc_58 VNB N_VGND_c_761_n 0.33739f $X=-0.19 $Y=-0.24 $X2=4.155 $Y2=1.96
cc_59 VNB N_A_1008_47#_c_860_n 0.00277337f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_60 VPB N_A_96_21#_c_123_n 0.019183f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_61 VPB N_A_96_21#_c_124_n 0.0158725f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=1.41
cc_62 VPB N_A_96_21#_c_125_n 0.0158895f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.41
cc_63 VPB N_A_96_21#_c_126_n 0.0191195f $X=-0.19 $Y=1.305 $X2=1.99 $Y2=1.41
cc_64 VPB N_A_96_21#_c_111_n 0.00827395f $X=-0.19 $Y=1.305 $X2=2.265 $Y2=1.785
cc_65 VPB N_A_96_21#_c_128_n 0.010722f $X=-0.19 $Y=1.305 $X2=3.09 $Y2=1.87
cc_66 VPB N_A_96_21#_c_129_n 0.00201536f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.87
cc_67 VPB N_A_96_21#_c_122_n 0.0467169f $X=-0.19 $Y=1.305 $X2=1.99 $Y2=1.202
cc_68 VPB N_B2_c_275_n 0.0301044f $X=-0.19 $Y=1.305 $X2=3.5 $Y2=0.235
cc_69 VPB N_B2_c_278_n 0.0256643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_B2_c_283_n 0.00683421f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_71 VPB N_B2_c_279_n 0.00272944f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_72 VPB B2 0.00314111f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=0.56
cc_73 VPB N_B1_c_359_n 0.0159948f $X=-0.19 $Y=1.305 $X2=4.01 $Y2=1.485
cc_74 VPB N_B1_c_360_n 0.0159958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_B1_c_358_n 0.0192932f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=0.56
cc_76 VPB N_A2_c_400_n 0.0256643f $X=-0.19 $Y=1.305 $X2=3.5 $Y2=0.235
cc_77 VPB N_A2_c_402_n 0.0331355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A2_c_410_n 0.00767987f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_79 VPB N_A2_c_404_n 0.00130718f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_80 VPB N_A2_c_405_n 0.00272944f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.985
cc_81 VPB N_A1_c_478_n 0.0159779f $X=-0.19 $Y=1.305 $X2=4.01 $Y2=1.485
cc_82 VPB N_A1_c_479_n 0.0159751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A1_c_477_n 0.0192923f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=0.56
cc_84 VPB N_VPWR_c_520_n 0.0140014f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_85 VPB N_VPWR_c_521_n 0.00518f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.985
cc_86 VPB N_VPWR_c_522_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=1.41
cc_87 VPB N_VPWR_c_523_n 0.00518f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=0.56
cc_88 VPB N_VPWR_c_524_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.985
cc_89 VPB N_VPWR_c_525_n 0.00516582f $X=-0.19 $Y=1.305 $X2=2.015 $Y2=0.995
cc_90 VPB N_VPWR_c_526_n 0.0195604f $X=-0.19 $Y=1.305 $X2=2.1 $Y2=1.175
cc_91 VPB N_VPWR_c_527_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.175
cc_92 VPB N_VPWR_c_528_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_93 VPB N_VPWR_c_529_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_530_n 0.064513f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.16
cc_95 VPB N_VPWR_c_531_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.16
cc_96 VPB N_VPWR_c_532_n 0.0195604f $X=-0.19 $Y=1.305 $X2=2.265 $Y2=1.785
cc_97 VPB N_VPWR_c_533_n 0.0047828f $X=-0.19 $Y=1.305 $X2=2.285 $Y2=0.905
cc_98 VPB N_VPWR_c_534_n 0.021236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_519_n 0.0546338f $X=-0.19 $Y=1.305 $X2=3.215 $Y2=1.96
cc_100 VPB N_X_c_621_n 0.00163065f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.56
cc_101 VPB N_X_c_622_n 0.0124524f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_102 VPB N_X_c_623_n 0.0037826f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=0.56
cc_103 VPB N_X_c_624_n 0.00150464f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.16
cc_104 VPB X 0.00761414f $X=-0.19 $Y=1.305 $X2=2.265 $Y2=1.275
cc_105 VPB N_A_524_297#_c_689_n 0.00341263f $X=-0.19 $Y=1.305 $X2=2.015
+ $Y2=0.995
cc_106 N_A_96_21#_c_111_n N_B2_c_275_n 0.00615701f $X=2.265 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_96_21#_c_112_n N_B2_c_275_n 0.00249961f $X=2.285 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_96_21#_c_128_n N_B2_c_275_n 0.0130414f $X=3.09 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_96_21#_c_118_n N_B2_c_275_n 0.00100694f $X=2.265 $Y=1.175 $X2=-0.19
+ $Y2=-0.24
cc_110 N_A_96_21#_c_119_n N_B2_c_275_n 0.00437142f $X=3.42 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_96_21#_c_112_n N_B2_c_276_n 0.00229864f $X=2.285 $Y=1.075 $X2=0 $Y2=0
cc_112 N_A_96_21#_c_115_n N_B2_c_276_n 4.83332e-19 $X=3.55 $Y=0.775 $X2=0 $Y2=0
cc_113 N_A_96_21#_c_119_n N_B2_c_276_n 0.0135212f $X=3.42 $Y=0.775 $X2=0 $Y2=0
cc_114 N_A_96_21#_c_120_n N_B2_c_277_n 4.42559e-19 $X=3.905 $Y=0.775 $X2=0 $Y2=0
cc_115 N_A_96_21#_c_121_n N_B2_c_277_n 0.0126763f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_116 N_A_96_21#_c_121_n N_B2_c_278_n 0.00437142f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_117 N_A_96_21#_M1012_d N_B2_c_283_n 0.00135043f $X=3.07 $Y=1.485 $X2=0 $Y2=0
cc_118 N_A_96_21#_M1006_d N_B2_c_283_n 0.00171997f $X=4.01 $Y=1.485 $X2=0 $Y2=0
cc_119 N_A_96_21#_c_144_p N_B2_c_283_n 0.0371166f $X=4.03 $Y=1.87 $X2=0 $Y2=0
cc_120 N_A_96_21#_c_145_p N_B2_c_283_n 0.00754343f $X=3.215 $Y=1.87 $X2=0 $Y2=0
cc_121 N_A_96_21#_c_119_n N_B2_c_283_n 0.0113406f $X=3.42 $Y=0.775 $X2=0 $Y2=0
cc_122 N_A_96_21#_c_147_p N_B2_c_283_n 0.0102375f $X=4.155 $Y=1.87 $X2=0 $Y2=0
cc_123 N_A_96_21#_M1006_d N_B2_c_279_n 7.75307e-19 $X=4.01 $Y=1.485 $X2=0 $Y2=0
cc_124 N_A_96_21#_c_147_p N_B2_c_279_n 0.00353817f $X=4.155 $Y=1.87 $X2=0 $Y2=0
cc_125 N_A_96_21#_c_121_n N_B2_c_279_n 0.0293526f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_126 N_A_96_21#_M1012_d B2 0.00115658f $X=3.07 $Y=1.485 $X2=0 $Y2=0
cc_127 N_A_96_21#_c_111_n B2 0.0270954f $X=2.265 $Y=1.785 $X2=0 $Y2=0
cc_128 N_A_96_21#_c_128_n B2 0.0303443f $X=3.09 $Y=1.87 $X2=0 $Y2=0
cc_129 N_A_96_21#_c_118_n B2 0.0170506f $X=2.265 $Y=1.175 $X2=0 $Y2=0
cc_130 N_A_96_21#_c_145_p B2 0.00648665f $X=3.215 $Y=1.87 $X2=0 $Y2=0
cc_131 N_A_96_21#_c_119_n B2 0.0463411f $X=3.42 $Y=0.775 $X2=0 $Y2=0
cc_132 N_A_96_21#_c_122_n B2 9.93151e-19 $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_133 N_A_96_21#_c_115_n N_B1_c_355_n 0.00578232f $X=3.55 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_96_21#_c_119_n N_B1_c_355_n 0.00539089f $X=3.42 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_96_21#_c_144_p N_B1_c_359_n 0.0108425f $X=4.03 $Y=1.87 $X2=0 $Y2=0
cc_136 N_A_96_21#_c_144_p N_B1_c_360_n 0.0108425f $X=4.03 $Y=1.87 $X2=0 $Y2=0
cc_137 N_A_96_21#_c_120_n N_B1_c_356_n 0.00351953f $X=3.905 $Y=0.775 $X2=0 $Y2=0
cc_138 N_A_96_21#_c_121_n N_B1_c_356_n 0.00720497f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_139 N_A_96_21#_c_119_n B1 0.0474637f $X=3.42 $Y=0.775 $X2=0 $Y2=0
cc_140 N_A_96_21#_c_114_n N_B1_c_358_n 0.00473056f $X=3.775 $Y=0.775 $X2=0 $Y2=0
cc_141 N_A_96_21#_c_121_n N_A2_c_400_n 0.00437142f $X=5.385 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_142 N_A_96_21#_c_116_n N_A2_c_401_n 4.7941e-19 $X=5.515 $Y=0.775 $X2=0 $Y2=0
cc_143 N_A_96_21#_c_121_n N_A2_c_401_n 0.0122477f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_144 N_A_96_21#_c_121_n N_A2_c_410_n 0.00717126f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_145 N_A_96_21#_c_121_n N_A2_c_405_n 0.0293526f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_146 N_A_96_21#_c_116_n N_A1_c_475_n 0.005477f $X=5.515 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_96_21#_c_121_n N_A1_c_475_n 0.00580546f $X=5.385 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_148 N_A_96_21#_c_117_n N_A1_c_476_n 4.134e-19 $X=5.645 $Y=0.73 $X2=0 $Y2=0
cc_149 N_A_96_21#_c_121_n A1 0.0338603f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_150 N_A_96_21#_c_117_n N_A1_c_477_n 0.0047334f $X=5.645 $Y=0.73 $X2=0 $Y2=0
cc_151 N_A_96_21#_c_111_n N_VPWR_M1022_s 0.00352509f $X=2.265 $Y=1.785 $X2=0
+ $Y2=0
cc_152 N_A_96_21#_c_129_n N_VPWR_M1022_s 0.00430391f $X=2.43 $Y=1.87 $X2=0 $Y2=0
cc_153 N_A_96_21#_c_123_n N_VPWR_c_521_n 0.00479105f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_96_21#_c_124_n N_VPWR_c_522_n 0.00300743f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_96_21#_c_125_n N_VPWR_c_522_n 0.00300743f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_96_21#_c_126_n N_VPWR_c_523_n 0.00479105f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_96_21#_c_129_n N_VPWR_c_523_n 0.0185141f $X=2.43 $Y=1.87 $X2=0 $Y2=0
cc_158 N_A_96_21#_c_123_n N_VPWR_c_526_n 0.00702461f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_96_21#_c_124_n N_VPWR_c_526_n 0.00702461f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_96_21#_c_125_n N_VPWR_c_528_n 0.00702461f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_96_21#_c_126_n N_VPWR_c_528_n 0.00702461f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_96_21#_M1012_d N_VPWR_c_519_n 0.00231289f $X=3.07 $Y=1.485 $X2=0
+ $Y2=0
cc_163 N_A_96_21#_M1006_d N_VPWR_c_519_n 0.00232092f $X=4.01 $Y=1.485 $X2=0
+ $Y2=0
cc_164 N_A_96_21#_c_123_n N_VPWR_c_519_n 0.0133906f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_96_21#_c_124_n N_VPWR_c_519_n 0.0124092f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_96_21#_c_125_n N_VPWR_c_519_n 0.0124092f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_96_21#_c_126_n N_VPWR_c_519_n 0.0136915f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_96_21#_c_128_n N_VPWR_c_519_n 0.0079376f $X=3.09 $Y=1.87 $X2=0 $Y2=0
cc_169 N_A_96_21#_c_129_n N_VPWR_c_519_n 0.00435471f $X=2.43 $Y=1.87 $X2=0 $Y2=0
cc_170 N_A_96_21#_c_144_p N_VPWR_c_519_n 0.00153883f $X=4.03 $Y=1.87 $X2=0 $Y2=0
cc_171 N_A_96_21#_c_106_n N_X_c_616_n 0.0111251f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_96_21#_c_110_n N_X_c_616_n 0.00410208f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_173 N_A_96_21#_c_123_n N_X_c_621_n 0.0178749f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_96_21#_c_110_n N_X_c_621_n 0.0103328f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_175 N_A_96_21#_c_122_n N_X_c_621_n 9.44081e-19 $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_176 N_A_96_21#_c_106_n N_X_c_631_n 0.0109499f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_96_21#_c_107_n N_X_c_631_n 0.00676224f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_96_21#_c_108_n N_X_c_631_n 5.42233e-19 $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_96_21#_c_124_n N_X_c_623_n 0.0157513f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_96_21#_c_125_n N_X_c_623_n 0.015669f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_96_21#_c_126_n N_X_c_623_n 4.00176e-19 $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_96_21#_c_110_n N_X_c_623_n 0.0689039f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_183 N_A_96_21#_c_111_n N_X_c_623_n 0.00287394f $X=2.265 $Y=1.785 $X2=0 $Y2=0
cc_184 N_A_96_21#_c_122_n N_X_c_623_n 0.0151889f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_185 N_A_96_21#_c_107_n N_X_c_618_n 0.00901745f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_96_21#_c_108_n N_X_c_618_n 0.010179f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_96_21#_c_109_n N_X_c_618_n 2.14781e-19 $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_96_21#_c_110_n N_X_c_618_n 0.0704813f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_189 N_A_96_21#_c_113_n N_X_c_618_n 0.00148154f $X=2.43 $Y=0.82 $X2=0 $Y2=0
cc_190 N_A_96_21#_c_122_n N_X_c_618_n 0.00831812f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_191 N_A_96_21#_c_107_n N_X_c_646_n 5.24597e-19 $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_96_21#_c_108_n N_X_c_646_n 0.00651696f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_96_21#_c_106_n N_X_c_619_n 0.00116607f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_96_21#_c_107_n N_X_c_619_n 0.00116607f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_96_21#_c_110_n N_X_c_619_n 0.0305614f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_196 N_A_96_21#_c_122_n N_X_c_619_n 0.00358132f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_197 N_A_96_21#_c_110_n N_X_c_624_n 0.020385f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_198 N_A_96_21#_c_122_n N_X_c_624_n 0.00664519f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_199 N_A_96_21#_c_106_n X 0.0186818f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_96_21#_c_123_n X 0.00133332f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_96_21#_c_110_n X 0.0164324f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_202 N_A_96_21#_c_128_n N_A_524_297#_M1012_s 0.00528269f $X=3.09 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_203 N_A_96_21#_c_144_p N_A_524_297#_M1003_s 0.00347905f $X=4.03 $Y=1.87 $X2=0
+ $Y2=0
cc_204 N_A_96_21#_M1012_d N_A_524_297#_c_692_n 0.0035039f $X=3.07 $Y=1.485 $X2=0
+ $Y2=0
cc_205 N_A_96_21#_c_128_n N_A_524_297#_c_692_n 0.00608347f $X=3.09 $Y=1.87 $X2=0
+ $Y2=0
cc_206 N_A_96_21#_c_144_p N_A_524_297#_c_692_n 0.00608347f $X=4.03 $Y=1.87 $X2=0
+ $Y2=0
cc_207 N_A_96_21#_c_145_p N_A_524_297#_c_692_n 0.0126551f $X=3.215 $Y=1.87 $X2=0
+ $Y2=0
cc_208 N_A_96_21#_M1006_d N_A_524_297#_c_696_n 0.0035039f $X=4.01 $Y=1.485 $X2=0
+ $Y2=0
cc_209 N_A_96_21#_c_144_p N_A_524_297#_c_696_n 0.00608347f $X=4.03 $Y=1.87 $X2=0
+ $Y2=0
cc_210 N_A_96_21#_c_147_p N_A_524_297#_c_696_n 0.0126551f $X=4.155 $Y=1.87 $X2=0
+ $Y2=0
cc_211 N_A_96_21#_c_128_n N_A_524_297#_c_699_n 0.0158267f $X=3.09 $Y=1.87 $X2=0
+ $Y2=0
cc_212 N_A_96_21#_c_144_p N_A_524_297#_c_700_n 0.0131392f $X=4.03 $Y=1.87 $X2=0
+ $Y2=0
cc_213 N_A_96_21#_c_113_n N_VGND_M1015_s 0.0054889f $X=2.43 $Y=0.82 $X2=0 $Y2=0
cc_214 N_A_96_21#_c_119_n N_VGND_M1015_s 0.00771529f $X=3.42 $Y=0.775 $X2=0
+ $Y2=0
cc_215 N_A_96_21#_c_121_n N_VGND_M1019_d 0.00574611f $X=5.385 $Y=0.775 $X2=0
+ $Y2=0
cc_216 N_A_96_21#_c_106_n N_VGND_c_748_n 0.00438629f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_217 N_A_96_21#_c_107_n N_VGND_c_749_n 0.00394736f $X=1.025 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_96_21#_c_108_n N_VGND_c_749_n 0.00276126f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_96_21#_c_121_n N_VGND_c_750_n 0.0125492f $X=5.385 $Y=0.775 $X2=0
+ $Y2=0
cc_220 N_A_96_21#_c_106_n N_VGND_c_753_n 0.00423737f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_96_21#_c_107_n N_VGND_c_753_n 0.00423737f $X=1.025 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_96_21#_c_119_n N_VGND_c_755_n 0.00195107f $X=3.42 $Y=0.775 $X2=0
+ $Y2=0
cc_223 N_A_96_21#_c_121_n N_VGND_c_755_n 0.00324501f $X=5.385 $Y=0.775 $X2=0
+ $Y2=0
cc_224 N_A_96_21#_c_121_n N_VGND_c_758_n 0.00244779f $X=5.385 $Y=0.775 $X2=0
+ $Y2=0
cc_225 N_A_96_21#_c_108_n N_VGND_c_759_n 0.00423334f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_96_21#_c_109_n N_VGND_c_759_n 0.00585385f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_96_21#_c_109_n N_VGND_c_760_n 0.00481673f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_96_21#_c_113_n N_VGND_c_760_n 0.0232224f $X=2.43 $Y=0.82 $X2=0 $Y2=0
cc_229 N_A_96_21#_c_119_n N_VGND_c_760_n 0.0297002f $X=3.42 $Y=0.775 $X2=0 $Y2=0
cc_230 N_A_96_21#_M1009_s N_VGND_c_761_n 0.00297142f $X=3.5 $Y=0.235 $X2=0 $Y2=0
cc_231 N_A_96_21#_M1011_s N_VGND_c_761_n 0.00297142f $X=5.46 $Y=0.235 $X2=0
+ $Y2=0
cc_232 N_A_96_21#_c_106_n N_VGND_c_761_n 0.00687004f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_96_21#_c_107_n N_VGND_c_761_n 0.0060934f $X=1.025 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_96_21#_c_108_n N_VGND_c_761_n 0.00608558f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_96_21#_c_109_n N_VGND_c_761_n 0.012103f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_96_21#_c_113_n N_VGND_c_761_n 0.00127084f $X=2.43 $Y=0.82 $X2=0 $Y2=0
cc_237 N_A_96_21#_c_119_n N_VGND_c_761_n 0.00655867f $X=3.42 $Y=0.775 $X2=0
+ $Y2=0
cc_238 N_A_96_21#_c_121_n N_VGND_c_761_n 0.0140014f $X=5.385 $Y=0.775 $X2=0
+ $Y2=0
cc_239 N_A_96_21#_c_119_n N_A_616_47#_M1014_s 0.00195168f $X=3.42 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_240 N_A_96_21#_c_121_n N_A_616_47#_M1016_d 0.00195168f $X=5.385 $Y=0.775
+ $X2=0 $Y2=0
cc_241 N_A_96_21#_M1009_s N_A_616_47#_c_846_n 0.00507817f $X=3.5 $Y=0.235 $X2=0
+ $Y2=0
cc_242 N_A_96_21#_c_115_n N_A_616_47#_c_846_n 0.0262985f $X=3.55 $Y=0.775 $X2=0
+ $Y2=0
cc_243 N_A_96_21#_c_119_n N_A_616_47#_c_846_n 0.0143855f $X=3.42 $Y=0.775 $X2=0
+ $Y2=0
cc_244 N_A_96_21#_c_121_n N_A_616_47#_c_846_n 0.0141607f $X=5.385 $Y=0.775 $X2=0
+ $Y2=0
cc_245 N_A_96_21#_c_121_n N_A_1008_47#_M1000_d 0.00195168f $X=5.385 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_246 N_A_96_21#_M1011_s N_A_1008_47#_c_862_n 0.00507817f $X=5.46 $Y=0.235
+ $X2=0 $Y2=0
cc_247 N_A_96_21#_c_116_n N_A_1008_47#_c_862_n 0.0236512f $X=5.515 $Y=0.775
+ $X2=0 $Y2=0
cc_248 N_A_96_21#_c_121_n N_A_1008_47#_c_862_n 0.0146102f $X=5.385 $Y=0.775
+ $X2=0 $Y2=0
cc_249 N_A_96_21#_c_117_n N_A_1008_47#_c_860_n 6.50328e-19 $X=5.645 $Y=0.73
+ $X2=0 $Y2=0
cc_250 N_B2_c_276_n N_B1_c_355_n 0.0268717f $X=3.005 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_251 N_B2_c_275_n N_B1_c_359_n 0.036701f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B2_c_283_n N_B1_c_359_n 0.0112877f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_253 B2 N_B1_c_359_n 0.00115622f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_254 N_B2_c_278_n N_B1_c_360_n 0.0367147f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B2_c_283_n N_B1_c_360_n 0.011241f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_256 N_B2_c_279_n N_B1_c_360_n 0.00101445f $X=4.365 $Y=1.16 $X2=0 $Y2=0
cc_257 N_B2_c_277_n N_B1_c_356_n 0.0269111f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B2_c_275_n B1 2.06946e-19 $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B2_c_278_n B1 6.86695e-19 $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B2_c_283_n B1 0.0461557f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_261 N_B2_c_279_n B1 0.0176354f $X=4.365 $Y=1.16 $X2=0 $Y2=0
cc_262 B2 B1 0.0173147f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_263 N_B2_c_275_n N_B1_c_358_n 0.0263618f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B2_c_278_n N_B1_c_358_n 0.0263033f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B2_c_283_n N_B1_c_358_n 0.00803891f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_266 N_B2_c_279_n N_B1_c_358_n 0.00392336f $X=4.365 $Y=1.16 $X2=0 $Y2=0
cc_267 B2 N_B1_c_358_n 0.00510434f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_268 N_B2_c_278_n N_A2_c_400_n 0.040024f $X=4.39 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_269 N_B2_c_279_n N_A2_c_400_n 0.00168165f $X=4.365 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_270 N_B2_c_277_n N_A2_c_401_n 0.0222335f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_271 N_B2_c_278_n N_A2_c_405_n 0.00168165f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B2_c_279_n N_A2_c_405_n 0.0455154f $X=4.365 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B2_c_275_n N_VPWR_c_523_n 0.00213395f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B2_c_275_n N_VPWR_c_530_n 0.00429453f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B2_c_278_n N_VPWR_c_530_n 0.00429453f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B2_c_275_n N_VPWR_c_519_n 0.00737353f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B2_c_278_n N_VPWR_c_519_n 0.00629441f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_278 B2 N_A_524_297#_M1012_s 0.00420446f $X=2.905 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_279 N_B2_c_283_n N_A_524_297#_M1003_s 0.00187547f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_280 N_B2_c_279_n N_A_524_297#_M1023_s 0.00161069f $X=4.365 $Y=1.16 $X2=0
+ $Y2=0
cc_281 N_B2_c_275_n N_A_524_297#_c_692_n 0.0099733f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_282 N_B2_c_278_n N_A_524_297#_c_696_n 0.0143148f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_283 N_B2_c_279_n N_A_524_297#_c_706_n 0.00372315f $X=4.365 $Y=1.16 $X2=0
+ $Y2=0
cc_284 N_B2_c_277_n N_VGND_c_750_n 0.00664414f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B2_c_276_n N_VGND_c_755_n 0.00395831f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B2_c_277_n N_VGND_c_755_n 0.0042294f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B2_c_276_n N_VGND_c_760_n 0.00770185f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B2_c_276_n N_VGND_c_761_n 0.0069348f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B2_c_277_n N_VGND_c_761_n 0.00636233f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B2_c_276_n N_A_616_47#_c_846_n 0.00518052f $X=3.005 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_B2_c_277_n N_A_616_47#_c_846_n 0.00359207f $X=4.365 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_B1_c_359_n N_VPWR_c_530_n 0.00429453f $X=3.45 $Y=1.41 $X2=0 $Y2=0
cc_293 N_B1_c_360_n N_VPWR_c_530_n 0.00429453f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_294 N_B1_c_359_n N_VPWR_c_519_n 0.00609118f $X=3.45 $Y=1.41 $X2=0 $Y2=0
cc_295 N_B1_c_360_n N_VPWR_c_519_n 0.00609118f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_296 N_B1_c_359_n N_A_524_297#_c_692_n 0.0099733f $X=3.45 $Y=1.41 $X2=0 $Y2=0
cc_297 N_B1_c_360_n N_A_524_297#_c_696_n 0.0099733f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_298 N_B1_c_355_n N_VGND_c_755_n 0.00357877f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B1_c_356_n N_VGND_c_755_n 0.00357877f $X=3.945 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B1_c_355_n N_VGND_c_761_n 0.005504f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B1_c_356_n N_VGND_c_761_n 0.005504f $X=3.945 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B1_c_355_n N_A_616_47#_c_846_n 0.00989193f $X=3.425 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_B1_c_356_n N_A_616_47#_c_846_n 0.0100513f $X=3.945 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A2_c_401_n N_A1_c_475_n 0.0268761f $X=4.965 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_305 N_A2_c_400_n N_A1_c_478_n 0.0371417f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A2_c_410_n N_A1_c_478_n 0.0116479f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_307 N_A2_c_405_n N_A1_c_478_n 0.00101445f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A2_c_402_n N_A1_c_479_n 0.0364739f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A2_c_410_n N_A1_c_479_n 0.0141145f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_310 N_A2_c_404_n N_A1_c_479_n 7.34002e-19 $X=6.2 $Y=1.445 $X2=0 $Y2=0
cc_311 N_A2_c_403_n N_A1_c_476_n 0.0103419f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A2_c_400_n A1 2.20488e-19 $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_313 N_A2_c_410_n A1 0.0384921f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_314 N_A2_c_405_n A1 0.0136034f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A2_c_406_n A1 0.0143347f $X=6.285 $Y=1.175 $X2=0 $Y2=0
cc_316 N_A2_c_400_n N_A1_c_477_n 0.0264727f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A2_c_402_n N_A1_c_477_n 0.026336f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A2_c_410_n N_A1_c_477_n 0.00821086f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_319 N_A2_c_404_n N_A1_c_477_n 0.0029218f $X=6.2 $Y=1.445 $X2=0 $Y2=0
cc_320 N_A2_c_405_n N_A1_c_477_n 0.00464862f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A2_c_406_n N_A1_c_477_n 0.00163966f $X=6.285 $Y=1.175 $X2=0 $Y2=0
cc_322 N_A2_c_410_n N_VPWR_M1002_d 0.00172342f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_323 N_A2_c_405_n N_VPWR_M1002_d 7.76441e-19 $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A2_c_410_n N_VPWR_M1021_d 0.00189646f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_325 N_A2_c_400_n N_VPWR_c_524_n 0.00300743f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A2_c_402_n N_VPWR_c_525_n 0.00300743f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A2_c_400_n N_VPWR_c_530_n 0.00702461f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A2_c_402_n N_VPWR_c_534_n 0.00702461f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_329 N_A2_c_400_n N_VPWR_c_519_n 0.00716301f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_330 N_A2_c_402_n N_VPWR_c_519_n 0.00791853f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_331 N_A2_c_405_n N_A_524_297#_M1023_s 0.00161069f $X=4.915 $Y=1.16 $X2=0
+ $Y2=0
cc_332 N_A2_c_410_n N_A_524_297#_M1017_s 0.00187091f $X=6.115 $Y=1.53 $X2=0
+ $Y2=0
cc_333 N_A2_c_400_n N_A_524_297#_c_711_n 0.011385f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_334 N_A2_c_410_n N_A_524_297#_c_711_n 0.0218268f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_335 N_A2_c_405_n N_A_524_297#_c_711_n 0.0167698f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A2_c_405_n N_A_524_297#_c_706_n 0.00372315f $X=4.915 $Y=1.16 $X2=0
+ $Y2=0
cc_337 N_A2_c_402_n N_A_524_297#_c_715_n 0.0139685f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_338 N_A2_c_410_n N_A_524_297#_c_715_n 0.0273762f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_339 A2 N_A_524_297#_c_715_n 0.00534422f $X=6.575 $Y=1.105 $X2=0 $Y2=0
cc_340 N_A2_c_402_n N_A_524_297#_c_689_n 0.004595f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A2_c_410_n N_A_524_297#_c_689_n 0.0104762f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_342 A2 N_A_524_297#_c_689_n 0.0166332f $X=6.575 $Y=1.105 $X2=0 $Y2=0
cc_343 N_A2_c_410_n N_A_524_297#_c_721_n 0.0143191f $X=6.115 $Y=1.53 $X2=0 $Y2=0
cc_344 N_A2_c_401_n N_VGND_c_750_n 0.00660142f $X=4.965 $Y=0.995 $X2=0 $Y2=0
cc_345 N_A2_c_402_n N_VGND_c_752_n 2.29969e-19 $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A2_c_403_n N_VGND_c_752_n 0.00461082f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_347 A2 N_VGND_c_752_n 0.0137431f $X=6.575 $Y=1.105 $X2=0 $Y2=0
cc_348 N_A2_c_401_n N_VGND_c_758_n 0.00395831f $X=4.965 $Y=0.995 $X2=0 $Y2=0
cc_349 N_A2_c_403_n N_VGND_c_758_n 0.00585385f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_350 N_A2_c_401_n N_VGND_c_761_n 0.00607592f $X=4.965 $Y=0.995 $X2=0 $Y2=0
cc_351 N_A2_c_403_n N_VGND_c_761_n 0.0116855f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_352 N_A2_c_401_n N_A_1008_47#_c_862_n 0.00530312f $X=4.965 $Y=0.995 $X2=0
+ $Y2=0
cc_353 N_A2_c_402_n N_A_1008_47#_c_860_n 0.00235635f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A2_c_410_n N_A_1008_47#_c_860_n 0.00310205f $X=6.115 $Y=1.53 $X2=0
+ $Y2=0
cc_355 N_A2_c_406_n N_A_1008_47#_c_860_n 0.014037f $X=6.285 $Y=1.175 $X2=0 $Y2=0
cc_356 N_A1_c_478_n N_VPWR_c_524_n 0.00300743f $X=5.41 $Y=1.41 $X2=0 $Y2=0
cc_357 N_A1_c_479_n N_VPWR_c_525_n 0.00300743f $X=5.88 $Y=1.41 $X2=0 $Y2=0
cc_358 N_A1_c_478_n N_VPWR_c_532_n 0.00702461f $X=5.41 $Y=1.41 $X2=0 $Y2=0
cc_359 N_A1_c_479_n N_VPWR_c_532_n 0.00702461f $X=5.88 $Y=1.41 $X2=0 $Y2=0
cc_360 N_A1_c_478_n N_VPWR_c_519_n 0.00695979f $X=5.41 $Y=1.41 $X2=0 $Y2=0
cc_361 N_A1_c_479_n N_VPWR_c_519_n 0.00695979f $X=5.88 $Y=1.41 $X2=0 $Y2=0
cc_362 N_A1_c_478_n N_A_524_297#_c_711_n 0.011229f $X=5.41 $Y=1.41 $X2=0 $Y2=0
cc_363 N_A1_c_479_n N_A_524_297#_c_715_n 0.011229f $X=5.88 $Y=1.41 $X2=0 $Y2=0
cc_364 N_A1_c_475_n N_VGND_c_758_n 0.00357877f $X=5.385 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A1_c_476_n N_VGND_c_758_n 0.00357877f $X=5.905 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A1_c_475_n N_VGND_c_761_n 0.005504f $X=5.385 $Y=0.995 $X2=0 $Y2=0
cc_367 N_A1_c_476_n N_VGND_c_761_n 0.00562222f $X=5.905 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A1_c_475_n N_A_1008_47#_c_862_n 0.00990963f $X=5.385 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A1_c_476_n N_A_1008_47#_c_862_n 0.0132083f $X=5.905 $Y=0.995 $X2=0
+ $Y2=0
cc_370 A1 N_A_1008_47#_c_862_n 0.00184847f $X=5.66 $Y=1.105 $X2=0 $Y2=0
cc_371 N_VPWR_c_519_n N_X_M1001_d 0.00370124f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_372 N_VPWR_c_519_n N_X_M1018_d 0.00370124f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_373 N_VPWR_M1001_s N_X_c_621_n 7.22239e-19 $X=0.2 $Y=1.485 $X2=0 $Y2=0
cc_374 N_VPWR_c_521_n N_X_c_621_n 0.00434858f $X=0.345 $Y=1.99 $X2=0 $Y2=0
cc_375 N_VPWR_M1001_s N_X_c_622_n 0.00354732f $X=0.2 $Y=1.485 $X2=0 $Y2=0
cc_376 N_VPWR_c_521_n N_X_c_622_n 0.011469f $X=0.345 $Y=1.99 $X2=0 $Y2=0
cc_377 N_VPWR_c_526_n N_X_c_663_n 0.0149311f $X=1.16 $Y=2.72 $X2=0 $Y2=0
cc_378 N_VPWR_c_519_n N_X_c_663_n 0.00955092f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_379 N_VPWR_M1005_s N_X_c_623_n 0.00191634f $X=1.14 $Y=1.485 $X2=0 $Y2=0
cc_380 N_VPWR_c_522_n N_X_c_623_n 0.0137198f $X=1.285 $Y=1.99 $X2=0 $Y2=0
cc_381 N_VPWR_c_528_n N_X_c_667_n 0.0149311f $X=2.1 $Y=2.72 $X2=0 $Y2=0
cc_382 N_VPWR_c_519_n N_X_c_667_n 0.00955092f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_c_519_n N_A_524_297#_M1012_s 0.00215913f $X=6.67 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_384 N_VPWR_c_519_n N_A_524_297#_M1003_s 0.00229658f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_519_n N_A_524_297#_M1023_s 0.00306083f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_519_n N_A_524_297#_M1017_s 0.00250817f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_519_n N_A_524_297#_M1010_s 0.00363111f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_530_n N_A_524_297#_c_692_n 0.0386534f $X=5.05 $Y=2.72 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_519_n N_A_524_297#_c_692_n 0.0239144f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_530_n N_A_524_297#_c_696_n 0.0592811f $X=5.05 $Y=2.72 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_519_n N_A_524_297#_c_696_n 0.0366233f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_392 N_VPWR_M1002_d N_A_524_297#_c_711_n 0.00367036f $X=5.03 $Y=1.485 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_524_n N_A_524_297#_c_711_n 0.0138319f $X=5.175 $Y=2.3 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_519_n N_A_524_297#_c_711_n 0.0141583f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_532_n N_A_524_297#_c_736_n 0.0149311f $X=5.99 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_519_n N_A_524_297#_c_736_n 0.00955092f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_397 N_VPWR_M1021_d N_A_524_297#_c_715_n 0.00369025f $X=5.97 $Y=1.485 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_525_n N_A_524_297#_c_715_n 0.0139109f $X=6.115 $Y=2.3 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_519_n N_A_524_297#_c_715_n 0.0158107f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_534_n N_A_524_297#_c_741_n 0.0142751f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_519_n N_A_524_297#_c_741_n 0.00781789f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_523_n N_A_524_297#_c_699_n 0.0186128f $X=2.225 $Y=2.3 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_530_n N_A_524_297#_c_699_n 0.0154637f $X=5.05 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_519_n N_A_524_297#_c_699_n 0.00938745f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_530_n N_A_524_297#_c_700_n 0.014332f $X=5.05 $Y=2.72 $X2=0 $Y2=0
cc_406 N_VPWR_c_519_n N_A_524_297#_c_700_n 0.00938745f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_X_c_616_n N_VGND_M1007_s 5.40298e-19 $X=0.6 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_408 N_X_c_617_n N_VGND_M1007_s 0.00329182f $X=0.37 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_409 N_X_c_618_n N_VGND_M1008_s 0.00251047f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_410 N_X_c_616_n N_VGND_c_748_n 0.00402428f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_411 N_X_c_617_n N_VGND_c_748_n 0.00920832f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_412 N_X_c_631_n N_VGND_c_749_n 0.0177507f $X=0.815 $Y=0.39 $X2=0 $Y2=0
cc_413 N_X_c_618_n N_VGND_c_749_n 0.0127273f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_414 N_X_c_631_n N_VGND_c_753_n 0.0210053f $X=0.815 $Y=0.39 $X2=0 $Y2=0
cc_415 N_X_c_618_n N_VGND_c_753_n 0.00266636f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_416 N_X_c_616_n N_VGND_c_757_n 0.0019947f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_417 N_X_c_617_n N_VGND_c_757_n 0.00293744f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_418 N_X_c_618_n N_VGND_c_759_n 0.00198695f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_419 N_X_c_646_n N_VGND_c_759_n 0.0231806f $X=1.755 $Y=0.39 $X2=0 $Y2=0
cc_420 N_X_M1007_d N_VGND_c_761_n 0.00255747f $X=0.63 $Y=0.235 $X2=0 $Y2=0
cc_421 N_X_M1013_d N_VGND_c_761_n 0.00364931f $X=1.57 $Y=0.235 $X2=0 $Y2=0
cc_422 N_X_c_616_n N_VGND_c_761_n 0.00407016f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_423 N_X_c_617_n N_VGND_c_761_n 0.00542613f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_424 N_X_c_631_n N_VGND_c_761_n 0.0140539f $X=0.815 $Y=0.39 $X2=0 $Y2=0
cc_425 N_X_c_618_n N_VGND_c_761_n 0.00972452f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_426 N_X_c_646_n N_VGND_c_761_n 0.0143352f $X=1.755 $Y=0.39 $X2=0 $Y2=0
cc_427 N_VGND_c_761_n N_A_616_47#_M1014_s 0.00215227f $X=6.67 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_428 N_VGND_c_761_n N_A_616_47#_M1016_d 0.00215227f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_750_n N_A_616_47#_c_846_n 0.0121537f $X=4.67 $Y=0.39 $X2=0 $Y2=0
cc_430 N_VGND_c_755_n N_A_616_47#_c_846_n 0.0742459f $X=4.585 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_760_n N_A_616_47#_c_846_n 0.0190752f $X=2.83 $Y=0.235 $X2=0
+ $Y2=0
cc_432 N_VGND_c_761_n N_A_616_47#_c_846_n 0.0472891f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_433 N_VGND_c_761_n N_A_1008_47#_M1000_d 0.00215227f $X=6.67 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_434 N_VGND_c_761_n N_A_1008_47#_M1020_d 0.00321315f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_750_n N_A_1008_47#_c_862_n 0.0148152f $X=4.67 $Y=0.39 $X2=0
+ $Y2=0
cc_436 N_VGND_c_758_n N_A_1008_47#_c_862_n 0.0600765f $X=6.5 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_761_n N_A_1008_47#_c_862_n 0.0381287f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_438 N_VGND_c_758_n N_A_1008_47#_c_878_n 0.015983f $X=6.5 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_c_761_n N_A_1008_47#_c_878_n 0.00961275f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_752_n N_A_1008_47#_c_860_n 5.82165e-19 $X=6.585 $Y=0.39 $X2=0
+ $Y2=0
