* File: sky130_fd_sc_hdll__nor2b_1.spice
* Created: Thu Aug 27 19:15:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor2b_1.pex.spice"
.subckt sky130_fd_sc_hdll__nor2b_1  VNB VPB B_N A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_B_N_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.113714 AS=0.1092 PD=0.918505 PS=1.36 NRD=55.704 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.175986 PD=0.92 PS=1.4215 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A_27_47#_M1002_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_B_N_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.108431 AS=0.1134 PD=0.887324 PS=1.38 NRD=95.2889 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1000 A_253_297# N_A_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.258169 PD=1.23 PS=2.11268 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90000.5
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1004 N_Y_M1004_d N_A_27_47#_M1004_g A_253_297# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.115 PD=2.54 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.9
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
pX7_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__nor2b_1.pxi.spice"
*
.ends
*
*
