* File: sky130_fd_sc_hdll__xor3_1.pxi.spice
* Created: Wed Sep  2 08:54:45 2020
* 
x_PM_SKY130_FD_SC_HDLL__XOR3_1%A_116_21# N_A_116_21#_M1007_d N_A_116_21#_M1005_d
+ N_A_116_21#_c_158_n N_A_116_21#_M1018_g N_A_116_21#_c_159_n
+ N_A_116_21#_M1019_g N_A_116_21#_c_160_n N_A_116_21#_c_171_p
+ N_A_116_21#_c_205_p N_A_116_21#_c_176_p N_A_116_21#_c_214_p
+ N_A_116_21#_c_161_n N_A_116_21#_c_166_n N_A_116_21#_c_162_n
+ N_A_116_21#_c_167_n N_A_116_21#_c_168_n N_A_116_21#_c_181_p
+ N_A_116_21#_c_163_n PM_SKY130_FD_SC_HDLL__XOR3_1%A_116_21#
x_PM_SKY130_FD_SC_HDLL__XOR3_1%C N_C_c_260_n N_C_M1002_g N_C_M1001_g N_C_c_261_n
+ N_C_c_262_n N_C_M1005_g N_C_c_263_n N_C_M1007_g N_C_c_264_n C N_C_c_265_n C
+ PM_SKY130_FD_SC_HDLL__XOR3_1%C
x_PM_SKY130_FD_SC_HDLL__XOR3_1%A_276_93# N_A_276_93#_M1002_d N_A_276_93#_M1001_d
+ N_A_276_93#_c_324_n N_A_276_93#_M1017_g N_A_276_93#_c_325_n
+ N_A_276_93#_M1020_g N_A_276_93#_c_340_n N_A_276_93#_c_326_n
+ N_A_276_93#_c_330_n N_A_276_93#_c_331_n N_A_276_93#_c_332_n
+ N_A_276_93#_c_327_n PM_SKY130_FD_SC_HDLL__XOR3_1%A_276_93#
x_PM_SKY130_FD_SC_HDLL__XOR3_1%A_875_297# N_A_875_297#_M1003_d
+ N_A_875_297#_M1006_d N_A_875_297#_c_413_n N_A_875_297#_M1015_g
+ N_A_875_297#_M1008_g N_A_875_297#_c_400_n N_A_875_297#_c_415_n
+ N_A_875_297#_M1010_g N_A_875_297#_M1014_g N_A_875_297#_c_401_n
+ N_A_875_297#_c_402_n N_A_875_297#_c_418_n N_A_875_297#_c_403_n
+ N_A_875_297#_c_404_n N_A_875_297#_c_422_p N_A_875_297#_c_405_n
+ N_A_875_297#_c_406_n N_A_875_297#_c_407_n N_A_875_297#_c_408_n
+ N_A_875_297#_c_409_n N_A_875_297#_c_410_n N_A_875_297#_c_411_n
+ N_A_875_297#_c_412_n PM_SKY130_FD_SC_HDLL__XOR3_1%A_875_297#
x_PM_SKY130_FD_SC_HDLL__XOR3_1%B N_B_c_588_n N_B_M1006_g N_B_M1003_g N_B_c_581_n
+ N_B_c_582_n N_B_M1011_g N_B_M1004_g N_B_c_591_n N_B_c_592_n N_B_M1009_g
+ N_B_c_593_n N_B_c_594_n N_B_M1012_g N_B_c_584_n N_B_c_597_n N_B_c_585_n
+ N_B_c_586_n B B N_B_c_587_n PM_SKY130_FD_SC_HDLL__XOR3_1%B
x_PM_SKY130_FD_SC_HDLL__XOR3_1%A N_A_c_717_n N_A_M1016_g N_A_c_718_n N_A_M1000_g
+ A A PM_SKY130_FD_SC_HDLL__XOR3_1%A
x_PM_SKY130_FD_SC_HDLL__XOR3_1%A_991_365# N_A_991_365#_M1004_s
+ N_A_991_365#_M1014_d N_A_991_365#_M1011_s N_A_991_365#_M1010_d
+ N_A_991_365#_c_754_n N_A_991_365#_M1013_g N_A_991_365#_c_755_n
+ N_A_991_365#_M1021_g N_A_991_365#_c_756_n N_A_991_365#_c_764_n
+ N_A_991_365#_c_757_n N_A_991_365#_c_758_n N_A_991_365#_c_759_n
+ N_A_991_365#_c_766_n N_A_991_365#_c_776_n N_A_991_365#_c_760_n
+ N_A_991_365#_c_761_n N_A_991_365#_c_789_n N_A_991_365#_c_790_n
+ PM_SKY130_FD_SC_HDLL__XOR3_1%A_991_365#
x_PM_SKY130_FD_SC_HDLL__XOR3_1%X N_X_M1018_s N_X_M1019_s N_X_c_883_n N_X_c_885_n
+ N_X_c_884_n X PM_SKY130_FD_SC_HDLL__XOR3_1%X
x_PM_SKY130_FD_SC_HDLL__XOR3_1%VPWR N_VPWR_M1019_d N_VPWR_M1006_s N_VPWR_M1016_d
+ N_VPWR_c_908_n N_VPWR_c_909_n N_VPWR_c_910_n VPWR N_VPWR_c_911_n
+ N_VPWR_c_912_n N_VPWR_c_907_n N_VPWR_c_914_n N_VPWR_c_915_n N_VPWR_c_916_n
+ N_VPWR_c_917_n PM_SKY130_FD_SC_HDLL__XOR3_1%VPWR
x_PM_SKY130_FD_SC_HDLL__XOR3_1%A_406_325# N_A_406_325#_M1020_d
+ N_A_406_325#_M1009_d N_A_406_325#_M1005_s N_A_406_325#_M1011_d
+ N_A_406_325#_c_1006_n N_A_406_325#_c_1026_n N_A_406_325#_c_1004_n
+ N_A_406_325#_c_1008_n N_A_406_325#_c_1043_n N_A_406_325#_c_1009_n
+ N_A_406_325#_c_1005_n N_A_406_325#_c_1137_p N_A_406_325#_c_1056_n
+ N_A_406_325#_c_1057_n N_A_406_325#_c_1078_n N_A_406_325#_c_1011_n
+ N_A_406_325#_c_1012_n N_A_406_325#_c_1013_n N_A_406_325#_c_1014_n
+ PM_SKY130_FD_SC_HDLL__XOR3_1%A_406_325#
x_PM_SKY130_FD_SC_HDLL__XOR3_1%A_424_49# N_A_424_49#_M1007_s N_A_424_49#_M1004_d
+ N_A_424_49#_M1017_d N_A_424_49#_M1012_d N_A_424_49#_c_1151_n
+ N_A_424_49#_c_1175_n N_A_424_49#_c_1152_n N_A_424_49#_c_1176_n
+ N_A_424_49#_c_1158_n N_A_424_49#_c_1159_n N_A_424_49#_c_1160_n
+ N_A_424_49#_c_1153_n N_A_424_49#_c_1154_n N_A_424_49#_c_1162_n
+ N_A_424_49#_c_1163_n N_A_424_49#_c_1164_n N_A_424_49#_c_1165_n
+ N_A_424_49#_c_1155_n N_A_424_49#_c_1167_n N_A_424_49#_c_1212_n
+ N_A_424_49#_c_1168_n N_A_424_49#_c_1156_n N_A_424_49#_c_1169_n
+ N_A_424_49#_c_1157_n N_A_424_49#_c_1170_n
+ PM_SKY130_FD_SC_HDLL__XOR3_1%A_424_49#
x_PM_SKY130_FD_SC_HDLL__XOR3_1%A_1276_297# N_A_1276_297#_M1008_d
+ N_A_1276_297#_M1021_d N_A_1276_297#_M1015_d N_A_1276_297#_M1013_d
+ N_A_1276_297#_c_1338_n N_A_1276_297#_c_1350_n N_A_1276_297#_c_1342_n
+ N_A_1276_297#_c_1339_n N_A_1276_297#_c_1351_n N_A_1276_297#_c_1344_n
+ N_A_1276_297#_c_1340_n PM_SKY130_FD_SC_HDLL__XOR3_1%A_1276_297#
x_PM_SKY130_FD_SC_HDLL__XOR3_1%VGND N_VGND_M1018_d N_VGND_M1003_s N_VGND_M1000_d
+ N_VGND_c_1404_n N_VGND_c_1405_n N_VGND_c_1406_n N_VGND_c_1407_n
+ N_VGND_c_1408_n N_VGND_c_1409_n N_VGND_c_1410_n VGND N_VGND_c_1411_n
+ N_VGND_c_1412_n N_VGND_c_1413_n N_VGND_c_1414_n
+ PM_SKY130_FD_SC_HDLL__XOR3_1%VGND
cc_1 VNB N_A_116_21#_c_158_n 0.0243567f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=0.995
cc_2 VNB N_A_116_21#_c_159_n 0.0374016f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.41
cc_3 VNB N_A_116_21#_c_160_n 0.00196712f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.16
cc_4 VNB N_A_116_21#_c_161_n 0.00138296f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.695
cc_5 VNB N_A_116_21#_c_162_n 0.00284376f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=0.34
cc_6 VNB N_A_116_21#_c_163_n 0.0162324f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.355
cc_7 VNB N_C_c_260_n 0.0199005f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=0.245
cc_8 VNB N_C_c_261_n 0.0556119f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=0.56
cc_9 VNB N_C_c_262_n 0.012954f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.41
cc_10 VNB N_C_c_263_n 0.0220325f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.865
cc_11 VNB N_C_c_264_n 0.0118441f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.16
cc_12 VNB N_C_c_265_n 0.00241009f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.425
cc_13 VNB N_A_276_93#_c_324_n 0.0267993f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=0.995
cc_14 VNB N_A_276_93#_c_325_n 0.021936f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.41
cc_15 VNB N_A_276_93#_c_326_n 0.00270273f $X=-0.19 $Y=-0.24 $X2=1.23 $Y2=0.78
cc_16 VNB N_A_276_93#_c_327_n 0.00242696f $X=-0.19 $Y=-0.24 $X2=1.57 $Y2=2.32
cc_17 VNB N_A_875_297#_M1008_g 0.0360507f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.985
cc_18 VNB N_A_875_297#_c_400_n 0.00170012f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.16
cc_19 VNB N_A_875_297#_c_401_n 0.0291447f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.425
cc_20 VNB N_A_875_297#_c_402_n 0.0176862f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.695
cc_21 VNB N_A_875_297#_c_403_n 0.00235412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_875_297#_c_404_n 0.00793619f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_875_297#_c_405_n 0.0128101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_875_297#_c_406_n 0.00135073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_875_297#_c_407_n 0.00305701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_875_297#_c_408_n 0.00216737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_875_297#_c_409_n 0.00613074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_875_297#_c_410_n 0.0286378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_875_297#_c_411_n 0.0195573f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_875_297#_c_412_n 0.00253923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_B_M1003_g 0.0302293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_B_c_581_n 0.0556994f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=0.56
cc_33 VNB N_B_c_582_n 0.0314753f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=0.56
cc_34 VNB N_B_M1004_g 0.0287687f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.16
cc_35 VNB N_B_c_584_n 0.0103656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_B_c_585_n 0.00131401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_B_c_586_n 0.0298429f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.16
cc_38 VNB N_B_c_587_n 0.0212173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_c_717_n 0.0263989f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=0.245
cc_40 VNB N_A_c_718_n 0.0204135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB A 0.0071675f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=0.995
cc_42 VNB N_A_991_365#_c_754_n 0.0299638f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.865
cc_43 VNB N_A_991_365#_c_755_n 0.0219208f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.16
cc_44 VNB N_A_991_365#_c_756_n 0.00635833f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.96
cc_45 VNB N_A_991_365#_c_757_n 0.00616113f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=0.34
cc_46 VNB N_A_991_365#_c_758_n 0.00201667f $X=-0.19 $Y=-0.24 $X2=1.57 $Y2=2.32
cc_47 VNB N_A_991_365#_c_759_n 0.00453988f $X=-0.19 $Y=-0.24 $X2=2.73 $Y2=2.32
cc_48 VNB N_A_991_365#_c_760_n 0.0020298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_991_365#_c_761_n 0.00505355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_X_c_883_n 0.0314184f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.41
cc_51 VNB N_X_c_884_n 0.0213326f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.16
cc_52 VNB N_VPWR_c_907_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_406_325#_c_1004_n 0.00971866f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.96
cc_54 VNB N_A_406_325#_c_1005_n 0.0097913f $X=-0.19 $Y=-0.24 $X2=2.73 $Y2=2.32
cc_55 VNB N_A_424_49#_c_1151_n 0.00264617f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.865
cc_56 VNB N_A_424_49#_c_1152_n 0.00850511f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.78
cc_57 VNB N_A_424_49#_c_1153_n 0.014051f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.34
cc_58 VNB N_A_424_49#_c_1154_n 0.00304946f $X=-0.19 $Y=-0.24 $X2=1.57 $Y2=2.32
cc_59 VNB N_A_424_49#_c_1155_n 0.00223545f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.16
cc_60 VNB N_A_424_49#_c_1156_n 0.0107916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_424_49#_c_1157_n 3.37974e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1276_297#_c_1338_n 0.00788636f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.16
cc_63 VNB N_A_1276_297#_c_1339_n 0.0307904f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.34
cc_64 VNB N_A_1276_297#_c_1340_n 0.0135316f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.16
cc_65 VNB N_VGND_c_1404_n 0.00516754f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.985
cc_66 VNB N_VGND_c_1405_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.16
cc_67 VNB N_VGND_c_1406_n 0.00630126f $X=-0.19 $Y=-0.24 $X2=1.35 $Y2=1.96
cc_68 VNB N_VGND_c_1407_n 0.0239542f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.695
cc_69 VNB N_VGND_c_1408_n 0.00478003f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=2.045
cc_70 VNB N_VGND_c_1409_n 0.0718762f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.34
cc_71 VNB N_VGND_c_1410_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=0.34
cc_72 VNB N_VGND_c_1411_n 0.109008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1412_n 0.0217413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1413_n 0.485301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1414_n 0.00862767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VPB N_A_116_21#_c_159_n 0.0395413f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.41
cc_77 VPB N_A_116_21#_c_160_n 0.00282905f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.16
cc_78 VPB N_A_116_21#_c_166_n 0.0038652f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=2.235
cc_79 VPB N_A_116_21#_c_167_n 0.00112766f $X=-0.19 $Y=1.305 $X2=1.57 $Y2=2.32
cc_80 VPB N_A_116_21#_c_168_n 0.0127396f $X=-0.19 $Y=1.305 $X2=2.73 $Y2=2.32
cc_81 VPB N_C_M1001_g 0.0323013f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=0.995
cc_82 VPB N_C_c_261_n 0.0253556f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=0.56
cc_83 VPB N_C_c_262_n 0.0395735f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.41
cc_84 VPB N_C_c_264_n 0.00718176f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.16
cc_85 VPB N_C_c_265_n 6.20239e-19 $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.425
cc_86 VPB N_A_276_93#_c_324_n 0.0399465f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=0.995
cc_87 VPB N_A_276_93#_c_326_n 0.00446988f $X=-0.19 $Y=1.305 $X2=1.23 $Y2=0.78
cc_88 VPB N_A_276_93#_c_330_n 0.0160663f $X=-0.19 $Y=1.305 $X2=1.35 $Y2=1.96
cc_89 VPB N_A_276_93#_c_331_n 0.00230347f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.695
cc_90 VPB N_A_276_93#_c_332_n 0.00173244f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=2.045
cc_91 VPB N_A_276_93#_c_327_n 2.71983e-19 $X=-0.19 $Y=1.305 $X2=1.57 $Y2=2.32
cc_92 VPB N_A_875_297#_c_413_n 0.0204741f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=0.995
cc_93 VPB N_A_875_297#_c_400_n 0.0104627f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.16
cc_94 VPB N_A_875_297#_c_415_n 0.0239536f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.16
cc_95 VPB N_A_875_297#_c_401_n 0.0105828f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.425
cc_96 VPB N_A_875_297#_c_402_n 0.00766961f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.695
cc_97 VPB N_A_875_297#_c_418_n 0.00591035f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=0.34
cc_98 VPB N_A_875_297#_c_412_n 0.0032041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_B_c_588_n 0.0216572f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=0.245
cc_100 VPB N_B_c_582_n 0.00747973f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=0.56
cc_101 VPB N_B_M1011_g 0.0155329f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.865
cc_102 VPB N_B_c_591_n 0.12486f $X=-0.19 $Y=1.305 $X2=1.23 $Y2=0.78
cc_103 VPB N_B_c_592_n 0.0170126f $X=-0.19 $Y=1.305 $X2=1 $Y2=0.78
cc_104 VPB N_B_c_593_n 0.0101708f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=2.045
cc_105 VPB N_B_c_594_n 0.00717497f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=2.235
cc_106 VPB N_B_M1012_g 0.0130358f $X=-0.19 $Y=1.305 $X2=1.57 $Y2=2.32
cc_107 VPB N_B_c_584_n 0.0087608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_B_c_597_n 0.00185689f $X=-0.19 $Y=1.305 $X2=2.725 $Y2=0.37
cc_109 VPB N_B_c_585_n 9.77983e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_B_c_586_n 0.0052573f $X=-0.19 $Y=1.305 $X2=0.8 $Y2=1.16
cc_111 VPB B 0.00366663f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_c_717_n 0.0298442f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=0.245
cc_113 VPB A 0.00364213f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=0.995
cc_114 VPB N_A_991_365#_c_754_n 0.0317993f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.865
cc_115 VPB N_A_991_365#_c_756_n 0.00273235f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.96
cc_116 VPB N_A_991_365#_c_764_n 0.00176559f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.695
cc_117 VPB N_A_991_365#_c_759_n 3.10649e-19 $X=-0.19 $Y=1.305 $X2=2.73 $Y2=2.32
cc_118 VPB N_A_991_365#_c_766_n 0.00206695f $X=-0.19 $Y=1.305 $X2=2.73 $Y2=2.32
cc_119 VPB N_X_c_885_n 0.0149648f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.16
cc_120 VPB N_X_c_884_n 0.00739754f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.16
cc_121 VPB X 0.0376478f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.16
cc_122 VPB N_VPWR_c_908_n 0.00957549f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.985
cc_123 VPB N_VPWR_c_909_n 0.0663405f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.875
cc_124 VPB N_VPWR_c_910_n 0.00804433f $X=-0.19 $Y=1.305 $X2=1.23 $Y2=0.78
cc_125 VPB N_VPWR_c_911_n 0.0233903f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.425
cc_126 VPB N_VPWR_c_912_n 0.0167157f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_907_n 0.073642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_914_n 0.00641289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_915_n 0.00513206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_916_n 0.096063f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_917_n 0.0124813f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_406_325#_c_1006_n 0.00306017f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.865
cc_133 VPB N_A_406_325#_c_1004_n 0.00164253f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.96
cc_134 VPB N_A_406_325#_c_1008_n 0.00270715f $X=-0.19 $Y=1.305 $X2=1.34
+ $Y2=0.695
cc_135 VPB N_A_406_325#_c_1009_n 8.62277e-19 $X=-0.19 $Y=1.305 $X2=1.45 $Y2=0.34
cc_136 VPB N_A_406_325#_c_1005_n 0.0021572f $X=-0.19 $Y=1.305 $X2=2.73 $Y2=2.32
cc_137 VPB N_A_406_325#_c_1011_n 0.0148089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_406_325#_c_1012_n 0.00318502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_406_325#_c_1013_n 0.0015478f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_406_325#_c_1014_n 0.0215932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_424_49#_c_1158_n 0.0026444f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.425
cc_142 VPB N_A_424_49#_c_1159_n 0.00579762f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.695
cc_143 VPB N_A_424_49#_c_1160_n 8.62166e-19 $X=-0.19 $Y=1.305 $X2=1.46 $Y2=2.045
cc_144 VPB N_A_424_49#_c_1154_n 0.00847729f $X=-0.19 $Y=1.305 $X2=1.57 $Y2=2.32
cc_145 VPB N_A_424_49#_c_1162_n 0.00306425f $X=-0.19 $Y=1.305 $X2=2.73 $Y2=2.32
cc_146 VPB N_A_424_49#_c_1163_n 0.00298222f $X=-0.19 $Y=1.305 $X2=2.725
+ $Y2=0.355
cc_147 VPB N_A_424_49#_c_1164_n 0.0103424f $X=-0.19 $Y=1.305 $X2=2.725 $Y2=0.37
cc_148 VPB N_A_424_49#_c_1165_n 0.00185607f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=0.355
cc_149 VPB N_A_424_49#_c_1155_n 0.00149669f $X=-0.19 $Y=1.305 $X2=0.8 $Y2=1.16
cc_150 VPB N_A_424_49#_c_1167_n 0.024688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_424_49#_c_1168_n 0.00221665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_424_49#_c_1169_n 2.86933e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_424_49#_c_1170_n 3.79061e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_1276_297#_c_1338_n 0.00457449f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.16
cc_155 VPB N_A_1276_297#_c_1342_n 0.0147295f $X=-0.19 $Y=1.305 $X2=1.34
+ $Y2=0.695
cc_156 VPB N_A_1276_297#_c_1339_n 0.0229985f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=0.34
cc_157 VPB N_A_1276_297#_c_1344_n 0.0101148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 N_A_116_21#_c_158_n N_C_c_260_n 0.0111306f $X=0.655 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_116_21#_c_160_n N_C_c_260_n 0.0014397f $X=0.885 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_116_21#_c_171_p N_C_c_260_n 0.0124376f $X=1.23 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A_116_21#_c_161_n N_C_c_260_n 0.0108052f $X=1.34 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_162 N_A_116_21#_c_162_n N_C_c_260_n 0.00580453f $X=1.45 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_163 N_A_116_21#_c_159_n N_C_M1001_g 0.0186386f $X=0.68 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_116_21#_c_160_n N_C_M1001_g 0.00568058f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_116_21#_c_176_p N_C_M1001_g 0.0133767f $X=1.35 $Y=1.96 $X2=0 $Y2=0
cc_166 N_A_116_21#_c_166_n N_C_M1001_g 0.00763977f $X=1.46 $Y=2.235 $X2=0 $Y2=0
cc_167 N_A_116_21#_c_167_n N_C_M1001_g 0.00747755f $X=1.57 $Y=2.32 $X2=0 $Y2=0
cc_168 N_A_116_21#_c_163_n N_C_c_261_n 0.010701f $X=2.49 $Y=0.355 $X2=0 $Y2=0
cc_169 N_A_116_21#_c_168_n N_C_c_262_n 0.0112964f $X=2.73 $Y=2.32 $X2=0 $Y2=0
cc_170 N_A_116_21#_c_181_p N_C_c_263_n 0.00537539f $X=2.725 $Y=0.37 $X2=0 $Y2=0
cc_171 N_A_116_21#_c_163_n N_C_c_263_n 0.00603149f $X=2.49 $Y=0.355 $X2=0 $Y2=0
cc_172 N_A_116_21#_c_159_n N_C_c_264_n 0.0248618f $X=0.68 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_116_21#_c_160_n N_C_c_264_n 0.00252038f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_116_21#_c_163_n N_C_c_265_n 0.00331115f $X=2.49 $Y=0.355 $X2=0 $Y2=0
cc_175 N_A_116_21#_c_171_p N_A_276_93#_M1002_d 0.00214828f $X=1.23 $Y=0.78
+ $X2=-0.19 $Y2=-0.24
cc_176 N_A_116_21#_c_161_n N_A_276_93#_M1002_d 0.00618081f $X=1.34 $Y=0.695
+ $X2=-0.19 $Y2=-0.24
cc_177 N_A_116_21#_c_176_p N_A_276_93#_M1001_d 0.00436734f $X=1.35 $Y=1.96 $X2=0
+ $Y2=0
cc_178 N_A_116_21#_c_166_n N_A_276_93#_M1001_d 0.00269214f $X=1.46 $Y=2.235
+ $X2=0 $Y2=0
cc_179 N_A_116_21#_c_168_n N_A_276_93#_c_324_n 0.00841967f $X=2.73 $Y=2.32 $X2=0
+ $Y2=0
cc_180 N_A_116_21#_c_181_p N_A_276_93#_c_325_n 0.00165143f $X=2.725 $Y=0.37
+ $X2=0 $Y2=0
cc_181 N_A_116_21#_c_171_p N_A_276_93#_c_340_n 0.00402121f $X=1.23 $Y=0.78 $X2=0
+ $Y2=0
cc_182 N_A_116_21#_c_176_p N_A_276_93#_c_340_n 0.0200253f $X=1.35 $Y=1.96 $X2=0
+ $Y2=0
cc_183 N_A_116_21#_c_168_n N_A_276_93#_c_340_n 0.00160427f $X=2.73 $Y=2.32 $X2=0
+ $Y2=0
cc_184 N_A_116_21#_c_159_n N_A_276_93#_c_326_n 6.8931e-19 $X=0.68 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_116_21#_c_160_n N_A_276_93#_c_326_n 0.0179148f $X=0.885 $Y=1.16 $X2=0
+ $Y2=0
cc_186 N_A_116_21#_c_171_p N_A_276_93#_c_326_n 0.0137799f $X=1.23 $Y=0.78 $X2=0
+ $Y2=0
cc_187 N_A_116_21#_c_161_n N_A_276_93#_c_326_n 0.00736858f $X=1.34 $Y=0.695
+ $X2=0 $Y2=0
cc_188 N_A_116_21#_c_163_n N_A_276_93#_c_326_n 0.0130244f $X=2.49 $Y=0.355 $X2=0
+ $Y2=0
cc_189 N_A_116_21#_M1005_d N_A_276_93#_c_330_n 0.00327687f $X=2.54 $Y=1.625
+ $X2=0 $Y2=0
cc_190 N_A_116_21#_c_168_n N_A_276_93#_c_330_n 0.00614909f $X=2.73 $Y=2.32 $X2=0
+ $Y2=0
cc_191 N_A_116_21#_c_168_n N_A_276_93#_c_332_n 0.00632099f $X=2.73 $Y=2.32 $X2=0
+ $Y2=0
cc_192 N_A_116_21#_c_158_n N_X_c_883_n 0.0119755f $X=0.655 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_116_21#_c_160_n N_X_c_883_n 0.00396341f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_116_21#_c_205_p N_X_c_883_n 0.012246f $X=1 $Y=0.78 $X2=0 $Y2=0
cc_195 N_A_116_21#_c_161_n N_X_c_883_n 0.00423537f $X=1.34 $Y=0.695 $X2=0 $Y2=0
cc_196 N_A_116_21#_c_159_n N_X_c_885_n 0.0053372f $X=0.68 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_116_21#_c_160_n N_X_c_885_n 0.0175614f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_116_21#_c_158_n N_X_c_884_n 0.0107344f $X=0.655 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_116_21#_c_160_n N_X_c_884_n 0.0170239f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_116_21#_c_159_n X 0.0108044f $X=0.68 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_116_21#_c_160_n N_VPWR_M1019_d 0.0080216f $X=0.885 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_202 N_A_116_21#_c_176_p N_VPWR_M1019_d 0.00908042f $X=1.35 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_203 N_A_116_21#_c_214_p N_VPWR_M1019_d 0.00342876f $X=1 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_204 N_A_116_21#_c_159_n N_VPWR_c_908_n 0.0086641f $X=0.68 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_116_21#_c_176_p N_VPWR_c_908_n 0.0126462f $X=1.35 $Y=1.96 $X2=0 $Y2=0
cc_206 N_A_116_21#_c_214_p N_VPWR_c_908_n 0.0143755f $X=1 $Y=1.96 $X2=0 $Y2=0
cc_207 N_A_116_21#_c_166_n N_VPWR_c_908_n 0.00141178f $X=1.46 $Y=2.235 $X2=0
+ $Y2=0
cc_208 N_A_116_21#_c_167_n N_VPWR_c_908_n 0.0133539f $X=1.57 $Y=2.32 $X2=0 $Y2=0
cc_209 N_A_116_21#_c_176_p N_VPWR_c_909_n 0.00241968f $X=1.35 $Y=1.96 $X2=0
+ $Y2=0
cc_210 N_A_116_21#_c_167_n N_VPWR_c_909_n 0.0109705f $X=1.57 $Y=2.32 $X2=0 $Y2=0
cc_211 N_A_116_21#_c_168_n N_VPWR_c_909_n 0.0642605f $X=2.73 $Y=2.32 $X2=0 $Y2=0
cc_212 N_A_116_21#_c_159_n N_VPWR_c_911_n 0.00673617f $X=0.68 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_116_21#_c_214_p N_VPWR_c_911_n 2.83092e-19 $X=1 $Y=1.96 $X2=0 $Y2=0
cc_214 N_A_116_21#_c_159_n N_VPWR_c_907_n 0.0142968f $X=0.68 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_116_21#_c_176_p N_VPWR_c_907_n 0.00567317f $X=1.35 $Y=1.96 $X2=0
+ $Y2=0
cc_216 N_A_116_21#_c_214_p N_VPWR_c_907_n 0.00170623f $X=1 $Y=1.96 $X2=0 $Y2=0
cc_217 N_A_116_21#_c_167_n N_VPWR_c_907_n 0.00809357f $X=1.57 $Y=2.32 $X2=0
+ $Y2=0
cc_218 N_A_116_21#_c_168_n N_VPWR_c_907_n 0.0515593f $X=2.73 $Y=2.32 $X2=0 $Y2=0
cc_219 N_A_116_21#_c_168_n N_A_406_325#_M1005_s 0.00721138f $X=2.73 $Y=2.32
+ $X2=0 $Y2=0
cc_220 N_A_116_21#_M1005_d N_A_406_325#_c_1006_n 0.00649326f $X=2.54 $Y=1.625
+ $X2=0 $Y2=0
cc_221 N_A_116_21#_c_176_p N_A_406_325#_c_1006_n 0.00740552f $X=1.35 $Y=1.96
+ $X2=0 $Y2=0
cc_222 N_A_116_21#_c_166_n N_A_406_325#_c_1006_n 8.52135e-19 $X=1.46 $Y=2.235
+ $X2=0 $Y2=0
cc_223 N_A_116_21#_c_168_n N_A_406_325#_c_1006_n 0.0612998f $X=2.73 $Y=2.32
+ $X2=0 $Y2=0
cc_224 N_A_116_21#_c_163_n N_A_424_49#_M1007_s 0.00669207f $X=2.49 $Y=0.355
+ $X2=-0.19 $Y2=-0.24
cc_225 N_A_116_21#_M1007_d N_A_424_49#_c_1151_n 0.0130594f $X=2.59 $Y=0.245
+ $X2=0 $Y2=0
cc_226 N_A_116_21#_c_181_p N_A_424_49#_c_1151_n 0.0203761f $X=2.725 $Y=0.37
+ $X2=0 $Y2=0
cc_227 N_A_116_21#_c_163_n N_A_424_49#_c_1151_n 0.0191047f $X=2.49 $Y=0.355
+ $X2=0 $Y2=0
cc_228 N_A_116_21#_c_181_p N_A_424_49#_c_1175_n 0.002195f $X=2.725 $Y=0.37 $X2=0
+ $Y2=0
cc_229 N_A_116_21#_c_181_p N_A_424_49#_c_1176_n 0.0147713f $X=2.725 $Y=0.37
+ $X2=0 $Y2=0
cc_230 N_A_116_21#_c_168_n N_A_424_49#_c_1168_n 0.0100105f $X=2.73 $Y=2.32 $X2=0
+ $Y2=0
cc_231 N_A_116_21#_c_160_n N_VGND_M1018_d 4.50328e-19 $X=0.885 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_232 N_A_116_21#_c_171_p N_VGND_M1018_d 0.00907954f $X=1.23 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_233 N_A_116_21#_c_205_p N_VGND_M1018_d 0.00512088f $X=1 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_234 N_A_116_21#_c_158_n N_VGND_c_1404_n 0.0103401f $X=0.655 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_116_21#_c_159_n N_VGND_c_1404_n 8.1672e-19 $X=0.68 $Y=1.41 $X2=0
+ $Y2=0
cc_236 N_A_116_21#_c_171_p N_VGND_c_1404_n 0.00454809f $X=1.23 $Y=0.78 $X2=0
+ $Y2=0
cc_237 N_A_116_21#_c_205_p N_VGND_c_1404_n 0.0162144f $X=1 $Y=0.78 $X2=0 $Y2=0
cc_238 N_A_116_21#_c_161_n N_VGND_c_1404_n 0.00733827f $X=1.34 $Y=0.695 $X2=0
+ $Y2=0
cc_239 N_A_116_21#_c_162_n N_VGND_c_1404_n 0.014093f $X=1.45 $Y=0.34 $X2=0 $Y2=0
cc_240 N_A_116_21#_c_158_n N_VGND_c_1407_n 0.00572867f $X=0.655 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_116_21#_c_171_p N_VGND_c_1409_n 0.0022086f $X=1.23 $Y=0.78 $X2=0
+ $Y2=0
cc_242 N_A_116_21#_c_162_n N_VGND_c_1409_n 0.0156439f $X=1.45 $Y=0.34 $X2=0
+ $Y2=0
cc_243 N_A_116_21#_c_163_n N_VGND_c_1409_n 0.0886428f $X=2.49 $Y=0.355 $X2=0
+ $Y2=0
cc_244 N_A_116_21#_c_158_n N_VGND_c_1413_n 0.0129442f $X=0.655 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_116_21#_c_171_p N_VGND_c_1413_n 0.00486519f $X=1.23 $Y=0.78 $X2=0
+ $Y2=0
cc_246 N_A_116_21#_c_205_p N_VGND_c_1413_n 0.00119066f $X=1 $Y=0.78 $X2=0 $Y2=0
cc_247 N_A_116_21#_c_162_n N_VGND_c_1413_n 0.00844855f $X=1.45 $Y=0.34 $X2=0
+ $Y2=0
cc_248 N_A_116_21#_c_163_n N_VGND_c_1413_n 0.0529876f $X=2.49 $Y=0.355 $X2=0
+ $Y2=0
cc_249 N_C_c_262_n N_A_276_93#_c_324_n 0.0495097f $X=2.45 $Y=1.55 $X2=0 $Y2=0
cc_250 N_C_c_265_n N_A_276_93#_c_324_n 0.001133f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_251 N_C_c_262_n N_A_276_93#_c_325_n 3.1776e-19 $X=2.45 $Y=1.55 $X2=0 $Y2=0
cc_252 N_C_c_263_n N_A_276_93#_c_325_n 0.0194799f $X=2.515 $Y=0.985 $X2=0 $Y2=0
cc_253 N_C_M1001_g N_A_276_93#_c_340_n 0.0115705f $X=1.33 $Y=1.805 $X2=0 $Y2=0
cc_254 N_C_c_261_n N_A_276_93#_c_340_n 0.00616727f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_255 N_C_c_260_n N_A_276_93#_c_326_n 0.00440154f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_256 N_C_M1001_g N_A_276_93#_c_326_n 0.00204947f $X=1.33 $Y=1.805 $X2=0 $Y2=0
cc_257 N_C_c_261_n N_A_276_93#_c_326_n 0.024119f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_258 N_C_c_262_n N_A_276_93#_c_326_n 0.00495404f $X=2.45 $Y=1.55 $X2=0 $Y2=0
cc_259 N_C_c_263_n N_A_276_93#_c_326_n 0.00292894f $X=2.515 $Y=0.985 $X2=0 $Y2=0
cc_260 N_C_c_264_n N_A_276_93#_c_326_n 0.00205064f $X=1.33 $Y=1.202 $X2=0 $Y2=0
cc_261 N_C_c_265_n N_A_276_93#_c_326_n 0.0250009f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_262 N_C_c_261_n N_A_276_93#_c_330_n 0.0145971f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_263 N_C_c_262_n N_A_276_93#_c_330_n 0.0166507f $X=2.45 $Y=1.55 $X2=0 $Y2=0
cc_264 N_C_c_265_n N_A_276_93#_c_330_n 0.0433481f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_265 N_C_c_262_n N_A_276_93#_c_331_n 0.00411747f $X=2.45 $Y=1.55 $X2=0 $Y2=0
cc_266 N_C_c_262_n N_A_276_93#_c_327_n 0.00100184f $X=2.45 $Y=1.55 $X2=0 $Y2=0
cc_267 N_C_c_265_n N_A_276_93#_c_327_n 0.0291268f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_268 N_C_c_260_n N_X_c_883_n 6.32235e-19 $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_269 N_C_M1001_g X 8.72575e-19 $X=1.33 $Y=1.805 $X2=0 $Y2=0
cc_270 N_C_M1001_g N_VPWR_c_908_n 0.00220316f $X=1.33 $Y=1.805 $X2=0 $Y2=0
cc_271 N_C_M1001_g N_VPWR_c_909_n 0.00514356f $X=1.33 $Y=1.805 $X2=0 $Y2=0
cc_272 N_C_c_262_n N_VPWR_c_909_n 0.00427564f $X=2.45 $Y=1.55 $X2=0 $Y2=0
cc_273 N_C_M1001_g N_VPWR_c_907_n 0.00682402f $X=1.33 $Y=1.805 $X2=0 $Y2=0
cc_274 N_C_c_262_n N_VPWR_c_907_n 0.00728509f $X=2.45 $Y=1.55 $X2=0 $Y2=0
cc_275 N_C_M1001_g N_A_406_325#_c_1006_n 9.28125e-19 $X=1.33 $Y=1.805 $X2=0
+ $Y2=0
cc_276 N_C_c_262_n N_A_406_325#_c_1006_n 0.0104309f $X=2.45 $Y=1.55 $X2=0 $Y2=0
cc_277 N_C_c_261_n N_A_424_49#_c_1151_n 0.00625753f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_278 N_C_c_263_n N_A_424_49#_c_1151_n 0.0094194f $X=2.515 $Y=0.985 $X2=0 $Y2=0
cc_279 N_C_c_265_n N_A_424_49#_c_1151_n 0.0382257f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_280 N_C_c_263_n N_A_424_49#_c_1175_n 7.51336e-19 $X=2.515 $Y=0.985 $X2=0
+ $Y2=0
cc_281 N_C_c_260_n N_VGND_c_1404_n 0.00114904f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_282 N_C_c_260_n N_VGND_c_1409_n 7.72982e-19 $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_283 N_C_c_263_n N_VGND_c_1409_n 0.00357877f $X=2.515 $Y=0.985 $X2=0 $Y2=0
cc_284 N_C_c_263_n N_VGND_c_1413_n 0.00706369f $X=2.515 $Y=0.985 $X2=0 $Y2=0
cc_285 N_A_276_93#_c_324_n N_VPWR_c_909_n 0.00455111f $X=3.03 $Y=1.55 $X2=0
+ $Y2=0
cc_286 N_A_276_93#_c_324_n N_VPWR_c_907_n 0.00760152f $X=3.03 $Y=1.55 $X2=0
+ $Y2=0
cc_287 N_A_276_93#_c_330_n N_A_406_325#_M1005_s 0.00366147f $X=2.815 $Y=1.62
+ $X2=0 $Y2=0
cc_288 N_A_276_93#_c_324_n N_A_406_325#_c_1006_n 0.0173326f $X=3.03 $Y=1.55
+ $X2=0 $Y2=0
cc_289 N_A_276_93#_c_330_n N_A_406_325#_c_1006_n 0.0559645f $X=2.815 $Y=1.62
+ $X2=0 $Y2=0
cc_290 N_A_276_93#_c_327_n N_A_406_325#_c_1006_n 0.00386917f $X=3.005 $Y=1.16
+ $X2=0 $Y2=0
cc_291 N_A_276_93#_c_324_n N_A_406_325#_c_1026_n 0.00748858f $X=3.03 $Y=1.55
+ $X2=0 $Y2=0
cc_292 N_A_276_93#_c_330_n N_A_406_325#_c_1026_n 6.13389e-19 $X=2.815 $Y=1.62
+ $X2=0 $Y2=0
cc_293 N_A_276_93#_c_324_n N_A_406_325#_c_1004_n 9.67237e-19 $X=3.03 $Y=1.55
+ $X2=0 $Y2=0
cc_294 N_A_276_93#_c_325_n N_A_406_325#_c_1004_n 0.0136697f $X=3.115 $Y=0.995
+ $X2=0 $Y2=0
cc_295 N_A_276_93#_c_331_n N_A_406_325#_c_1004_n 0.00166649f $X=2.9 $Y=1.535
+ $X2=0 $Y2=0
cc_296 N_A_276_93#_c_327_n N_A_406_325#_c_1004_n 0.015773f $X=3.005 $Y=1.16
+ $X2=0 $Y2=0
cc_297 N_A_276_93#_c_330_n N_A_406_325#_c_1012_n 4.56942e-19 $X=2.815 $Y=1.62
+ $X2=0 $Y2=0
cc_298 N_A_276_93#_c_331_n N_A_406_325#_c_1012_n 6.00479e-19 $X=2.9 $Y=1.535
+ $X2=0 $Y2=0
cc_299 N_A_276_93#_c_324_n N_A_406_325#_c_1014_n 0.00700676f $X=3.03 $Y=1.55
+ $X2=0 $Y2=0
cc_300 N_A_276_93#_c_330_n N_A_406_325#_c_1014_n 0.0109044f $X=2.815 $Y=1.62
+ $X2=0 $Y2=0
cc_301 N_A_276_93#_c_331_n N_A_406_325#_c_1014_n 0.00528578f $X=2.9 $Y=1.535
+ $X2=0 $Y2=0
cc_302 N_A_276_93#_c_324_n N_A_424_49#_c_1151_n 0.0041059f $X=3.03 $Y=1.55 $X2=0
+ $Y2=0
cc_303 N_A_276_93#_c_325_n N_A_424_49#_c_1151_n 0.0121256f $X=3.115 $Y=0.995
+ $X2=0 $Y2=0
cc_304 N_A_276_93#_c_326_n N_A_424_49#_c_1151_n 0.00977033f $X=1.705 $Y=0.76
+ $X2=0 $Y2=0
cc_305 N_A_276_93#_c_327_n N_A_424_49#_c_1151_n 0.0224608f $X=3.005 $Y=1.16
+ $X2=0 $Y2=0
cc_306 N_A_276_93#_c_325_n N_A_424_49#_c_1175_n 0.00969442f $X=3.115 $Y=0.995
+ $X2=0 $Y2=0
cc_307 N_A_276_93#_c_325_n N_A_424_49#_c_1176_n 0.00814783f $X=3.115 $Y=0.995
+ $X2=0 $Y2=0
cc_308 N_A_276_93#_c_324_n N_A_424_49#_c_1158_n 0.00452598f $X=3.03 $Y=1.55
+ $X2=0 $Y2=0
cc_309 N_A_276_93#_c_324_n N_A_424_49#_c_1160_n 7.6183e-19 $X=3.03 $Y=1.55 $X2=0
+ $Y2=0
cc_310 N_A_276_93#_c_325_n N_A_424_49#_c_1153_n 0.00103799f $X=3.115 $Y=0.995
+ $X2=0 $Y2=0
cc_311 N_A_276_93#_c_324_n N_A_424_49#_c_1168_n 0.00354471f $X=3.03 $Y=1.55
+ $X2=0 $Y2=0
cc_312 N_A_276_93#_c_325_n N_VGND_c_1409_n 0.00367048f $X=3.115 $Y=0.995 $X2=0
+ $Y2=0
cc_313 N_A_276_93#_c_325_n N_VGND_c_1413_n 0.00715174f $X=3.115 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_A_875_297#_c_418_n N_B_c_588_n 0.00851867f $X=4.675 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_315 N_A_875_297#_c_412_n N_B_c_588_n 8.21886e-19 $X=4.735 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_316 N_A_875_297#_c_422_p N_B_M1003_g 0.00371022f $X=4.765 $Y=0.85 $X2=0 $Y2=0
cc_317 N_A_875_297#_c_412_n N_B_M1003_g 0.0174461f $X=4.735 $Y=0.72 $X2=0 $Y2=0
cc_318 N_A_875_297#_c_404_n N_B_c_581_n 0.00502253f $X=5.955 $Y=0.85 $X2=0 $Y2=0
cc_319 N_A_875_297#_c_412_n N_B_c_581_n 0.0123135f $X=4.735 $Y=0.72 $X2=0 $Y2=0
cc_320 N_A_875_297#_c_418_n N_B_c_582_n 0.00731407f $X=4.675 $Y=1.58 $X2=0 $Y2=0
cc_321 N_A_875_297#_c_412_n N_B_c_582_n 0.00954146f $X=4.735 $Y=0.72 $X2=0 $Y2=0
cc_322 N_A_875_297#_c_413_n N_B_M1011_g 0.0117988f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A_875_297#_M1008_g N_B_M1004_g 0.0101671f $X=6.315 $Y=0.455 $X2=0 $Y2=0
cc_324 N_A_875_297#_c_401_n N_B_M1004_g 0.0212291f $X=6.19 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_875_297#_c_403_n N_B_M1004_g 0.00190447f $X=6.077 $Y=0.995 $X2=0
+ $Y2=0
cc_326 N_A_875_297#_c_404_n N_B_M1004_g 0.00156951f $X=5.955 $Y=0.85 $X2=0 $Y2=0
cc_327 N_A_875_297#_c_406_n N_B_M1004_g 6.73467e-19 $X=6.245 $Y=0.85 $X2=0 $Y2=0
cc_328 N_A_875_297#_c_407_n N_B_M1004_g 0.00123519f $X=6.1 $Y=0.85 $X2=0 $Y2=0
cc_329 N_A_875_297#_c_413_n N_B_c_591_n 0.0105804f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_330 N_A_875_297#_c_415_n N_B_c_591_n 0.00616735f $X=7.78 $Y=1.57 $X2=0 $Y2=0
cc_331 N_A_875_297#_c_400_n N_B_c_593_n 0.00407979f $X=7.78 $Y=1.47 $X2=0 $Y2=0
cc_332 N_A_875_297#_c_415_n N_B_c_594_n 0.00407979f $X=7.78 $Y=1.57 $X2=0 $Y2=0
cc_333 N_A_875_297#_c_415_n N_B_M1012_g 0.0242934f $X=7.78 $Y=1.57 $X2=0 $Y2=0
cc_334 N_A_875_297#_c_402_n N_B_c_584_n 0.00179713f $X=6.29 $Y=1.202 $X2=0 $Y2=0
cc_335 N_A_875_297#_c_400_n N_B_c_585_n 9.96285e-19 $X=7.78 $Y=1.47 $X2=0 $Y2=0
cc_336 N_A_875_297#_c_405_n N_B_c_585_n 0.00735944f $X=7.435 $Y=0.85 $X2=0 $Y2=0
cc_337 N_A_875_297#_c_409_n N_B_c_585_n 0.021521f $X=7.58 $Y=0.85 $X2=0 $Y2=0
cc_338 N_A_875_297#_c_410_n N_B_c_585_n 2.70696e-19 $X=7.7 $Y=1.11 $X2=0 $Y2=0
cc_339 N_A_875_297#_c_400_n N_B_c_586_n 0.00187722f $X=7.78 $Y=1.47 $X2=0 $Y2=0
cc_340 N_A_875_297#_c_402_n N_B_c_586_n 0.00774829f $X=6.29 $Y=1.202 $X2=0 $Y2=0
cc_341 N_A_875_297#_c_405_n N_B_c_586_n 0.00133312f $X=7.435 $Y=0.85 $X2=0 $Y2=0
cc_342 N_A_875_297#_c_409_n N_B_c_586_n 0.00172718f $X=7.58 $Y=0.85 $X2=0 $Y2=0
cc_343 N_A_875_297#_c_410_n N_B_c_586_n 0.0173414f $X=7.7 $Y=1.11 $X2=0 $Y2=0
cc_344 N_A_875_297#_c_400_n B 0.00134318f $X=7.78 $Y=1.47 $X2=0 $Y2=0
cc_345 N_A_875_297#_c_415_n B 0.00796231f $X=7.78 $Y=1.57 $X2=0 $Y2=0
cc_346 N_A_875_297#_c_405_n B 0.004363f $X=7.435 $Y=0.85 $X2=0 $Y2=0
cc_347 N_A_875_297#_c_408_n B 0.00246368f $X=7.58 $Y=0.85 $X2=0 $Y2=0
cc_348 N_A_875_297#_c_409_n B 0.0189884f $X=7.58 $Y=0.85 $X2=0 $Y2=0
cc_349 N_A_875_297#_c_410_n B 8.41241e-19 $X=7.7 $Y=1.11 $X2=0 $Y2=0
cc_350 N_A_875_297#_M1008_g N_B_c_587_n 0.00774829f $X=6.315 $Y=0.455 $X2=0
+ $Y2=0
cc_351 N_A_875_297#_c_405_n N_B_c_587_n 0.0073961f $X=7.435 $Y=0.85 $X2=0 $Y2=0
cc_352 N_A_875_297#_c_408_n N_B_c_587_n 0.00141075f $X=7.58 $Y=0.85 $X2=0 $Y2=0
cc_353 N_A_875_297#_c_409_n N_B_c_587_n 0.00206736f $X=7.58 $Y=0.85 $X2=0 $Y2=0
cc_354 N_A_875_297#_c_410_n N_B_c_587_n 0.00135765f $X=7.7 $Y=1.11 $X2=0 $Y2=0
cc_355 N_A_875_297#_c_411_n N_B_c_587_n 0.0136423f $X=7.722 $Y=0.945 $X2=0 $Y2=0
cc_356 N_A_875_297#_c_400_n N_A_c_717_n 0.00765017f $X=7.78 $Y=1.47 $X2=-0.19
+ $Y2=-0.24
cc_357 N_A_875_297#_c_415_n N_A_c_717_n 0.031553f $X=7.78 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_358 N_A_875_297#_c_409_n N_A_c_717_n 6.51299e-19 $X=7.58 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_359 N_A_875_297#_c_410_n N_A_c_717_n 0.0202732f $X=7.7 $Y=1.11 $X2=-0.19
+ $Y2=-0.24
cc_360 N_A_875_297#_c_409_n N_A_c_718_n 2.39914e-19 $X=7.58 $Y=0.85 $X2=0 $Y2=0
cc_361 N_A_875_297#_c_411_n N_A_c_718_n 0.0185553f $X=7.722 $Y=0.945 $X2=0 $Y2=0
cc_362 N_A_875_297#_c_409_n A 0.0138459f $X=7.58 $Y=0.85 $X2=0 $Y2=0
cc_363 N_A_875_297#_c_410_n A 0.00288931f $X=7.7 $Y=1.11 $X2=0 $Y2=0
cc_364 N_A_875_297#_c_404_n N_A_991_365#_M1004_s 8.50051e-19 $X=5.955 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_365 N_A_875_297#_c_418_n N_A_991_365#_c_756_n 0.0199218f $X=4.675 $Y=1.58
+ $X2=0 $Y2=0
cc_366 N_A_875_297#_c_404_n N_A_991_365#_c_756_n 0.0123662f $X=5.955 $Y=0.85
+ $X2=0 $Y2=0
cc_367 N_A_875_297#_c_422_p N_A_991_365#_c_756_n 5.85147e-19 $X=4.765 $Y=0.85
+ $X2=0 $Y2=0
cc_368 N_A_875_297#_c_412_n N_A_991_365#_c_756_n 0.0617741f $X=4.735 $Y=0.72
+ $X2=0 $Y2=0
cc_369 N_A_875_297#_c_415_n N_A_991_365#_c_764_n 0.00215422f $X=7.78 $Y=1.57
+ $X2=0 $Y2=0
cc_370 N_A_875_297#_c_408_n N_A_991_365#_c_758_n 0.00537182f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_371 N_A_875_297#_c_409_n N_A_991_365#_c_758_n 0.0052004f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_372 N_A_875_297#_c_411_n N_A_991_365#_c_758_n 0.00186387f $X=7.722 $Y=0.945
+ $X2=0 $Y2=0
cc_373 N_A_875_297#_M1008_g N_A_991_365#_c_776_n 0.00614563f $X=6.315 $Y=0.455
+ $X2=0 $Y2=0
cc_374 N_A_875_297#_c_403_n N_A_991_365#_c_776_n 3.7129e-19 $X=6.077 $Y=0.995
+ $X2=0 $Y2=0
cc_375 N_A_875_297#_c_404_n N_A_991_365#_c_776_n 0.0529545f $X=5.955 $Y=0.85
+ $X2=0 $Y2=0
cc_376 N_A_875_297#_c_405_n N_A_991_365#_c_776_n 0.0955498f $X=7.435 $Y=0.85
+ $X2=0 $Y2=0
cc_377 N_A_875_297#_c_406_n N_A_991_365#_c_776_n 0.0266362f $X=6.245 $Y=0.85
+ $X2=0 $Y2=0
cc_378 N_A_875_297#_c_407_n N_A_991_365#_c_776_n 0.00318096f $X=6.1 $Y=0.85
+ $X2=0 $Y2=0
cc_379 N_A_875_297#_c_408_n N_A_991_365#_c_776_n 0.0266136f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_380 N_A_875_297#_c_409_n N_A_991_365#_c_776_n 0.00475925f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_381 N_A_875_297#_c_411_n N_A_991_365#_c_776_n 0.00868614f $X=7.722 $Y=0.945
+ $X2=0 $Y2=0
cc_382 N_A_875_297#_c_404_n N_A_991_365#_c_760_n 0.0261136f $X=5.955 $Y=0.85
+ $X2=0 $Y2=0
cc_383 N_A_875_297#_c_412_n N_A_991_365#_c_760_n 0.00677952f $X=4.735 $Y=0.72
+ $X2=0 $Y2=0
cc_384 N_A_875_297#_c_404_n N_A_991_365#_c_761_n 0.00110106f $X=5.955 $Y=0.85
+ $X2=0 $Y2=0
cc_385 N_A_875_297#_c_412_n N_A_991_365#_c_761_n 0.0118823f $X=4.735 $Y=0.72
+ $X2=0 $Y2=0
cc_386 N_A_875_297#_c_411_n N_A_991_365#_c_789_n 0.00156339f $X=7.722 $Y=0.945
+ $X2=0 $Y2=0
cc_387 N_A_875_297#_c_411_n N_A_991_365#_c_790_n 0.00805147f $X=7.722 $Y=0.945
+ $X2=0 $Y2=0
cc_388 N_A_875_297#_M1006_d N_VPWR_c_907_n 0.00359518f $X=4.375 $Y=1.485 $X2=0
+ $Y2=0
cc_389 N_A_875_297#_c_415_n N_VPWR_c_907_n 0.00650675f $X=7.78 $Y=1.57 $X2=0
+ $Y2=0
cc_390 N_A_875_297#_c_415_n N_VPWR_c_916_n 0.00434439f $X=7.78 $Y=1.57 $X2=0
+ $Y2=0
cc_391 N_A_875_297#_c_415_n N_VPWR_c_917_n 0.00134203f $X=7.78 $Y=1.57 $X2=0
+ $Y2=0
cc_392 N_A_875_297#_c_405_n N_A_406_325#_M1009_d 0.00140408f $X=7.435 $Y=0.85
+ $X2=0 $Y2=0
cc_393 N_A_875_297#_c_408_n N_A_406_325#_M1009_d 0.00214439f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_394 N_A_875_297#_c_409_n N_A_406_325#_M1009_d 0.0050343f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_395 N_A_875_297#_c_401_n N_A_406_325#_c_1008_n 0.00894291f $X=6.19 $Y=1.16
+ $X2=0 $Y2=0
cc_396 N_A_875_297#_c_403_n N_A_406_325#_c_1008_n 0.0270839f $X=6.077 $Y=0.995
+ $X2=0 $Y2=0
cc_397 N_A_875_297#_c_404_n N_A_406_325#_c_1008_n 5.63647e-19 $X=5.955 $Y=0.85
+ $X2=0 $Y2=0
cc_398 N_A_875_297#_c_413_n N_A_406_325#_c_1043_n 0.00385601f $X=6.29 $Y=1.41
+ $X2=0 $Y2=0
cc_399 N_A_875_297#_c_413_n N_A_406_325#_c_1009_n 0.0175866f $X=6.29 $Y=1.41
+ $X2=0 $Y2=0
cc_400 N_A_875_297#_c_401_n N_A_406_325#_c_1009_n 7.42472e-19 $X=6.19 $Y=1.16
+ $X2=0 $Y2=0
cc_401 N_A_875_297#_c_402_n N_A_406_325#_c_1009_n 9.0109e-19 $X=6.29 $Y=1.202
+ $X2=0 $Y2=0
cc_402 N_A_875_297#_c_403_n N_A_406_325#_c_1009_n 0.00152864f $X=6.077 $Y=0.995
+ $X2=0 $Y2=0
cc_403 N_A_875_297#_c_405_n N_A_406_325#_c_1009_n 0.00419686f $X=7.435 $Y=0.85
+ $X2=0 $Y2=0
cc_404 N_A_875_297#_c_406_n N_A_406_325#_c_1009_n 6.55203e-19 $X=6.245 $Y=0.85
+ $X2=0 $Y2=0
cc_405 N_A_875_297#_c_413_n N_A_406_325#_c_1005_n 0.00139259f $X=6.29 $Y=1.41
+ $X2=0 $Y2=0
cc_406 N_A_875_297#_M1008_g N_A_406_325#_c_1005_n 0.0164123f $X=6.315 $Y=0.455
+ $X2=0 $Y2=0
cc_407 N_A_875_297#_c_403_n N_A_406_325#_c_1005_n 0.0173003f $X=6.077 $Y=0.995
+ $X2=0 $Y2=0
cc_408 N_A_875_297#_c_405_n N_A_406_325#_c_1005_n 0.0173494f $X=7.435 $Y=0.85
+ $X2=0 $Y2=0
cc_409 N_A_875_297#_c_406_n N_A_406_325#_c_1005_n 0.00232583f $X=6.245 $Y=0.85
+ $X2=0 $Y2=0
cc_410 N_A_875_297#_c_407_n N_A_406_325#_c_1005_n 0.0185429f $X=6.1 $Y=0.85
+ $X2=0 $Y2=0
cc_411 N_A_875_297#_c_405_n N_A_406_325#_c_1056_n 0.00166303f $X=7.435 $Y=0.85
+ $X2=0 $Y2=0
cc_412 N_A_875_297#_c_408_n N_A_406_325#_c_1057_n 3.55136e-19 $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_413 N_A_875_297#_c_409_n N_A_406_325#_c_1057_n 0.00528249f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_414 N_A_875_297#_c_411_n N_A_406_325#_c_1057_n 0.00335197f $X=7.722 $Y=0.945
+ $X2=0 $Y2=0
cc_415 N_A_875_297#_c_418_n N_A_406_325#_c_1011_n 0.0271848f $X=4.675 $Y=1.58
+ $X2=0 $Y2=0
cc_416 N_A_875_297#_c_403_n N_A_406_325#_c_1011_n 8.37577e-19 $X=6.077 $Y=0.995
+ $X2=0 $Y2=0
cc_417 N_A_875_297#_c_404_n N_A_406_325#_c_1011_n 0.0525503f $X=5.955 $Y=0.85
+ $X2=0 $Y2=0
cc_418 N_A_875_297#_c_422_p N_A_406_325#_c_1011_n 0.0124517f $X=4.765 $Y=0.85
+ $X2=0 $Y2=0
cc_419 N_A_875_297#_c_412_n N_A_406_325#_c_1011_n 0.00234408f $X=4.735 $Y=0.72
+ $X2=0 $Y2=0
cc_420 N_A_875_297#_c_413_n N_A_406_325#_c_1013_n 0.00348597f $X=6.29 $Y=1.41
+ $X2=0 $Y2=0
cc_421 N_A_875_297#_c_401_n N_A_406_325#_c_1013_n 0.00431105f $X=6.19 $Y=1.16
+ $X2=0 $Y2=0
cc_422 N_A_875_297#_c_402_n N_A_406_325#_c_1013_n 2.0806e-19 $X=6.29 $Y=1.202
+ $X2=0 $Y2=0
cc_423 N_A_875_297#_c_403_n N_A_406_325#_c_1013_n 0.00243787f $X=6.077 $Y=0.995
+ $X2=0 $Y2=0
cc_424 N_A_875_297#_c_406_n N_A_406_325#_c_1013_n 0.0154521f $X=6.245 $Y=0.85
+ $X2=0 $Y2=0
cc_425 N_A_875_297#_c_404_n N_A_424_49#_M1004_d 0.00139415f $X=5.955 $Y=0.85
+ $X2=0 $Y2=0
cc_426 N_A_875_297#_c_406_n N_A_424_49#_M1004_d 5.07779e-19 $X=6.245 $Y=0.85
+ $X2=0 $Y2=0
cc_427 N_A_875_297#_c_407_n N_A_424_49#_M1004_d 0.00662486f $X=6.1 $Y=0.85 $X2=0
+ $Y2=0
cc_428 N_A_875_297#_c_422_p N_A_424_49#_c_1153_n 0.00233211f $X=4.765 $Y=0.85
+ $X2=0 $Y2=0
cc_429 N_A_875_297#_c_412_n N_A_424_49#_c_1153_n 0.00359007f $X=4.735 $Y=0.72
+ $X2=0 $Y2=0
cc_430 N_A_875_297#_c_418_n N_A_424_49#_c_1154_n 0.0144112f $X=4.675 $Y=1.58
+ $X2=0 $Y2=0
cc_431 N_A_875_297#_c_412_n N_A_424_49#_c_1154_n 0.00935491f $X=4.735 $Y=0.72
+ $X2=0 $Y2=0
cc_432 N_A_875_297#_M1006_d N_A_424_49#_c_1162_n 0.0074794f $X=4.375 $Y=1.485
+ $X2=0 $Y2=0
cc_433 N_A_875_297#_c_418_n N_A_424_49#_c_1162_n 0.0314935f $X=4.675 $Y=1.58
+ $X2=0 $Y2=0
cc_434 N_A_875_297#_M1006_d N_A_424_49#_c_1163_n 0.00302314f $X=4.375 $Y=1.485
+ $X2=0 $Y2=0
cc_435 N_A_875_297#_M1006_d N_A_424_49#_c_1165_n 0.00298868f $X=4.375 $Y=1.485
+ $X2=0 $Y2=0
cc_436 N_A_875_297#_c_413_n N_A_424_49#_c_1155_n 0.00130504f $X=6.29 $Y=1.41
+ $X2=0 $Y2=0
cc_437 N_A_875_297#_c_401_n N_A_424_49#_c_1155_n 6.50075e-19 $X=6.19 $Y=1.16
+ $X2=0 $Y2=0
cc_438 N_A_875_297#_c_402_n N_A_424_49#_c_1155_n 3.92684e-19 $X=6.29 $Y=1.202
+ $X2=0 $Y2=0
cc_439 N_A_875_297#_c_403_n N_A_424_49#_c_1155_n 0.0156137f $X=6.077 $Y=0.995
+ $X2=0 $Y2=0
cc_440 N_A_875_297#_c_404_n N_A_424_49#_c_1155_n 0.00605333f $X=5.955 $Y=0.85
+ $X2=0 $Y2=0
cc_441 N_A_875_297#_c_406_n N_A_424_49#_c_1155_n 0.00104191f $X=6.245 $Y=0.85
+ $X2=0 $Y2=0
cc_442 N_A_875_297#_c_407_n N_A_424_49#_c_1155_n 0.00261896f $X=6.1 $Y=0.85
+ $X2=0 $Y2=0
cc_443 N_A_875_297#_c_413_n N_A_424_49#_c_1167_n 0.00258134f $X=6.29 $Y=1.41
+ $X2=0 $Y2=0
cc_444 N_A_875_297#_c_415_n N_A_424_49#_c_1167_n 0.00822576f $X=7.78 $Y=1.57
+ $X2=0 $Y2=0
cc_445 N_A_875_297#_M1008_g N_A_424_49#_c_1212_n 0.0022242f $X=6.315 $Y=0.455
+ $X2=0 $Y2=0
cc_446 N_A_875_297#_c_407_n N_A_424_49#_c_1212_n 0.00181204f $X=6.1 $Y=0.85
+ $X2=0 $Y2=0
cc_447 N_A_875_297#_c_412_n N_A_424_49#_c_1156_n 0.00622512f $X=4.735 $Y=0.72
+ $X2=0 $Y2=0
cc_448 N_A_875_297#_c_401_n N_A_424_49#_c_1157_n 2.22283e-19 $X=6.19 $Y=1.16
+ $X2=0 $Y2=0
cc_449 N_A_875_297#_c_403_n N_A_424_49#_c_1157_n 0.00265833f $X=6.077 $Y=0.995
+ $X2=0 $Y2=0
cc_450 N_A_875_297#_c_404_n N_A_424_49#_c_1157_n 0.0174471f $X=5.955 $Y=0.85
+ $X2=0 $Y2=0
cc_451 N_A_875_297#_c_406_n N_A_424_49#_c_1157_n 0.00133974f $X=6.245 $Y=0.85
+ $X2=0 $Y2=0
cc_452 N_A_875_297#_c_407_n N_A_424_49#_c_1157_n 0.0142042f $X=6.1 $Y=0.85 $X2=0
+ $Y2=0
cc_453 N_A_875_297#_c_405_n N_A_1276_297#_M1008_d 0.00166227f $X=7.435 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_454 N_A_875_297#_c_413_n N_A_1276_297#_c_1338_n 0.00686704f $X=6.29 $Y=1.41
+ $X2=0 $Y2=0
cc_455 N_A_875_297#_c_405_n N_A_1276_297#_c_1338_n 0.0181022f $X=7.435 $Y=0.85
+ $X2=0 $Y2=0
cc_456 N_A_875_297#_c_408_n N_A_1276_297#_c_1338_n 0.0020738f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_457 N_A_875_297#_c_409_n N_A_1276_297#_c_1338_n 0.00517339f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_458 N_A_875_297#_c_413_n N_A_1276_297#_c_1350_n 0.00431165f $X=6.29 $Y=1.41
+ $X2=0 $Y2=0
cc_459 N_A_875_297#_c_415_n N_A_1276_297#_c_1351_n 0.0164032f $X=7.78 $Y=1.57
+ $X2=0 $Y2=0
cc_460 N_A_875_297#_c_409_n N_A_1276_297#_c_1351_n 0.00161448f $X=7.58 $Y=0.85
+ $X2=0 $Y2=0
cc_461 N_A_875_297#_c_422_p N_VGND_c_1405_n 0.00369072f $X=4.765 $Y=0.85 $X2=0
+ $Y2=0
cc_462 N_A_875_297#_c_412_n N_VGND_c_1405_n 0.0242508f $X=4.735 $Y=0.72 $X2=0
+ $Y2=0
cc_463 N_A_875_297#_M1008_g N_VGND_c_1411_n 0.00575161f $X=6.315 $Y=0.455 $X2=0
+ $Y2=0
cc_464 N_A_875_297#_c_407_n N_VGND_c_1411_n 0.00348958f $X=6.1 $Y=0.85 $X2=0
+ $Y2=0
cc_465 N_A_875_297#_c_409_n N_VGND_c_1411_n 0.00102193f $X=7.58 $Y=0.85 $X2=0
+ $Y2=0
cc_466 N_A_875_297#_c_411_n N_VGND_c_1411_n 0.00585385f $X=7.722 $Y=0.945 $X2=0
+ $Y2=0
cc_467 N_A_875_297#_c_412_n N_VGND_c_1411_n 0.0088551f $X=4.735 $Y=0.72 $X2=0
+ $Y2=0
cc_468 N_A_875_297#_M1003_d N_VGND_c_1413_n 0.00198683f $X=4.6 $Y=0.235 $X2=0
+ $Y2=0
cc_469 N_A_875_297#_M1008_g N_VGND_c_1413_n 0.00669445f $X=6.315 $Y=0.455 $X2=0
+ $Y2=0
cc_470 N_A_875_297#_c_404_n N_VGND_c_1413_n 0.0112971f $X=5.955 $Y=0.85 $X2=0
+ $Y2=0
cc_471 N_A_875_297#_c_422_p N_VGND_c_1413_n 0.0147993f $X=4.765 $Y=0.85 $X2=0
+ $Y2=0
cc_472 N_A_875_297#_c_411_n N_VGND_c_1413_n 0.00635691f $X=7.722 $Y=0.945 $X2=0
+ $Y2=0
cc_473 N_A_875_297#_c_412_n N_VGND_c_1413_n 0.00448337f $X=4.735 $Y=0.72 $X2=0
+ $Y2=0
cc_474 N_B_c_588_n N_A_991_365#_c_756_n 0.00363086f $X=4.285 $Y=1.41 $X2=0 $Y2=0
cc_475 N_B_M1003_g N_A_991_365#_c_756_n 0.00120086f $X=4.525 $Y=0.56 $X2=0 $Y2=0
cc_476 N_B_c_581_n N_A_991_365#_c_756_n 0.0145436f $X=5.38 $Y=1.16 $X2=0 $Y2=0
cc_477 N_B_M1011_g N_A_991_365#_c_756_n 0.00419529f $X=5.48 $Y=1.905 $X2=0 $Y2=0
cc_478 N_B_M1004_g N_A_991_365#_c_756_n 0.00351927f $X=5.505 $Y=0.565 $X2=0
+ $Y2=0
cc_479 N_B_c_584_n N_A_991_365#_c_756_n 0.00110014f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_480 B N_A_991_365#_c_764_n 0.015034f $X=7.495 $Y=1.5 $X2=0 $Y2=0
cc_481 N_B_M1004_g N_A_991_365#_c_776_n 0.00201366f $X=5.505 $Y=0.565 $X2=0
+ $Y2=0
cc_482 N_B_c_587_n N_A_991_365#_c_776_n 0.0032563f $X=7.195 $Y=0.995 $X2=0 $Y2=0
cc_483 N_B_M1003_g N_A_991_365#_c_760_n 4.1997e-19 $X=4.525 $Y=0.56 $X2=0 $Y2=0
cc_484 N_B_M1004_g N_A_991_365#_c_760_n 9.1979e-19 $X=5.505 $Y=0.565 $X2=0 $Y2=0
cc_485 N_B_M1003_g N_A_991_365#_c_761_n 0.00489085f $X=4.525 $Y=0.56 $X2=0 $Y2=0
cc_486 N_B_c_581_n N_A_991_365#_c_761_n 0.00313752f $X=5.38 $Y=1.16 $X2=0 $Y2=0
cc_487 N_B_c_588_n N_VPWR_c_910_n 0.0113699f $X=4.285 $Y=1.41 $X2=0 $Y2=0
cc_488 N_B_c_588_n N_VPWR_c_907_n 0.00656627f $X=4.285 $Y=1.41 $X2=0 $Y2=0
cc_489 N_B_c_591_n N_VPWR_c_907_n 0.0413158f $X=7.115 $Y=2.54 $X2=0 $Y2=0
cc_490 N_B_c_592_n N_VPWR_c_907_n 0.00712081f $X=5.58 $Y=2.54 $X2=0 $Y2=0
cc_491 N_B_c_588_n N_VPWR_c_916_n 0.00455828f $X=4.285 $Y=1.41 $X2=0 $Y2=0
cc_492 N_B_c_592_n N_VPWR_c_916_n 0.0408109f $X=5.58 $Y=2.54 $X2=0 $Y2=0
cc_493 N_B_c_582_n N_A_406_325#_c_1004_n 4.45781e-19 $X=4.6 $Y=1.16 $X2=0 $Y2=0
cc_494 N_B_M1011_g N_A_406_325#_c_1008_n 0.00146463f $X=5.48 $Y=1.905 $X2=0
+ $Y2=0
cc_495 N_B_M1011_g N_A_406_325#_c_1043_n 0.0044998f $X=5.48 $Y=1.905 $X2=0 $Y2=0
cc_496 N_B_c_587_n N_A_406_325#_c_1005_n 0.0026019f $X=7.195 $Y=0.995 $X2=0
+ $Y2=0
cc_497 N_B_c_585_n N_A_406_325#_c_1056_n 0.00294871f $X=7.17 $Y=1.16 $X2=0 $Y2=0
cc_498 N_B_c_586_n N_A_406_325#_c_1056_n 4.30216e-19 $X=7.17 $Y=1.16 $X2=0 $Y2=0
cc_499 N_B_c_587_n N_A_406_325#_c_1056_n 0.00498906f $X=7.195 $Y=0.995 $X2=0
+ $Y2=0
cc_500 N_B_c_586_n N_A_406_325#_c_1057_n 0.00110831f $X=7.17 $Y=1.16 $X2=0 $Y2=0
cc_501 N_B_c_587_n N_A_406_325#_c_1078_n 0.00521263f $X=7.195 $Y=0.995 $X2=0
+ $Y2=0
cc_502 N_B_c_588_n N_A_406_325#_c_1011_n 0.00484975f $X=4.285 $Y=1.41 $X2=0
+ $Y2=0
cc_503 N_B_c_581_n N_A_406_325#_c_1011_n 0.00478884f $X=5.38 $Y=1.16 $X2=0 $Y2=0
cc_504 N_B_c_582_n N_A_406_325#_c_1011_n 2.58451e-19 $X=4.6 $Y=1.16 $X2=0 $Y2=0
cc_505 N_B_M1011_g N_A_406_325#_c_1011_n 0.00508939f $X=5.48 $Y=1.905 $X2=0
+ $Y2=0
cc_506 N_B_c_584_n N_A_406_325#_c_1011_n 2.29578e-19 $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_507 N_B_M1011_g N_A_406_325#_c_1013_n 4.47596e-19 $X=5.48 $Y=1.905 $X2=0
+ $Y2=0
cc_508 B N_A_424_49#_M1012_d 0.00323521f $X=7.495 $Y=1.5 $X2=0 $Y2=0
cc_509 N_B_c_588_n N_A_424_49#_c_1158_n 0.00287893f $X=4.285 $Y=1.41 $X2=0 $Y2=0
cc_510 N_B_M1003_g N_A_424_49#_c_1153_n 0.00319704f $X=4.525 $Y=0.56 $X2=0 $Y2=0
cc_511 N_B_c_588_n N_A_424_49#_c_1154_n 0.0127864f $X=4.285 $Y=1.41 $X2=0 $Y2=0
cc_512 N_B_c_582_n N_A_424_49#_c_1154_n 0.00534802f $X=4.6 $Y=1.16 $X2=0 $Y2=0
cc_513 N_B_c_588_n N_A_424_49#_c_1162_n 0.0174362f $X=4.285 $Y=1.41 $X2=0 $Y2=0
cc_514 N_B_c_588_n N_A_424_49#_c_1163_n 0.00608631f $X=4.285 $Y=1.41 $X2=0 $Y2=0
cc_515 N_B_M1011_g N_A_424_49#_c_1163_n 8.91158e-19 $X=5.48 $Y=1.905 $X2=0 $Y2=0
cc_516 N_B_c_588_n N_A_424_49#_c_1165_n 0.00366198f $X=4.285 $Y=1.41 $X2=0 $Y2=0
cc_517 N_B_c_581_n N_A_424_49#_c_1155_n 0.00364094f $X=5.38 $Y=1.16 $X2=0 $Y2=0
cc_518 N_B_M1011_g N_A_424_49#_c_1155_n 0.0315702f $X=5.48 $Y=1.905 $X2=0 $Y2=0
cc_519 N_B_M1004_g N_A_424_49#_c_1155_n 0.00650642f $X=5.505 $Y=0.565 $X2=0
+ $Y2=0
cc_520 N_B_c_584_n N_A_424_49#_c_1155_n 0.0104909f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_521 N_B_M1011_g N_A_424_49#_c_1167_n 0.00851955f $X=5.48 $Y=1.905 $X2=0 $Y2=0
cc_522 N_B_c_591_n N_A_424_49#_c_1167_n 0.0365765f $X=7.115 $Y=2.54 $X2=0 $Y2=0
cc_523 N_B_c_592_n N_A_424_49#_c_1167_n 2.38151e-19 $X=5.58 $Y=2.54 $X2=0 $Y2=0
cc_524 N_B_M1012_g N_A_424_49#_c_1167_n 0.0102069f $X=7.215 $Y=1.965 $X2=0 $Y2=0
cc_525 N_B_M1004_g N_A_424_49#_c_1212_n 5.72667e-19 $X=5.505 $Y=0.565 $X2=0
+ $Y2=0
cc_526 N_B_M1003_g N_A_424_49#_c_1156_n 8.52685e-19 $X=4.525 $Y=0.56 $X2=0 $Y2=0
cc_527 N_B_c_582_n N_A_424_49#_c_1156_n 0.00386142f $X=4.6 $Y=1.16 $X2=0 $Y2=0
cc_528 N_B_M1004_g N_A_424_49#_c_1157_n 0.013823f $X=5.505 $Y=0.565 $X2=0 $Y2=0
cc_529 N_B_M1011_g N_A_424_49#_c_1170_n 0.00703655f $X=5.48 $Y=1.905 $X2=0 $Y2=0
cc_530 N_B_c_592_n N_A_424_49#_c_1170_n 2.51585e-19 $X=5.58 $Y=2.54 $X2=0 $Y2=0
cc_531 N_B_c_593_n N_A_1276_297#_c_1338_n 0.00160527f $X=7.215 $Y=1.47 $X2=0
+ $Y2=0
cc_532 N_B_M1012_g N_A_1276_297#_c_1338_n 0.00614132f $X=7.215 $Y=1.965 $X2=0
+ $Y2=0
cc_533 N_B_c_597_n N_A_1276_297#_c_1338_n 0.0196555f $X=7.195 $Y=1.445 $X2=0
+ $Y2=0
cc_534 N_B_c_585_n N_A_1276_297#_c_1338_n 0.0332296f $X=7.17 $Y=1.16 $X2=0 $Y2=0
cc_535 N_B_c_587_n N_A_1276_297#_c_1338_n 0.0105486f $X=7.195 $Y=0.995 $X2=0
+ $Y2=0
cc_536 N_B_M1012_g N_A_1276_297#_c_1351_n 0.0104919f $X=7.215 $Y=1.965 $X2=0
+ $Y2=0
cc_537 N_B_c_597_n N_A_1276_297#_c_1351_n 0.0115397f $X=7.195 $Y=1.445 $X2=0
+ $Y2=0
cc_538 N_B_c_586_n N_A_1276_297#_c_1351_n 0.00114355f $X=7.17 $Y=1.16 $X2=0
+ $Y2=0
cc_539 B N_A_1276_297#_c_1351_n 0.0189751f $X=7.495 $Y=1.5 $X2=0 $Y2=0
cc_540 N_B_M1003_g N_VGND_c_1405_n 0.0190364f $X=4.525 $Y=0.56 $X2=0 $Y2=0
cc_541 N_B_c_582_n N_VGND_c_1405_n 0.00518895f $X=4.6 $Y=1.16 $X2=0 $Y2=0
cc_542 N_B_M1003_g N_VGND_c_1411_n 0.00494995f $X=4.525 $Y=0.56 $X2=0 $Y2=0
cc_543 N_B_M1004_g N_VGND_c_1411_n 0.00427876f $X=5.505 $Y=0.565 $X2=0 $Y2=0
cc_544 N_B_c_587_n N_VGND_c_1411_n 0.00357877f $X=7.195 $Y=0.995 $X2=0 $Y2=0
cc_545 N_B_M1003_g N_VGND_c_1413_n 0.00933567f $X=4.525 $Y=0.56 $X2=0 $Y2=0
cc_546 N_B_M1004_g N_VGND_c_1413_n 0.00718941f $X=5.505 $Y=0.565 $X2=0 $Y2=0
cc_547 N_B_c_587_n N_VGND_c_1413_n 0.00612424f $X=7.195 $Y=0.995 $X2=0 $Y2=0
cc_548 N_A_c_717_n N_A_991_365#_c_754_n 0.0284366f $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_549 A N_A_991_365#_c_754_n 0.00118453f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_550 N_A_c_718_n N_A_991_365#_c_755_n 0.0129172f $X=8.36 $Y=0.995 $X2=0 $Y2=0
cc_551 N_A_c_717_n N_A_991_365#_c_764_n 0.015957f $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_552 A N_A_991_365#_c_764_n 0.0473094f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_553 N_A_c_717_n N_A_991_365#_c_757_n 5.76324e-19 $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_554 N_A_c_718_n N_A_991_365#_c_757_n 0.0126007f $X=8.36 $Y=0.995 $X2=0 $Y2=0
cc_555 A N_A_991_365#_c_757_n 0.0320801f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_556 N_A_c_717_n N_A_991_365#_c_758_n 0.00444032f $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_557 A N_A_991_365#_c_758_n 0.0205785f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_558 N_A_c_717_n N_A_991_365#_c_759_n 6.12146e-19 $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_559 N_A_c_718_n N_A_991_365#_c_759_n 0.00283691f $X=8.36 $Y=0.995 $X2=0 $Y2=0
cc_560 A N_A_991_365#_c_759_n 0.0166196f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_561 N_A_c_717_n N_A_991_365#_c_766_n 0.00264548f $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_562 A N_A_991_365#_c_789_n 9.51454e-19 $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_563 N_A_c_717_n N_VPWR_c_907_n 0.00392692f $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_564 N_A_c_717_n N_VPWR_c_916_n 0.0030886f $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_565 N_A_c_717_n N_VPWR_c_917_n 0.0165091f $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_566 N_A_c_717_n N_A_424_49#_c_1167_n 0.00147486f $X=8.335 $Y=1.41 $X2=0 $Y2=0
cc_567 N_A_c_717_n N_A_1276_297#_c_1351_n 0.0148572f $X=8.335 $Y=1.41 $X2=0
+ $Y2=0
cc_568 N_A_c_717_n N_A_1276_297#_c_1344_n 2.98504e-19 $X=8.335 $Y=1.41 $X2=0
+ $Y2=0
cc_569 N_A_c_718_n N_VGND_c_1406_n 0.00616303f $X=8.36 $Y=0.995 $X2=0 $Y2=0
cc_570 N_A_c_718_n N_VGND_c_1411_n 0.00439206f $X=8.36 $Y=0.995 $X2=0 $Y2=0
cc_571 N_A_c_718_n N_VGND_c_1413_n 0.00704273f $X=8.36 $Y=0.995 $X2=0 $Y2=0
cc_572 N_A_991_365#_c_764_n N_VPWR_M1016_d 0.0155096f $X=8.945 $Y=1.6 $X2=0
+ $Y2=0
cc_573 N_A_991_365#_c_754_n N_VPWR_c_912_n 0.00435494f $X=9.115 $Y=1.41 $X2=0
+ $Y2=0
cc_574 N_A_991_365#_M1010_d N_VPWR_c_907_n 0.00402227f $X=7.87 $Y=1.645 $X2=0
+ $Y2=0
cc_575 N_A_991_365#_c_754_n N_VPWR_c_907_n 0.00588473f $X=9.115 $Y=1.41 $X2=0
+ $Y2=0
cc_576 N_A_991_365#_c_754_n N_VPWR_c_917_n 0.0135108f $X=9.115 $Y=1.41 $X2=0
+ $Y2=0
cc_577 N_A_991_365#_c_776_n N_A_406_325#_M1009_d 0.00419658f $X=7.945 $Y=0.51
+ $X2=0 $Y2=0
cc_578 N_A_991_365#_c_776_n N_A_406_325#_c_1005_n 0.014738f $X=7.945 $Y=0.51
+ $X2=0 $Y2=0
cc_579 N_A_991_365#_c_776_n N_A_406_325#_c_1056_n 0.00610486f $X=7.945 $Y=0.51
+ $X2=0 $Y2=0
cc_580 N_A_991_365#_c_776_n N_A_406_325#_c_1057_n 0.00980954f $X=7.945 $Y=0.51
+ $X2=0 $Y2=0
cc_581 N_A_991_365#_c_789_n N_A_406_325#_c_1057_n 0.0012274f $X=8.09 $Y=0.51
+ $X2=0 $Y2=0
cc_582 N_A_991_365#_c_790_n N_A_406_325#_c_1057_n 0.00676871f $X=8.09 $Y=0.51
+ $X2=0 $Y2=0
cc_583 N_A_991_365#_c_776_n N_A_406_325#_c_1078_n 0.0119237f $X=7.945 $Y=0.51
+ $X2=0 $Y2=0
cc_584 N_A_991_365#_M1011_s N_A_406_325#_c_1011_n 0.00764502f $X=4.955 $Y=1.825
+ $X2=0 $Y2=0
cc_585 N_A_991_365#_c_756_n N_A_406_325#_c_1011_n 0.0182772f $X=5.08 $Y=1.94
+ $X2=0 $Y2=0
cc_586 N_A_991_365#_c_776_n N_A_424_49#_M1004_d 0.00606718f $X=7.945 $Y=0.51
+ $X2=0 $Y2=0
cc_587 N_A_991_365#_c_756_n N_A_424_49#_c_1162_n 0.0138372f $X=5.08 $Y=1.94
+ $X2=0 $Y2=0
cc_588 N_A_991_365#_c_756_n N_A_424_49#_c_1163_n 0.0028603f $X=5.08 $Y=1.94
+ $X2=0 $Y2=0
cc_589 N_A_991_365#_M1011_s N_A_424_49#_c_1164_n 0.0104901f $X=4.955 $Y=1.825
+ $X2=0 $Y2=0
cc_590 N_A_991_365#_c_756_n N_A_424_49#_c_1164_n 0.0128549f $X=5.08 $Y=1.94
+ $X2=0 $Y2=0
cc_591 N_A_991_365#_c_756_n N_A_424_49#_c_1155_n 0.067594f $X=5.08 $Y=1.94 $X2=0
+ $Y2=0
cc_592 N_A_991_365#_M1010_d N_A_424_49#_c_1167_n 0.0026089f $X=7.87 $Y=1.645
+ $X2=0 $Y2=0
cc_593 N_A_991_365#_c_776_n N_A_424_49#_c_1212_n 0.0125744f $X=7.945 $Y=0.51
+ $X2=0 $Y2=0
cc_594 N_A_991_365#_c_760_n N_A_424_49#_c_1212_n 0.00143452f $X=5.275 $Y=0.51
+ $X2=0 $Y2=0
cc_595 N_A_991_365#_c_761_n N_A_424_49#_c_1212_n 0.00335094f $X=5.13 $Y=0.51
+ $X2=0 $Y2=0
cc_596 N_A_991_365#_M1004_s N_A_424_49#_c_1157_n 0.00157756f $X=5.12 $Y=0.245
+ $X2=0 $Y2=0
cc_597 N_A_991_365#_c_756_n N_A_424_49#_c_1157_n 0.0123139f $X=5.08 $Y=1.94
+ $X2=0 $Y2=0
cc_598 N_A_991_365#_c_776_n N_A_424_49#_c_1157_n 0.00370418f $X=7.945 $Y=0.51
+ $X2=0 $Y2=0
cc_599 N_A_991_365#_c_761_n N_A_424_49#_c_1157_n 0.0020377f $X=5.13 $Y=0.51
+ $X2=0 $Y2=0
cc_600 N_A_991_365#_c_776_n N_A_1276_297#_M1008_d 0.00653094f $X=7.945 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_601 N_A_991_365#_c_776_n N_A_1276_297#_c_1338_n 0.00162336f $X=7.945 $Y=0.51
+ $X2=0 $Y2=0
cc_602 N_A_991_365#_c_754_n N_A_1276_297#_c_1339_n 0.0195627f $X=9.115 $Y=1.41
+ $X2=0 $Y2=0
cc_603 N_A_991_365#_c_755_n N_A_1276_297#_c_1339_n 0.0097849f $X=9.14 $Y=0.995
+ $X2=0 $Y2=0
cc_604 N_A_991_365#_c_764_n N_A_1276_297#_c_1339_n 0.0112214f $X=8.945 $Y=1.6
+ $X2=0 $Y2=0
cc_605 N_A_991_365#_c_759_n N_A_1276_297#_c_1339_n 0.0381742f $X=9.03 $Y=1.325
+ $X2=0 $Y2=0
cc_606 N_A_991_365#_c_766_n N_A_1276_297#_c_1339_n 0.00830381f $X=9.03 $Y=1.495
+ $X2=0 $Y2=0
cc_607 N_A_991_365#_M1010_d N_A_1276_297#_c_1351_n 0.00774465f $X=7.87 $Y=1.645
+ $X2=0 $Y2=0
cc_608 N_A_991_365#_c_754_n N_A_1276_297#_c_1351_n 0.00344895f $X=9.115 $Y=1.41
+ $X2=0 $Y2=0
cc_609 N_A_991_365#_c_764_n N_A_1276_297#_c_1351_n 0.0536865f $X=8.945 $Y=1.6
+ $X2=0 $Y2=0
cc_610 N_A_991_365#_c_754_n N_A_1276_297#_c_1344_n 0.0129179f $X=9.115 $Y=1.41
+ $X2=0 $Y2=0
cc_611 N_A_991_365#_c_764_n N_A_1276_297#_c_1344_n 0.00653478f $X=8.945 $Y=1.6
+ $X2=0 $Y2=0
cc_612 N_A_991_365#_c_759_n N_A_1276_297#_c_1344_n 0.00278512f $X=9.03 $Y=1.325
+ $X2=0 $Y2=0
cc_613 N_A_991_365#_c_754_n N_A_1276_297#_c_1340_n 2.03932e-19 $X=9.115 $Y=1.41
+ $X2=0 $Y2=0
cc_614 N_A_991_365#_c_757_n N_VGND_M1000_d 0.00647663f $X=8.945 $Y=0.82 $X2=0
+ $Y2=0
cc_615 N_A_991_365#_c_759_n N_VGND_M1000_d 0.00128228f $X=9.03 $Y=1.325 $X2=0
+ $Y2=0
cc_616 N_A_991_365#_c_755_n N_VGND_c_1406_n 0.00734879f $X=9.14 $Y=0.995 $X2=0
+ $Y2=0
cc_617 N_A_991_365#_c_757_n N_VGND_c_1406_n 0.0346839f $X=8.945 $Y=0.82 $X2=0
+ $Y2=0
cc_618 N_A_991_365#_c_789_n N_VGND_c_1406_n 0.00124328f $X=8.09 $Y=0.51 $X2=0
+ $Y2=0
cc_619 N_A_991_365#_c_757_n N_VGND_c_1411_n 0.00248202f $X=8.945 $Y=0.82 $X2=0
+ $Y2=0
cc_620 N_A_991_365#_c_776_n N_VGND_c_1411_n 0.00575847f $X=7.945 $Y=0.51 $X2=0
+ $Y2=0
cc_621 N_A_991_365#_c_760_n N_VGND_c_1411_n 2.49898e-19 $X=5.275 $Y=0.51 $X2=0
+ $Y2=0
cc_622 N_A_991_365#_c_761_n N_VGND_c_1411_n 0.0254286f $X=5.13 $Y=0.51 $X2=0
+ $Y2=0
cc_623 N_A_991_365#_c_789_n N_VGND_c_1411_n 3.63685e-19 $X=8.09 $Y=0.51 $X2=0
+ $Y2=0
cc_624 N_A_991_365#_c_790_n N_VGND_c_1411_n 0.0149689f $X=8.09 $Y=0.51 $X2=0
+ $Y2=0
cc_625 N_A_991_365#_c_755_n N_VGND_c_1412_n 0.00536613f $X=9.14 $Y=0.995 $X2=0
+ $Y2=0
cc_626 N_A_991_365#_c_759_n N_VGND_c_1412_n 0.00214688f $X=9.03 $Y=1.325 $X2=0
+ $Y2=0
cc_627 N_A_991_365#_M1014_d N_VGND_c_1413_n 0.00244776f $X=7.88 $Y=0.235 $X2=0
+ $Y2=0
cc_628 N_A_991_365#_c_755_n N_VGND_c_1413_n 0.0108777f $X=9.14 $Y=0.995 $X2=0
+ $Y2=0
cc_629 N_A_991_365#_c_757_n N_VGND_c_1413_n 0.00697395f $X=8.945 $Y=0.82 $X2=0
+ $Y2=0
cc_630 N_A_991_365#_c_759_n N_VGND_c_1413_n 0.00449391f $X=9.03 $Y=1.325 $X2=0
+ $Y2=0
cc_631 N_A_991_365#_c_776_n N_VGND_c_1413_n 0.232956f $X=7.945 $Y=0.51 $X2=0
+ $Y2=0
cc_632 N_A_991_365#_c_760_n N_VGND_c_1413_n 0.0285546f $X=5.275 $Y=0.51 $X2=0
+ $Y2=0
cc_633 N_A_991_365#_c_761_n N_VGND_c_1413_n 0.00396297f $X=5.13 $Y=0.51 $X2=0
+ $Y2=0
cc_634 N_A_991_365#_c_789_n N_VGND_c_1413_n 0.0285254f $X=8.09 $Y=0.51 $X2=0
+ $Y2=0
cc_635 N_A_991_365#_c_790_n N_VGND_c_1413_n 0.0036194f $X=8.09 $Y=0.51 $X2=0
+ $Y2=0
cc_636 X N_VPWR_c_908_n 0.0164984f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_637 X N_VPWR_c_911_n 0.0350126f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_638 N_X_M1019_s N_VPWR_c_907_n 0.00233913f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_639 X N_VPWR_c_907_n 0.0199823f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_640 N_X_c_883_n N_VGND_c_1404_n 0.0112664f $X=0.425 $Y=0.56 $X2=0 $Y2=0
cc_641 N_X_c_883_n N_VGND_c_1407_n 0.0208694f $X=0.425 $Y=0.56 $X2=0 $Y2=0
cc_642 N_X_M1018_s N_VGND_c_1413_n 0.00236581f $X=0.3 $Y=0.235 $X2=0 $Y2=0
cc_643 N_X_c_883_n N_VGND_c_1413_n 0.018324f $X=0.425 $Y=0.56 $X2=0 $Y2=0
cc_644 N_VPWR_c_909_n N_A_406_325#_c_1006_n 0.00407465f $X=3.885 $Y=2.72 $X2=0
+ $Y2=0
cc_645 N_VPWR_c_907_n N_A_406_325#_c_1006_n 0.0092333f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_646 N_VPWR_M1006_s N_A_406_325#_c_1011_n 0.00109947f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_647 N_VPWR_c_907_n N_A_424_49#_M1012_d 0.00241089f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_648 N_VPWR_c_909_n N_A_424_49#_c_1159_n 0.00296166f $X=3.885 $Y=2.72 $X2=0
+ $Y2=0
cc_649 N_VPWR_c_910_n N_A_424_49#_c_1159_n 0.00147971f $X=4.05 $Y=2.32 $X2=0
+ $Y2=0
cc_650 N_VPWR_c_907_n N_A_424_49#_c_1159_n 0.00485654f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_651 N_VPWR_M1006_s N_A_424_49#_c_1154_n 0.00659923f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_652 N_VPWR_M1006_s N_A_424_49#_c_1162_n 0.00155527f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_653 N_VPWR_c_910_n N_A_424_49#_c_1162_n 0.00612755f $X=4.05 $Y=2.32 $X2=0
+ $Y2=0
cc_654 N_VPWR_c_907_n N_A_424_49#_c_1162_n 0.0119497f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_655 N_VPWR_c_916_n N_A_424_49#_c_1162_n 0.00666556f $X=8.355 $Y=2.54 $X2=0
+ $Y2=0
cc_656 N_VPWR_c_910_n N_A_424_49#_c_1163_n 0.00140976f $X=4.05 $Y=2.32 $X2=0
+ $Y2=0
cc_657 N_VPWR_c_907_n N_A_424_49#_c_1164_n 0.0189426f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_658 N_VPWR_c_916_n N_A_424_49#_c_1164_n 0.0294498f $X=8.355 $Y=2.54 $X2=0
+ $Y2=0
cc_659 N_VPWR_c_910_n N_A_424_49#_c_1165_n 0.00679194f $X=4.05 $Y=2.32 $X2=0
+ $Y2=0
cc_660 N_VPWR_c_907_n N_A_424_49#_c_1165_n 0.00644066f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_661 N_VPWR_c_916_n N_A_424_49#_c_1165_n 0.0105745f $X=8.355 $Y=2.54 $X2=0
+ $Y2=0
cc_662 N_VPWR_c_907_n N_A_424_49#_c_1167_n 0.0814431f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_916_n N_A_424_49#_c_1167_n 0.135241f $X=8.355 $Y=2.54 $X2=0
+ $Y2=0
cc_664 N_VPWR_c_917_n N_A_424_49#_c_1167_n 0.00742618f $X=9.05 $Y=2.54 $X2=0
+ $Y2=0
cc_665 N_VPWR_c_909_n N_A_424_49#_c_1168_n 0.0186431f $X=3.885 $Y=2.72 $X2=0
+ $Y2=0
cc_666 N_VPWR_c_910_n N_A_424_49#_c_1168_n 0.0142739f $X=4.05 $Y=2.32 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_907_n N_A_424_49#_c_1168_n 0.0145279f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_668 N_VPWR_M1006_s N_A_424_49#_c_1169_n 0.00243878f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_910_n N_A_424_49#_c_1169_n 0.0143988f $X=4.05 $Y=2.32 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_907_n N_A_424_49#_c_1169_n 8.22076e-19 $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_907_n N_A_424_49#_c_1170_n 0.00590105f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_672 N_VPWR_c_916_n N_A_424_49#_c_1170_n 0.010368f $X=8.355 $Y=2.54 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_907_n N_A_1276_297#_M1013_d 0.00259864f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_674 N_VPWR_c_912_n N_A_1276_297#_c_1342_n 0.0197624f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_675 N_VPWR_c_907_n N_A_1276_297#_c_1342_n 0.0111058f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_917_n N_A_1276_297#_c_1342_n 0.0126729f $X=9.05 $Y=2.54 $X2=0
+ $Y2=0
cc_677 N_VPWR_M1016_d N_A_1276_297#_c_1351_n 0.0130816f $X=8.425 $Y=1.485 $X2=0
+ $Y2=0
cc_678 N_VPWR_c_907_n N_A_1276_297#_c_1351_n 0.0163551f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_679 N_VPWR_c_916_n N_A_1276_297#_c_1351_n 0.00691204f $X=8.355 $Y=2.54 $X2=0
+ $Y2=0
cc_680 N_VPWR_c_917_n N_A_1276_297#_c_1351_n 0.0433445f $X=9.05 $Y=2.54 $X2=0
+ $Y2=0
cc_681 N_VPWR_c_912_n N_A_1276_297#_c_1344_n 0.0034505f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_682 N_VPWR_c_907_n N_A_1276_297#_c_1344_n 0.00562459f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_683 N_A_406_325#_c_1006_n N_A_424_49#_M1017_d 0.00645539f $X=3.205 $Y=1.98
+ $X2=0 $Y2=0
cc_684 N_A_406_325#_c_1026_n N_A_424_49#_M1017_d 0.00677252f $X=3.29 $Y=1.895
+ $X2=0 $Y2=0
cc_685 N_A_406_325#_c_1014_n N_A_424_49#_M1017_d 0.00697789f $X=3.535 $Y=1.535
+ $X2=0 $Y2=0
cc_686 N_A_406_325#_M1020_d N_A_424_49#_c_1151_n 0.00334341f $X=3.19 $Y=0.245
+ $X2=0 $Y2=0
cc_687 N_A_406_325#_c_1004_n N_A_424_49#_c_1151_n 0.0138308f $X=3.535 $Y=0.76
+ $X2=0 $Y2=0
cc_688 N_A_406_325#_M1020_d N_A_424_49#_c_1175_n 0.00348437f $X=3.19 $Y=0.245
+ $X2=0 $Y2=0
cc_689 N_A_406_325#_c_1004_n N_A_424_49#_c_1175_n 0.00440606f $X=3.535 $Y=0.76
+ $X2=0 $Y2=0
cc_690 N_A_406_325#_M1020_d N_A_424_49#_c_1152_n 0.0175141f $X=3.19 $Y=0.245
+ $X2=0 $Y2=0
cc_691 N_A_406_325#_c_1004_n N_A_424_49#_c_1152_n 0.0128008f $X=3.535 $Y=0.76
+ $X2=0 $Y2=0
cc_692 N_A_406_325#_M1020_d N_A_424_49#_c_1176_n 3.2099e-19 $X=3.19 $Y=0.245
+ $X2=0 $Y2=0
cc_693 N_A_406_325#_c_1011_n N_A_424_49#_c_1159_n 0.00437461f $X=5.955 $Y=1.53
+ $X2=0 $Y2=0
cc_694 N_A_406_325#_c_1012_n N_A_424_49#_c_1159_n 0.00277011f $X=3.795 $Y=1.53
+ $X2=0 $Y2=0
cc_695 N_A_406_325#_c_1014_n N_A_424_49#_c_1159_n 0.00125154f $X=3.535 $Y=1.535
+ $X2=0 $Y2=0
cc_696 N_A_406_325#_c_1006_n N_A_424_49#_c_1160_n 0.0153275f $X=3.205 $Y=1.98
+ $X2=0 $Y2=0
cc_697 N_A_406_325#_c_1012_n N_A_424_49#_c_1160_n 0.00119193f $X=3.795 $Y=1.53
+ $X2=0 $Y2=0
cc_698 N_A_406_325#_c_1014_n N_A_424_49#_c_1160_n 0.0114314f $X=3.535 $Y=1.535
+ $X2=0 $Y2=0
cc_699 N_A_406_325#_c_1004_n N_A_424_49#_c_1153_n 0.0327455f $X=3.535 $Y=0.76
+ $X2=0 $Y2=0
cc_700 N_A_406_325#_c_1026_n N_A_424_49#_c_1154_n 0.00649967f $X=3.29 $Y=1.895
+ $X2=0 $Y2=0
cc_701 N_A_406_325#_c_1004_n N_A_424_49#_c_1154_n 0.00891656f $X=3.535 $Y=0.76
+ $X2=0 $Y2=0
cc_702 N_A_406_325#_c_1011_n N_A_424_49#_c_1154_n 0.0161183f $X=5.955 $Y=1.53
+ $X2=0 $Y2=0
cc_703 N_A_406_325#_c_1012_n N_A_424_49#_c_1154_n 0.00275249f $X=3.795 $Y=1.53
+ $X2=0 $Y2=0
cc_704 N_A_406_325#_c_1014_n N_A_424_49#_c_1154_n 0.0233325f $X=3.535 $Y=1.535
+ $X2=0 $Y2=0
cc_705 N_A_406_325#_c_1011_n N_A_424_49#_c_1162_n 0.011487f $X=5.955 $Y=1.53
+ $X2=0 $Y2=0
cc_706 N_A_406_325#_c_1008_n N_A_424_49#_c_1155_n 0.00833378f $X=5.952 $Y=1.615
+ $X2=0 $Y2=0
cc_707 N_A_406_325#_c_1043_n N_A_424_49#_c_1155_n 0.0247324f $X=5.92 $Y=1.62
+ $X2=0 $Y2=0
cc_708 N_A_406_325#_c_1011_n N_A_424_49#_c_1155_n 0.0194987f $X=5.955 $Y=1.53
+ $X2=0 $Y2=0
cc_709 N_A_406_325#_c_1013_n N_A_424_49#_c_1155_n 0.00126802f $X=6.1 $Y=1.53
+ $X2=0 $Y2=0
cc_710 N_A_406_325#_M1011_d N_A_424_49#_c_1167_n 0.0094538f $X=5.57 $Y=1.485
+ $X2=0 $Y2=0
cc_711 N_A_406_325#_c_1043_n N_A_424_49#_c_1167_n 0.0238103f $X=5.92 $Y=1.62
+ $X2=0 $Y2=0
cc_712 N_A_406_325#_c_1009_n N_A_424_49#_c_1167_n 0.0100462f $X=6.405 $Y=1.53
+ $X2=0 $Y2=0
cc_713 N_A_406_325#_c_1005_n N_A_424_49#_c_1212_n 0.00250545f $X=6.49 $Y=1.445
+ $X2=0 $Y2=0
cc_714 N_A_406_325#_c_1006_n N_A_424_49#_c_1168_n 0.0049241f $X=3.205 $Y=1.98
+ $X2=0 $Y2=0
cc_715 N_A_406_325#_c_1012_n N_A_424_49#_c_1168_n 2.48159e-19 $X=3.795 $Y=1.53
+ $X2=0 $Y2=0
cc_716 N_A_406_325#_c_1014_n N_A_424_49#_c_1168_n 0.00535873f $X=3.535 $Y=1.535
+ $X2=0 $Y2=0
cc_717 N_A_406_325#_c_1004_n N_A_424_49#_c_1156_n 0.0132287f $X=3.535 $Y=0.76
+ $X2=0 $Y2=0
cc_718 N_A_406_325#_c_1011_n N_A_424_49#_c_1156_n 0.0052436f $X=5.955 $Y=1.53
+ $X2=0 $Y2=0
cc_719 N_A_406_325#_c_1012_n N_A_424_49#_c_1156_n 2.29009e-19 $X=3.795 $Y=1.53
+ $X2=0 $Y2=0
cc_720 N_A_406_325#_c_1008_n N_A_424_49#_c_1157_n 2.53366e-19 $X=5.952 $Y=1.615
+ $X2=0 $Y2=0
cc_721 N_A_406_325#_c_1011_n N_A_424_49#_c_1157_n 9.70582e-19 $X=5.955 $Y=1.53
+ $X2=0 $Y2=0
cc_722 N_A_406_325#_c_1005_n N_A_1276_297#_M1008_d 0.00729398f $X=6.49 $Y=1.445
+ $X2=-0.19 $Y2=-0.24
cc_723 N_A_406_325#_c_1137_p N_A_1276_297#_M1008_d 0.0024562f $X=6.575 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_724 N_A_406_325#_c_1078_n N_A_1276_297#_M1008_d 0.0107136f $X=7.085 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_725 N_A_406_325#_c_1009_n N_A_1276_297#_M1015_d 0.00444096f $X=6.405 $Y=1.53
+ $X2=0 $Y2=0
cc_726 N_A_406_325#_c_1043_n N_A_1276_297#_c_1338_n 0.00453141f $X=5.92 $Y=1.62
+ $X2=0 $Y2=0
cc_727 N_A_406_325#_c_1009_n N_A_1276_297#_c_1338_n 0.013519f $X=6.405 $Y=1.53
+ $X2=0 $Y2=0
cc_728 N_A_406_325#_c_1005_n N_A_1276_297#_c_1338_n 0.062318f $X=6.49 $Y=1.445
+ $X2=0 $Y2=0
cc_729 N_A_406_325#_c_1078_n N_A_1276_297#_c_1338_n 0.0106102f $X=7.085 $Y=0.36
+ $X2=0 $Y2=0
cc_730 N_A_406_325#_c_1013_n N_A_1276_297#_c_1338_n 0.00130235f $X=6.1 $Y=1.53
+ $X2=0 $Y2=0
cc_731 N_A_406_325#_c_1011_n N_VGND_c_1405_n 0.00558664f $X=5.955 $Y=1.53 $X2=0
+ $Y2=0
cc_732 N_A_406_325#_c_1137_p N_VGND_c_1411_n 0.0104913f $X=6.575 $Y=0.34 $X2=0
+ $Y2=0
cc_733 N_A_406_325#_c_1078_n N_VGND_c_1411_n 0.0617902f $X=7.085 $Y=0.36 $X2=0
+ $Y2=0
cc_734 N_A_406_325#_M1009_d N_VGND_c_1413_n 0.00226821f $X=7.185 $Y=0.245 $X2=0
+ $Y2=0
cc_735 N_A_406_325#_c_1137_p N_VGND_c_1413_n 0.00184693f $X=6.575 $Y=0.34 $X2=0
+ $Y2=0
cc_736 N_A_406_325#_c_1078_n N_VGND_c_1413_n 0.00974346f $X=7.085 $Y=0.36 $X2=0
+ $Y2=0
cc_737 N_A_424_49#_c_1167_n N_A_1276_297#_M1015_d 0.00563686f $X=7.535 $Y=2.36
+ $X2=0 $Y2=0
cc_738 N_A_424_49#_c_1167_n N_A_1276_297#_c_1350_n 0.0129278f $X=7.535 $Y=2.36
+ $X2=0 $Y2=0
cc_739 N_A_424_49#_M1012_d N_A_1276_297#_c_1351_n 0.00610222f $X=7.305 $Y=1.645
+ $X2=0 $Y2=0
cc_740 N_A_424_49#_c_1167_n N_A_1276_297#_c_1351_n 0.0533312f $X=7.535 $Y=2.36
+ $X2=0 $Y2=0
cc_741 N_A_424_49#_c_1152_n N_VGND_c_1405_n 0.0141318f $X=3.79 $Y=0.34 $X2=0
+ $Y2=0
cc_742 N_A_424_49#_c_1153_n N_VGND_c_1405_n 0.0321795f $X=3.875 $Y=1.035 $X2=0
+ $Y2=0
cc_743 N_A_424_49#_c_1151_n N_VGND_c_1409_n 0.00239374f $X=3.06 $Y=0.74 $X2=0
+ $Y2=0
cc_744 N_A_424_49#_c_1152_n N_VGND_c_1409_n 0.0445697f $X=3.79 $Y=0.34 $X2=0
+ $Y2=0
cc_745 N_A_424_49#_c_1176_n N_VGND_c_1409_n 0.0130641f $X=3.28 $Y=0.34 $X2=0
+ $Y2=0
cc_746 N_A_424_49#_c_1212_n N_VGND_c_1411_n 0.00800682f $X=5.715 $Y=0.545 $X2=0
+ $Y2=0
cc_747 N_A_424_49#_c_1157_n N_VGND_c_1411_n 0.0028353f $X=5.42 $Y=0.772 $X2=0
+ $Y2=0
cc_748 N_A_424_49#_c_1151_n N_VGND_c_1413_n 0.00649067f $X=3.06 $Y=0.74 $X2=0
+ $Y2=0
cc_749 N_A_424_49#_c_1152_n N_VGND_c_1413_n 0.0255342f $X=3.79 $Y=0.34 $X2=0
+ $Y2=0
cc_750 N_A_424_49#_c_1176_n N_VGND_c_1413_n 0.00783952f $X=3.28 $Y=0.34 $X2=0
+ $Y2=0
cc_751 N_A_424_49#_c_1212_n N_VGND_c_1413_n 0.0018012f $X=5.715 $Y=0.545 $X2=0
+ $Y2=0
cc_752 N_A_1276_297#_c_1340_n N_VGND_c_1412_n 0.0197576f $X=9.48 $Y=0.42 $X2=0
+ $Y2=0
cc_753 N_A_1276_297#_M1021_d N_VGND_c_1413_n 0.00399944f $X=9.215 $Y=0.235 $X2=0
+ $Y2=0
cc_754 N_A_1276_297#_c_1340_n N_VGND_c_1413_n 0.0113402f $X=9.48 $Y=0.42 $X2=0
+ $Y2=0
