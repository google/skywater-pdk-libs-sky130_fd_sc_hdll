* File: sky130_fd_sc_hdll__or2_2.pex.spice
* Created: Thu Aug 27 19:23:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR2_2%B 3 5 7 8 9 15
r27 15 16 4.66022 $w=3.62e-07 $l=3.5e-08 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.555 $Y2=1.202
r28 13 15 34.6188 $w=3.62e-07 $l=2.6e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.52 $Y2=1.202
r29 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r30 8 9 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=0.235 $Y=0.85 $X2=0.235
+ $Y2=1.16
r31 5 16 19.0988 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.555 $Y=1.41
+ $X2=0.555 $Y2=1.202
r32 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.555 $Y=1.41
+ $X2=0.555 $Y2=1.695
r33 1 15 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_2%A 3 5 7 8 9
r33 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r34 9 14 0.780051 $w=4.58e-07 $l=3e-08 $layer=LI1_cond $X=1.145 $Y=1.19
+ $X2=1.145 $Y2=1.16
r35 8 14 8.06053 $w=4.58e-07 $l=3.1e-07 $layer=LI1_cond $X=1.145 $Y=0.85
+ $X2=1.145 $Y2=1.16
r36 5 13 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=1.025 $Y2=1.16
r37 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.695
r38 1 13 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=1.025 $Y2=1.16
r39 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_2%A_39_297# 1 2 7 9 10 12 13 15 16 18 20 21 22
+ 25 32 38
c71 25 0 7.50958e-20 $X=1.63 $Y=1.16
c72 20 0 1.05688e-19 $X=0.63 $Y=1.495
r73 38 39 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.99 $Y=1.202
+ $X2=2.015 $Y2=1.202
r74 35 36 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.495 $Y=1.202
+ $X2=1.52 $Y2=1.202
r75 32 34 6.80499 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.685 $Y=0.43
+ $X2=0.685 $Y2=0.595
r76 26 38 45.6632 $w=3.8e-07 $l=3.6e-07 $layer=POLY_cond $X=1.63 $Y=1.202
+ $X2=1.99 $Y2=1.202
r77 26 36 13.9526 $w=3.8e-07 $l=1.1e-07 $layer=POLY_cond $X=1.63 $Y=1.202
+ $X2=1.52 $Y2=1.202
r78 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.16 $X2=1.63 $Y2=1.16
r79 23 25 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=1.655 $Y=1.495
+ $X2=1.655 $Y2=1.16
r80 21 23 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.545 $Y=1.58
+ $X2=1.655 $Y2=1.495
r81 21 22 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.545 $Y=1.58
+ $X2=0.745 $Y2=1.58
r82 20 22 6.87116 $w=2.76e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.63 $Y=1.495
+ $X2=0.745 $Y2=1.58
r83 20 29 13.7029 $w=2.76e-07 $l=3.86549e-07 $layer=LI1_cond $X=0.63 $Y=1.495
+ $X2=0.32 $Y2=1.667
r84 20 34 45.0956 $w=2.28e-07 $l=9e-07 $layer=LI1_cond $X=0.63 $Y=1.495 $X2=0.63
+ $Y2=0.595
r85 16 39 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=1.202
r86 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=0.56
r87 13 38 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.202
r88 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.985
r89 10 36 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.52 $Y=1.41
+ $X2=1.52 $Y2=1.202
r90 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.52 $Y=1.41
+ $X2=1.52 $Y2=1.985
r91 7 35 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=1.202
r92 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=0.56
r93 2 29 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.485 $X2=0.32 $Y2=1.66
r94 1 32 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_2%VPWR 1 2 9 13 16 17 19 20 21 34 35
r34 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r35 32 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r38 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r39 24 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r40 21 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r41 21 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r42 19 31 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.14 $Y=2.72 $X2=2.07
+ $Y2=2.72
r43 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.72
+ $X2=2.225 $Y2=2.72
r44 18 34 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.225 $Y2=2.72
r46 16 28 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=2.72 $X2=1.15
+ $Y2=2.72
r47 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.72 $X2=1.285
+ $Y2=2.72
r48 15 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.37 $Y=2.72 $X2=2.07
+ $Y2=2.72
r49 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.72
+ $X2=1.285 $Y2=2.72
r50 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.72
r51 11 13 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.34
r52 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=2.72
r53 7 9 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=2.01
r54 2 13 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.485 $X2=2.225 $Y2=2.34
r55 1 9 300 $w=1.7e-07 $l=6.29583e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.285 $Y2=2.01
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_2%X 1 2 7 10 13 16
c43 2 0 7.50958e-20 $X=1.61 $Y=1.485
r44 13 16 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=1.92
+ $X2=2.175 $Y2=1.92
r45 13 16 0.622958 $w=4.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.175 $Y=1.81
+ $X2=2.175 $Y2=1.835
r46 12 13 24.5445 $w=4.78e-07 $l=9.85e-07 $layer=LI1_cond $X=2.175 $Y=0.825
+ $X2=2.175 $Y2=1.81
r47 10 12 22.1818 $w=2.31e-07 $l=4.2e-07 $layer=LI1_cond $X=1.755 $Y=0.655
+ $X2=2.175 $Y2=0.655
r48 7 13 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.73 $Y=1.92 $X2=2.07
+ $Y2=1.92
r49 2 7 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.61
+ $Y=1.485 $X2=1.755 $Y2=2
r50 1 10 182 $w=1.7e-07 $l=4.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.235 $X2=1.755 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_2%VGND 1 2 3 10 12 14 18 20 24 26 30 31 37 40
r43 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r44 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r45 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r46 31 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r47 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r48 28 40 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.2
+ $Y2=0
r49 28 30 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.53
+ $Y2=0
r50 26 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r51 26 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r52 22 40 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0.085 $X2=2.2
+ $Y2=0
r53 22 24 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=2.2 $Y=0.085
+ $X2=2.2 $Y2=0.39
r54 21 37 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.292
+ $Y2=0
r55 20 40 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.2
+ $Y2=0
r56 20 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.45
+ $Y2=0
r57 16 37 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.292 $Y=0.085
+ $X2=1.292 $Y2=0
r58 16 18 12.622 $w=3.13e-07 $l=3.45e-07 $layer=LI1_cond $X=1.292 $Y=0.085
+ $X2=1.292 $Y2=0.43
r59 15 34 3.93736 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r60 14 37 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.292
+ $Y2=0
r61 14 15 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.345
+ $Y2=0
r62 10 34 3.14078 $w=2.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.172 $Y2=0
r63 10 12 16.5664 $w=2.38e-07 $l=3.45e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.43
r64 3 24 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.235 $X2=2.225 $Y2=0.39
r65 2 18 182 $w=1.7e-07 $l=3.49142e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.28 $Y2=0.43
r66 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

