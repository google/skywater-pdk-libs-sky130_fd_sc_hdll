* File: sky130_fd_sc_hdll__a22oi_1.pex.spice
* Created: Thu Aug 27 18:54:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A22OI_1%B2 1 3 4 6 7 8
c28 1 0 7.47939e-20 $X=0.495 $Y=1.41
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r30 8 13 0.717647 $w=4.98e-07 $l=3e-08 $layer=LI1_cond $X=0.375 $Y=1.19
+ $X2=0.375 $Y2=1.16
r31 7 13 7.41569 $w=4.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.375 $Y=0.85
+ $X2=0.375 $Y2=1.16
r32 4 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.435 $Y2=1.16
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r34 1 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.435 $Y2=1.16
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_1%B1 1 3 4 6 7 8 22
c35 7 0 2.28009e-19 $X=1.13 $Y=0.85
c36 4 0 1.67017e-19 $X=0.965 $Y=1.41
r37 14 22 1.94091 $w=1.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.19 $Y=1.175
+ $X2=1.155 $Y2=1.175
r38 13 22 8.59545 $w=1.98e-07 $l=1.55e-07 $layer=LI1_cond $X=1 $Y=1.175
+ $X2=1.155 $Y2=1.175
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r40 8 14 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=1.23 $Y=1.175 $X2=1.19
+ $Y2=1.175
r41 7 14 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=1.19 $Y=0.85 $X2=1.19
+ $Y2=1.075
r42 4 12 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=1 $Y2=1.16
r43 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r44 1 12 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=1 $Y2=1.16
r45 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_1%A1 1 3 4 6 7 8 14 15
c32 7 0 1.67017e-19 $X=1.635 $Y=0.85
c33 1 0 1.93103e-19 $X=1.955 $Y=1.41
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.16 $X2=1.92 $Y2=1.16
r35 8 15 3.48996 $w=2.1e-07 $l=1.1e-07 $layer=LI1_cond $X=1.63 $Y=1.165 $X2=1.63
+ $Y2=1.055
r36 8 14 7.63857 $w=3.88e-07 $l=1.85e-07 $layer=LI1_cond $X=1.735 $Y=1.165
+ $X2=1.92 $Y2=1.165
r37 7 15 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=1.63 $Y=0.85
+ $X2=1.63 $Y2=1.055
r38 4 13 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.92 $Y2=1.16
r39 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.98 $Y=0.995 $X2=1.98
+ $Y2=0.56
r40 1 13 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.92 $Y2=1.16
r41 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_1%A2 1 3 4 6 7
r27 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r28 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.46 $Y2=1.16
r29 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
r30 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.46 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995 $X2=2.4
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_1%Y 1 2 3 4 15 23 24 26 27 31 32 34 35 36 42
+ 47
r78 40 42 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=0.425 $Y=1.53
+ $X2=1.615 $Y2=1.53
r79 36 42 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.715 $Y=1.53
+ $X2=1.615 $Y2=1.53
r80 35 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=1.53
+ $X2=0.425 $Y2=1.53
r81 35 47 2.46016 $w=4.98e-07 $l=4.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.66
r82 34 36 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=2.795 $Y=1.53
+ $X2=1.715 $Y2=1.53
r83 31 32 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=2.33
+ $X2=1.035 $Y2=2.33
r84 27 47 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=1.66
r85 27 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.295 $X2=0.26
+ $Y2=2.38
r86 26 34 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.965 $Y=1.445
+ $X2=2.795 $Y2=1.53
r87 25 26 21.0151 $w=3.38e-07 $l=6.2e-07 $layer=LI1_cond $X=2.965 $Y=0.825
+ $X2=2.965 $Y2=1.445
r88 23 25 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.795 $Y=0.74
+ $X2=2.965 $Y2=0.825
r89 23 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.795 $Y=0.74
+ $X2=2.275 $Y2=0.74
r90 22 24 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.185 $Y=0.655
+ $X2=2.275 $Y2=0.74
r91 21 22 9.24242 $w=1.78e-07 $l=1.5e-07 $layer=LI1_cond $X=2.185 $Y=0.505
+ $X2=2.185 $Y2=0.655
r92 17 20 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=1.16 $Y=0.38
+ $X2=1.72 $Y2=0.38
r93 15 21 7.0541 $w=2.5e-07 $l=1.63936e-07 $layer=LI1_cond $X=2.095 $Y=0.38
+ $X2=2.185 $Y2=0.505
r94 15 20 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=2.095 $Y=0.38
+ $X2=1.72 $Y2=0.38
r95 14 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.26 $Y2=2.38
r96 14 32 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=1.035 $Y2=2.38
r97 4 31 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r98 3 47 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r99 3 29 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r100 2 20 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.42
r101 1 17 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.16 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_1%A_117_297# 1 2 7 8
c21 7 0 3.98882e-20 $X=2.105 $Y=1.882
r22 7 16 7.6984 $w=1.68e-07 $l=1.18e-07 $layer=LI1_cond $X=2.19 $Y=1.882
+ $X2=2.19 $Y2=2
r23 7 8 73.3706 $w=1.93e-07 $l=1.29e-06 $layer=LI1_cond $X=2.105 $Y=1.882
+ $X2=0.815 $Y2=1.882
r24 2 16 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2
r25 1 8 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_1%VPWR 1 2 9 13 16 17 18 20 30 31 34
r38 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r39 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r40 28 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r41 28 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r42 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 25 34 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.91 $Y=2.72
+ $X2=1.732 $Y2=2.72
r44 25 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.91 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 20 34 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=1.732 $Y2=2.72
r46 20 22 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=0.23 $Y2=2.72
r47 18 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 18 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r49 16 27 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.56 $Y=2.72 $X2=2.53
+ $Y2=2.72
r50 16 17 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.56 $Y=2.72
+ $X2=2.692 $Y2=2.72
r51 15 30 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 15 17 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=2.692 $Y2=2.72
r53 11 17 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.692 $Y=2.635
+ $X2=2.692 $Y2=2.72
r54 11 13 26.7454 $w=2.63e-07 $l=6.15e-07 $layer=LI1_cond $X=2.692 $Y=2.635
+ $X2=2.692 $Y2=2.02
r55 7 34 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.732 $Y=2.635
+ $X2=1.732 $Y2=2.72
r56 7 9 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.732 $Y=2.635
+ $X2=1.732 $Y2=2.34
r57 2 13 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=2.02
r58 1 9 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.485 $X2=1.72 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22OI_1%VGND 1 2 7 9 13 15 17 24 25 31
r34 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r35 25 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r36 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r37 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=0 $X2=2.67
+ $Y2=0
r38 22 24 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.835 $Y=0 $X2=2.99
+ $Y2=0
r39 21 32 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r40 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r41 18 28 6.38223 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.297
+ $Y2=0
r42 18 20 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.69
+ $Y2=0
r43 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=0 $X2=2.67
+ $Y2=0
r44 17 20 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=2.505 $Y=0
+ $X2=0.69 $Y2=0
r45 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r46 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r47 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=0.085
+ $X2=2.67 $Y2=0
r48 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.67 $Y=0.085
+ $X2=2.67 $Y2=0.4
r49 7 28 2.84844 $w=5e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.297 $Y2=0
r50 7 9 10.1667 $w=4.98e-07 $l=4.25e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0.51
r51 2 13 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.67 $Y2=0.4
r52 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

