* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A3 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_493_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_485_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_1194_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_695_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_493_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND B2 a_1194_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_485_47# A2 a_695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VGND A3 a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_79_21# A1 a_695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_1194_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_79_21# B1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_79_21# B1 a_1194_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_493_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_493_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_79_21# B2 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_695_47# A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_493_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 VPWR A2 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
