* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xnor3_4 A B C VGND VNB VPB VPWR X
X0 a_1207_297# B a_657_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_101_21# a_532_93# a_681_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X2 a_657_325# C a_101_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X3 a_1490_297# B a_657_325# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X4 X a_101_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_1207_297# a_1490_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_1207_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 a_101_21# a_532_93# a_657_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 VGND B a_1089_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR C a_532_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X10 VPWR a_101_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_657_325# a_1089_297# a_1490_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 X a_101_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_1207_297# B a_681_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X14 VGND a_101_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_101_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_1207_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_681_49# C a_101_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_657_325# a_1089_297# a_1207_297# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X19 X a_101_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 X a_101_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND C a_532_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR a_101_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_681_49# a_1089_297# a_1207_297# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X24 a_1490_297# B a_681_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_681_49# a_1089_297# a_1490_297# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X26 VGND a_1207_297# a_1490_297# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 VPWR B a_1089_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
