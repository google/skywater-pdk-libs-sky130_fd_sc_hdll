* File: sky130_fd_sc_hdll__or4bb_1.spice
* Created: Wed Sep  2 08:49:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or4bb_1.pex.spice"
.subckt sky130_fd_sc_hdll__or4bb_1  VNB VPB C_N D_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_C_N_M1006_g N_A_27_410#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.1302 PD=0.72 PS=1.46 NRD=5.712 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_216_93#_M1003_d N_D_N_M1003_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1281 AS=0.063 PD=1.45 PS=0.72 NRD=11.424 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_331_413#_M1010_d N_A_216_93#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.42 AD=0.07035 AS=0.1302 PD=0.755 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_27_410#_M1007_g N_A_331_413#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.06405 AS=0.07035 PD=0.725 PS=0.755 NRD=0 NRS=17.136 M=1 R=2.8
+ SA=75000.7 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_331_413#_M1004_d N_B_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.06405 PD=0.755 PS=0.725 NRD=2.856 NRS=8.568 M=1 R=2.8
+ SA=75001.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_331_413#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0927336 AS=0.07035 PD=0.816449 PS=0.755 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75001.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_331_413#_M1009_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.143516 PD=1.85 PS=1.26355 NRD=0 NRS=11.988 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_C_N_M1011_g N_A_27_410#_M1011_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.126812 AS=0.1134 PD=1.34 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1012 N_A_216_93#_M1012_d N_D_N_M1012_g N_VPWR_M1011_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1218 AS=0.126812 PD=1.42 PS=1.34 NRD=2.3443 NRS=115.816 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1002 A_421_413# N_A_216_93#_M1002_g N_A_331_413#_M1002_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1257 AS=0.1134 PD=1.35 PS=1.38 NRD=114.575 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1013 A_527_297# N_A_27_410#_M1013_g A_421_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0483 AS=0.1257 PD=0.65 PS=1.35 NRD=28.1316 NRS=114.575 M=1 R=2.33333
+ SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1001 A_609_297# N_B_M1001_g A_527_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.06405
+ AS=0.0483 PD=0.725 PS=0.65 NRD=45.7237 NRS=28.1316 M=1 R=2.33333 SA=90000.6
+ SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g A_609_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0918972 AS=0.06405 PD=0.804507 PS=0.725 NRD=76.83 NRS=45.7237 M=1
+ R=2.33333 SA=90001.1 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1000 N_X_M1000_d N_A_331_413#_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.285 AS=0.218803 PD=2.57 PS=1.91549 NRD=0.9653 NRS=1.9503 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX15_noxref noxref_16 D_N D_N PROBETYPE=1
pX16_noxref noxref_17 A A PROBETYPE=1
pX17_noxref noxref_18 B B PROBETYPE=1
c_92 VPB 0 2.01548e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__or4bb_1.pxi.spice"
*
.ends
*
*
