* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xnor3_1 A B C VGND VNB VPB VPWR X
M1000 VPWR a_83_21# X VPB phighvt w=1e+06u l=180000u
+  ad=1.22595e+12p pd=8.52e+06u as=2.9e+11p ps=2.58e+06u
M1001 a_901_297# a_783_297# a_375_49# VNB nshort w=600000u l=150000u
+  ad=4.4975e+11p pd=3.99e+06u as=5.4545e+11p ps=4.31e+06u
M1002 a_83_21# C a_375_49# VNB nshort w=640000u l=150000u
+  ad=2.176e+11p pd=1.96e+06u as=0p ps=0u
M1003 a_1184_297# a_901_297# VGND VNB nshort w=640000u l=150000u
+  ad=5.677e+11p pd=4.42e+06u as=9.124e+11p ps=6.76e+06u
M1004 a_783_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
M1005 a_901_297# a_783_297# a_351_325# VPB phighvt w=840000u l=180000u
+  ad=7.226e+11p pd=5.29e+06u as=5.878e+11p ps=4.8e+06u
M1006 a_351_325# B a_901_297# VNB nshort w=640000u l=150000u
+  ad=6.091e+11p pd=4.57e+06u as=0p ps=0u
M1007 a_1184_297# a_901_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.998e+11p pd=5.68e+06u as=0p ps=0u
M1008 a_783_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.6515e+11p pd=1.82e+06u as=0p ps=0u
M1009 VGND A a_901_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_375_49# B a_901_297# VPB phighvt w=840000u l=180000u
+  ad=8.3175e+11p pd=5.4e+06u as=0p ps=0u
M1011 a_351_325# B a_1184_297# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_83_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.82e+11p ps=1.86e+06u
M1013 a_351_325# a_226_93# a_83_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A a_901_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_83_21# C a_351_325# VPB phighvt w=840000u l=180000u
+  ad=3.227e+11p pd=2.67e+06u as=0p ps=0u
M1016 a_1184_297# a_783_297# a_351_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_226_93# C VPWR VPB phighvt w=640000u l=180000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1018 a_1184_297# a_783_297# a_375_49# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_375_49# B a_1184_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_226_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=0p ps=0u
M1021 a_375_49# a_226_93# a_83_21# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
