* NGSPICE file created from sky130_fd_sc_hdll__dfrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 a_436_413# D VPWR VPB phighvt w=420000u l=180000u
+  ad=1.428e+11p pd=1.52e+06u as=1.3145e+12p ps=1.289e+07u
M1001 VPWR a_1323_21# a_1330_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1002 a_211_363# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.1789e+12p ps=1.006e+07u
M1003 Q a_1323_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1004 a_649_413# a_27_47# a_534_47# VPB phighvt w=420000u l=180000u
+  ad=3.318e+11p pd=3.26e+06u as=1.533e+11p ps=1.57e+06u
M1005 a_805_47# a_751_289# a_642_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.748e+11p ps=2.17e+06u
M1006 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1007 VGND RESET_B a_805_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_436_413# D VGND VNB nshort w=420000u l=150000u
+  ad=1.338e+11p pd=1.5e+06u as=0p ps=0u
M1009 VGND a_1323_21# a_1237_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.698e+11p ps=1.7e+06u
M1010 VPWR a_751_289# a_649_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_751_289# a_534_47# VGND VNB nshort w=640000u l=150000u
+  ad=1.998e+11p pd=1.97e+06u as=0p ps=0u
M1012 Q a_1323_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1013 VPWR a_1128_47# a_1323_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1014 a_1128_47# a_211_363# a_751_289# VNB nshort w=360000u l=150000u
+  ad=1.422e+11p pd=1.51e+06u as=0p ps=0u
M1015 a_534_47# a_27_47# a_436_413# VNB nshort w=360000u l=150000u
+  ad=1.404e+11p pd=1.5e+06u as=0p ps=0u
M1016 a_751_289# a_534_47# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.709e+11p pd=2.41e+06u as=0p ps=0u
M1017 a_1128_47# a_27_47# a_751_289# VPB phighvt w=420000u l=180000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1018 a_642_47# a_211_363# a_534_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1237_47# a_27_47# a_1128_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1542_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1021 a_1323_21# a_1128_47# a_1542_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1022 a_649_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1024 a_1323_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_211_363# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1026 a_534_47# a_211_363# a_436_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1330_413# a_211_363# a_1128_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

