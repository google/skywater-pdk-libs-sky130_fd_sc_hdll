* File: sky130_fd_sc_hdll__nand2_6.pex.spice
* Created: Thu Aug 27 19:13:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2_6%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 54 55
r126 55 56 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=2.87 $Y2=1.202
r127 53 55 31.9162 $w=3.7e-07 $l=2.45e-07 $layer=POLY_cond $X=2.6 $Y=1.202
+ $X2=2.845 $Y2=1.202
r128 53 54 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=2.6
+ $Y=1.16 $X2=2.6 $Y2=1.16
r129 51 53 29.3108 $w=3.7e-07 $l=2.25e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.6 $Y2=1.202
r130 50 51 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r131 49 50 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.93 $Y=1.202
+ $X2=2.35 $Y2=1.202
r132 48 49 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r133 47 48 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.905 $Y2=1.202
r134 46 47 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r135 45 46 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.41 $Y2=1.202
r136 44 45 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r137 42 44 52.7595 $w=3.7e-07 $l=4.05e-07 $layer=POLY_cond $X=0.56 $Y=1.202
+ $X2=0.965 $Y2=1.202
r138 42 43 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=0.56
+ $Y=1.16 $X2=0.56 $Y2=1.16
r139 40 42 8.46757 $w=3.7e-07 $l=6.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.56 $Y2=1.202
r140 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r141 37 54 42.2562 $w=2.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.61 $Y=1.19
+ $X2=2.6 $Y2=1.19
r142 37 43 44.8172 $w=2.68e-07 $l=1.05e-06 $layer=LI1_cond $X=1.61 $Y=1.19
+ $X2=0.56 $Y2=1.19
r143 34 56 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=1.202
r144 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=0.56
r145 31 55 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r146 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r147 28 51 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r148 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r149 25 50 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r150 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
r151 22 49 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r152 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r153 19 48 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r154 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r155 16 47 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r156 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r157 13 46 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r158 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r159 10 45 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r160 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r161 7 44 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r162 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r163 4 40 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r164 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r165 1 39 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r166 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_6%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 52 55
r105 55 56 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.665 $Y=1.202
+ $X2=5.69 $Y2=1.202
r106 54 55 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=5.195 $Y=1.202
+ $X2=5.665 $Y2=1.202
r107 53 54 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.202
+ $X2=5.195 $Y2=1.202
r108 51 53 23.4486 $w=3.7e-07 $l=1.8e-07 $layer=POLY_cond $X=4.99 $Y=1.202
+ $X2=5.17 $Y2=1.202
r109 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.99
+ $Y=1.16 $X2=4.99 $Y2=1.16
r110 49 51 31.2649 $w=3.7e-07 $l=2.4e-07 $layer=POLY_cond $X=4.75 $Y=1.202
+ $X2=4.99 $Y2=1.202
r111 48 49 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.725 $Y=1.202
+ $X2=4.75 $Y2=1.202
r112 47 48 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=4.255 $Y=1.202
+ $X2=4.725 $Y2=1.202
r113 46 47 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.202
+ $X2=4.255 $Y2=1.202
r114 44 46 33.8703 $w=3.7e-07 $l=2.6e-07 $layer=POLY_cond $X=3.97 $Y=1.202
+ $X2=4.23 $Y2=1.202
r115 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.97
+ $Y=1.16 $X2=3.97 $Y2=1.16
r116 42 44 24.1 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.97 $Y2=1.202
r117 41 42 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.202
+ $X2=3.785 $Y2=1.202
r118 40 41 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.76 $Y2=1.202
r119 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r120 37 52 26.4635 $w=2.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.37 $Y=1.19
+ $X2=4.99 $Y2=1.19
r121 37 45 17.0732 $w=2.68e-07 $l=4e-07 $layer=LI1_cond $X=4.37 $Y=1.19 $X2=3.97
+ $Y2=1.19
r122 34 56 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r123 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.56
r124 31 55 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.202
r125 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r126 28 54 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.202
r127 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r128 25 53 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=1.202
r129 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=0.56
r130 22 49 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=1.202
r131 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=0.56
r132 19 48 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.202
r133 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r134 16 47 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.202
r135 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r136 13 46 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=1.202
r137 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=0.56
r138 10 42 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r139 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r140 7 41 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=1.202
r141 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=0.56
r142 4 40 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r143 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r144 1 39 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r145 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_6%VPWR 1 2 3 4 5 6 7 22 24 30 32 36 38 42 44
+ 48 50 54 58 63 64 65 67 77 78 84 87 90 93 96
r90 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r91 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r92 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r93 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r94 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r95 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r96 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r97 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r98 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r99 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r100 75 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r101 75 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=4.83 $Y2=2.72
r102 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r103 72 96 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.095 $Y=2.72
+ $X2=4.96 $Y2=2.72
r104 72 74 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.095 $Y=2.72
+ $X2=5.75 $Y2=2.72
r105 71 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r106 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r107 68 81 4.1687 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r108 68 70 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r109 67 84 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.2 $Y2=2.72
r110 67 70 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 65 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r112 65 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r113 63 74 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=5.75 $Y2=2.72
r114 63 64 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=5.9 $Y2=2.72
r115 62 77 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.035 $Y=2.72
+ $X2=6.21 $Y2=2.72
r116 62 64 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.035 $Y=2.72
+ $X2=5.9 $Y2=2.72
r117 58 61 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.9 $Y=1.66 $X2=5.9
+ $Y2=2.34
r118 56 64 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2.72
r119 56 61 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2.34
r120 52 96 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2.72
r121 52 54 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2
r122 51 93 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.02 $Y2=2.72
r123 50 96 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=4.96 $Y2=2.72
r124 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=4.155 $Y2=2.72
r125 46 93 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r126 46 48 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2
r127 45 90 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.08 $Y2=2.72
r128 44 93 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=4.02 $Y2=2.72
r129 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=3.215 $Y2=2.72
r130 40 90 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r131 40 42 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r132 39 87 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.14 $Y2=2.72
r133 38 90 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=3.08 $Y2=2.72
r134 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.275 $Y2=2.72
r135 34 87 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r136 34 36 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r137 33 84 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.2 $Y2=2.72
r138 32 87 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.14 $Y2=2.72
r139 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=1.335 $Y2=2.72
r140 28 84 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r141 28 30 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r142 24 27 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r143 22 81 3.116 $w=2.7e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.197 $Y2=2.72
r144 22 27 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r145 7 61 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=2.34
r146 7 58 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=1.66
r147 6 54 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=2
r148 5 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2
r149 4 42 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r150 3 36 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r151 2 30 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r152 1 27 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r153 1 24 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_6%Y 1 2 3 4 5 6 7 8 9 28 30 32 36 38 42 44
+ 48 50 54 58 60 64 66 67 69 75 77 78 83 85 87 90 91
r135 81 91 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=3.485 $Y=1.495
+ $X2=3.485 $Y2=1.19
r136 81 83 1.40534 $w=3e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.485 $Y=1.495
+ $X2=3.525 $Y2=1.58
r137 78 91 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=3.485 $Y=0.885
+ $X2=3.485 $Y2=1.19
r138 78 80 3.13183 $w=3e-07 $l=1.25e-07 $layer=LI1_cond $X=3.485 $Y=0.885
+ $X2=3.485 $Y2=0.76
r139 69 87 3.14896 $w=3e-07 $l=9.88686e-08 $layer=LI1_cond $X=5.46 $Y=1.495
+ $X2=5.43 $Y2=1.58
r140 68 90 5.16603 $w=2.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.46 $Y=1.325
+ $X2=5.46 $Y2=1.19
r141 68 69 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.46 $Y=1.325
+ $X2=5.46 $Y2=1.495
r142 67 90 5.16603 $w=2.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.46 $Y=1.055
+ $X2=5.46 $Y2=1.19
r143 66 89 3.28347 $w=2.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.46 $Y=0.885
+ $X2=5.46 $Y2=0.76
r144 66 67 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.46 $Y=0.885
+ $X2=5.46 $Y2=1.055
r145 62 87 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=1.665 $X2=5.43
+ $Y2=1.58
r146 62 64 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.43 $Y=1.665
+ $X2=5.43 $Y2=2.34
r147 61 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.655 $Y=1.58
+ $X2=4.49 $Y2=1.58
r148 60 87 3.44808 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=1.58
+ $X2=5.43 $Y2=1.58
r149 60 61 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.265 $Y=1.58
+ $X2=4.655 $Y2=1.58
r150 56 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=1.665
+ $X2=4.49 $Y2=1.58
r151 56 58 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.49 $Y=1.665
+ $X2=4.49 $Y2=2.34
r152 55 83 5.10667 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=1.58
+ $X2=3.525 $Y2=1.58
r153 54 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=1.58
+ $X2=4.49 $Y2=1.58
r154 54 55 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.325 $Y=1.58
+ $X2=3.715 $Y2=1.58
r155 51 80 3.75819 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=3.635 $Y=0.76
+ $X2=3.485 $Y2=0.76
r156 51 53 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=3.635 $Y=0.76
+ $X2=4.49 $Y2=0.76
r157 50 89 3.54615 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=5.325 $Y=0.76
+ $X2=5.46 $Y2=0.76
r158 50 53 38.4916 $w=2.48e-07 $l=8.35e-07 $layer=LI1_cond $X=5.325 $Y=0.76
+ $X2=4.49 $Y2=0.76
r159 46 83 1.40534 $w=3.3e-07 $l=9.66954e-08 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.525 $Y2=1.58
r160 46 48 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=2.34
r161 45 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=1.58
+ $X2=2.61 $Y2=1.58
r162 44 83 5.10667 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=1.58
+ $X2=3.525 $Y2=1.58
r163 44 45 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.335 $Y=1.58
+ $X2=2.775 $Y2=1.58
r164 40 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.58
r165 40 42 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=2.34
r166 39 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.67 $Y2=1.58
r167 38 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=2.61 $Y2=1.58
r168 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=1.835 $Y2=1.58
r169 34 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.58
r170 34 36 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=2.34
r171 33 73 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.73 $Y2=1.58
r172 32 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=1.67 $Y2=1.58
r173 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=0.895 $Y2=1.58
r174 28 73 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.58
r175 28 30 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.34
r176 9 87 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.66
r177 9 64 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.34
r178 8 85 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.66
r179 8 58 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2.34
r180 7 83 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.66
r181 7 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.34
r182 6 77 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r183 6 42 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r184 5 75 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r185 5 36 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r186 4 73 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r187 4 30 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r188 3 89 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=5.245
+ $Y=0.235 $X2=5.43 $Y2=0.72
r189 2 53 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.72
r190 1 80 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_6%A_27_47# 1 2 3 4 5 6 7 24 26 27 30 32 36
+ 38 40 41 42 50 51 57
r96 45 47 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=4.02 $Y=0.36 $X2=4.96
+ $Y2=0.36
r97 43 53 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.165 $Y=0.36
+ $X2=3.04 $Y2=0.36
r98 43 45 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=3.165 $Y=0.36
+ $X2=4.02 $Y2=0.36
r99 42 57 4.17428 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=5.765 $Y=0.36
+ $X2=5.915 $Y2=0.36
r100 42 47 42.5152 $w=2.08e-07 $l=8.05e-07 $layer=LI1_cond $X=5.765 $Y=0.36
+ $X2=4.96 $Y2=0.36
r101 41 55 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=0.715
+ $X2=3.04 $Y2=0.8
r102 40 53 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.04 $Y=0.465
+ $X2=3.04 $Y2=0.36
r103 40 41 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=3.04 $Y=0.465
+ $X2=3.04 $Y2=0.715
r104 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.8
+ $X2=2.14 $Y2=0.8
r105 38 55 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.915 $Y=0.8
+ $X2=3.04 $Y2=0.8
r106 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=0.8
+ $X2=2.305 $Y2=0.8
r107 34 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.715
+ $X2=2.14 $Y2=0.8
r108 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.14 $Y=0.715
+ $X2=2.14 $Y2=0.38
r109 33 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0.8
+ $X2=1.2 $Y2=0.8
r110 32 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0.8
+ $X2=2.14 $Y2=0.8
r111 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.975 $Y=0.8
+ $X2=1.365 $Y2=0.8
r112 28 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.715 $X2=1.2
+ $Y2=0.8
r113 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.2 $Y=0.715
+ $X2=1.2 $Y2=0.38
r114 26 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0.8
+ $X2=1.2 $Y2=0.8
r115 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.035 $Y=0.8
+ $X2=0.425 $Y2=0.8
r116 22 27 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.425 $Y2=0.8
r117 22 24 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.257 $Y2=0.38
r118 7 57 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.765
+ $Y=0.235 $X2=5.9 $Y2=0.38
r119 6 47 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.235 $X2=4.96 $Y2=0.38
r120 5 45 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.38
r121 4 55 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.72
r122 4 53 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.38
r123 3 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r124 2 30 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r125 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_6%VGND 1 2 3 12 14 18 20 24 26 28 38 39 42
+ 45 48
r78 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r79 46 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r80 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r81 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r82 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r83 38 39 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r84 36 39 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=6.21
+ $Y2=0
r85 36 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r86 35 38 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=6.21
+ $Y2=0
r87 35 36 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r88 33 48 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.61
+ $Y2=0
r89 33 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.99
+ $Y2=0
r90 28 42 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.73
+ $Y2=0
r91 28 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r92 26 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r93 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r94 22 48 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r95 22 24 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.38
r96 21 45 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.67
+ $Y2=0
r97 20 48 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.61
+ $Y2=0
r98 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=1.805
+ $Y2=0
r99 16 45 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r100 16 18 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.38
r101 15 42 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.73
+ $Y2=0
r102 14 45 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.67
+ $Y2=0
r103 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=0.865 $Y2=0
r104 10 42 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r105 10 12 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r106 3 24 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.38
r107 2 18 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.38
r108 1 12 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

