* NGSPICE file created from sky130_fd_sc_hdll__nor3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nor3b_2 A B C_N VGND VNB VPB VPWR Y
M1000 Y a_571_21# a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u
M1001 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=4.034e+11p pd=3.96e+06u as=8.7e+11p ps=7.74e+06u
M1002 VGND C_N a_571_21# VNB nshort w=420000u l=150000u
+  ad=1.0662e+12p pd=1.084e+07u as=1.092e+11p ps=1.36e+06u
M1003 a_27_297# B a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_309_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_571_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=6.89e+11p ps=6.02e+06u
M1006 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_571_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR C_N a_571_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1010 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_309_297# a_571_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

