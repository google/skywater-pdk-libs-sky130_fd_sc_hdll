* File: sky130_fd_sc_hdll__nand2b_1.pex.spice
* Created: Thu Aug 27 19:13:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2B_1%A_N 1 3 4 6 7 12
c26 7 0 1.53383e-19 $X=0.235 $Y=1.19
c27 4 0 1.40223e-19 $X=0.52 $Y=0.995
r28 12 13 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r29 10 12 31.6932 $w=3.65e-07 $l=2.4e-07 $layer=POLY_cond $X=0.255 $Y=1.202
+ $X2=0.495 $Y2=1.202
r30 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r31 4 13 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r32 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.675
r33 1 12 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r34 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_1%B 1 3 4 6 7 11 13
c28 1 0 1.53383e-19 $X=1.03 $Y=1.41
r29 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.16 $X2=0.995 $Y2=1.16
r30 7 11 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=0.745 $Y=1.195
+ $X2=0.995 $Y2=1.195
r31 7 13 2.40092 $w=2.38e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.195
+ $X2=0.695 $Y2=1.195
r32 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=0.995 $Y2=1.16
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=0.56
r34 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=0.995 $Y2=1.16
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41 $X2=1.03
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_1%A_27_93# 1 2 7 9 10 12 13 15 20 23 27
c56 23 0 1.40223e-19 $X=0.26 $Y=0.69
r57 27 30 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=0.23 $Y=1.58 $X2=0.23
+ $Y2=1.66
r58 23 25 5.5488 $w=2.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.225 $Y=0.69
+ $X2=0.225 $Y2=0.82
r59 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.535
+ $Y=1.16 $X2=1.535 $Y2=1.16
r60 18 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=1.495
+ $X2=1.535 $Y2=1.16
r61 17 20 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.535 $Y=0.905
+ $X2=1.535 $Y2=1.16
r62 16 27 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.37 $Y=1.58 $X2=0.23
+ $Y2=1.58
r63 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.45 $Y=1.58
+ $X2=1.535 $Y2=1.495
r64 15 16 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=1.45 $Y=1.58
+ $X2=0.37 $Y2=1.58
r65 14 25 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.36 $Y=0.82
+ $X2=0.225 $Y2=0.82
r66 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.45 $Y=0.82
+ $X2=1.535 $Y2=0.905
r67 13 14 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=1.45 $Y=0.82
+ $X2=0.36 $Y2=0.82
r68 10 21 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.535 $Y2=1.16
r69 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.5 $Y=1.41 $X2=1.5
+ $Y2=1.985
r70 7 21 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.535 $Y2=1.16
r71 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=0.56
r72 2 30 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r73 1 23 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_1%VPWR 1 2 11 15 18 19 20 27 28 31 34
r33 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r34 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r35 25 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r36 25 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r37 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r38 22 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.88 $Y=2.72
+ $X2=0.755 $Y2=2.72
r39 22 24 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=0.88 $Y=2.72
+ $X2=1.61 $Y2=2.72
r40 20 32 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 20 34 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r42 18 24 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.65 $Y=2.72 $X2=1.61
+ $Y2=2.72
r43 18 19 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.65 $Y=2.72
+ $X2=1.757 $Y2=2.72
r44 17 27 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.865 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 17 19 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.865 $Y=2.72
+ $X2=1.757 $Y2=2.72
r46 13 19 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.757 $Y=2.635
+ $X2=1.757 $Y2=2.72
r47 13 15 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=1.757 $Y=2.635
+ $X2=1.757 $Y2=2.34
r48 9 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=2.635
+ $X2=0.755 $Y2=2.72
r49 9 11 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.755 $Y=2.635
+ $X2=0.755 $Y2=2
r50 2 15 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.485 $X2=1.735 $Y2=2.34
r51 1 11 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.795 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_1%Y 1 2 9 12 15 16 17 18 19 20 28 29
r37 20 29 2.55307 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=1.92
+ $X2=2.005 $Y2=1.835
r38 20 29 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.005 $Y=1.81
+ $X2=2.005 $Y2=1.835
r39 19 20 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.005 $Y=1.53
+ $X2=2.005 $Y2=1.81
r40 18 19 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.005 $Y=1.19
+ $X2=2.005 $Y2=1.53
r41 17 18 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.005 $Y=0.85
+ $X2=2.005 $Y2=1.19
r42 16 28 3.05272 $w=3.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.005 $Y=0.4
+ $X2=2.005 $Y2=0.545
r43 16 17 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.005 $Y=0.57
+ $X2=2.005 $Y2=0.85
r44 16 28 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.005 $Y=0.57
+ $X2=2.005 $Y2=0.545
r45 13 15 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.43 $Y=1.92 $X2=1.24
+ $Y2=1.92
r46 12 20 5.55669 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.82 $Y=1.92
+ $X2=2.005 $Y2=1.92
r47 12 13 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.82 $Y=1.92
+ $X2=1.43 $Y2=1.92
r48 9 16 3.89485 $w=2.9e-07 $l=1.85e-07 $layer=LI1_cond $X=1.82 $Y=0.4 $X2=2.005
+ $Y2=0.4
r49 9 11 3.57586 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.82 $Y=0.4 $X2=1.735
+ $Y2=0.4
r50 2 15 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=2
r51 1 11 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.235 $X2=1.735 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_1%VGND 1 8 10 17 18 21 24
r25 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r26 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r27 15 18 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r28 15 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r29 14 17 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r30 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r31 12 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.795
+ $Y2=0
r32 12 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.15
+ $Y2=0
r33 10 22 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r34 10 24 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r35 6 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r36 6 8 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.38
r37 1 8 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.465 $X2=0.795 $Y2=0.38
.ends

