* NGSPICE file created from sky130_fd_sc_hdll__sdfstp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 VPWR SET_B a_1229_21# VPB phighvt w=420000u l=180000u
+  ad=2.0718e+12p pd=1.868e+07u as=1.722e+11p ps=1.66e+06u
M1001 VGND a_349_21# a_295_47# VNB nshort w=420000u l=150000u
+  ad=1.50395e+12p pd=1.505e+07u as=1.134e+11p ps=1.38e+06u
M1002 a_2067_47# a_1951_295# a_1995_47# VNB nshort w=420000u l=150000u
+  ad=2.016e+11p pd=1.8e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_1745_329# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=4.746e+11p pd=4.26e+06u as=0p ps=0u
M1004 a_1951_295# a_1745_329# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1005 a_1995_47# a_693_369# a_1745_329# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.332e+11p ps=2.5e+06u
M1006 a_1891_413# a_877_369# a_1745_329# VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1007 VGND SCE a_349_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1008 a_1075_413# a_877_369# a_201_47# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.99e+11p ps=3.24e+06u
M1009 VPWR SCD a_27_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=3.456e+11p ps=3.64e+06u
M1010 a_1229_21# a_1075_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR SCE a_349_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1012 VGND SET_B a_2067_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_2447_47# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1014 VGND SET_B a_1467_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1015 a_877_369# a_693_369# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1016 VGND a_1229_21# a_1177_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1017 VPWR a_1951_295# a_1891_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND CLK a_693_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1019 a_1951_295# a_1745_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1020 a_1654_47# a_1075_413# VGND VNB nshort w=640000u l=150000u
+  ad=5.088e+11p pd=2.87e+06u as=0p ps=0u
M1021 a_1467_47# a_1075_413# a_1229_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.512e+11p ps=1.56e+06u
M1022 Q a_2447_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_369# a_349_21# a_201_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_119_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1025 a_1177_47# a_877_369# a_1075_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1026 VGND a_1745_329# a_2447_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1027 a_877_369# a_693_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1028 a_1663_329# a_1075_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=1.932e+11p pd=2.14e+06u as=0p ps=0u
M1029 VPWR a_1745_329# a_2447_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1030 a_1075_413# a_693_369# a_201_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1031 a_1745_329# a_693_369# a_1663_329# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_295_47# D a_201_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_2447_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1034 a_201_47# SCE a_119_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Q a_2447_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_211_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=0p ps=0u
M1037 a_201_47# D a_211_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1169_413# a_693_369# a_1075_413# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1039 VPWR a_1229_21# a_1169_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VPWR CLK a_693_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1041 a_1745_329# a_877_369# a_1654_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

