* File: sky130_fd_sc_hdll__sdfsbp_2.spice
* Created: Thu Aug 27 19:27:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdfsbp_2.pex.spice"
.subckt sky130_fd_sc_hdll__sdfsbp_2  VNB VPB SCD SCE D CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* SCE	SCE
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1038 A_109_47# N_SCD_M1038_g N_VGND_M1038_s VNB NSHORT L=0.15 W=0.42 AD=0.063
+ AS=0.1092 PD=0.72 PS=1.36 NRD=27.132 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1028 N_A_199_47#_M1028_d N_SCE_M1028_g A_109_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.063 PD=0.75 PS=0.72 NRD=15.708 NRS=27.132 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1032 A_295_47# N_D_M1032_g N_A_199_47#_M1028_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0693 PD=0.69 PS=0.75 NRD=22.848 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_349_21#_M1000_g A_295_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1428 AS=0.0567 PD=1.52 PS=0.69 NRD=21.42 NRS=22.848 M=1 R=2.8 SA=75001.5
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_SCE_M1004_g N_A_349_21#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1218 AS=0.1176 PD=1.42 PS=1.4 NRD=7.14 NRS=4.284 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_CLK_M1017_g N_A_693_369#_M1017_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0609 AS=0.1302 PD=0.71 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1018 N_A_877_369#_M1018_d N_A_693_369#_M1018_g N_VGND_M1017_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1218 AS=0.0609 PD=1.42 PS=0.71 NRD=7.14 NRS=4.284 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_A_1075_413#_M1031_d N_A_693_369#_M1031_g N_A_199_47#_M1031_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1024 A_1177_47# N_A_877_369#_M1024_g N_A_1075_413#_M1031_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=14.28 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1219_21#_M1029_g A_1177_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0441 PD=1.46 PS=0.63 NRD=12.852 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 A_1467_47# N_A_1075_413#_M1021_g N_A_1219_21#_M1021_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1512 PD=0.63 PS=1.56 NRD=14.28 NRS=27.132 M=1 R=2.8
+ SA=75000.3 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_SET_B_M1025_g A_1467_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0981453 AS=0.0441 PD=0.847925 PS=0.63 NRD=12.852 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1010 A_1655_47# N_A_1075_413#_M1010_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.64
+ AD=0.2368 AS=0.149555 PD=1.38 PS=1.29208 NRD=59.052 NRS=19.68 M=1 R=4.26667
+ SA=75000.9 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1005 N_A_1735_329#_M1005_d N_A_877_369#_M1005_g A_1655_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.184392 AS=0.2368 PD=1.46113 PS=1.38 NRD=13.116 NRS=59.052 M=1
+ R=4.26667 SA=75001.8 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1045 A_1977_47# N_A_693_369#_M1045_g N_A_1735_329#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.121008 PD=0.63 PS=0.958868 NRD=14.28 NRS=62.856 M=1
+ R=2.8 SA=75002.8 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1039 A_2049_47# N_A_1930_295#_M1039_g A_1977_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1344 AS=0.0441 PD=1.06 PS=0.63 NRD=75.708 NRS=14.28 M=1 R=2.8 SA=75003.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1043 N_VGND_M1043_d N_SET_B_M1043_g A_2049_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.09555 AS=0.1344 PD=0.875 PS=1.06 NRD=37.14 NRS=75.708 M=1 R=2.8 SA=75004
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_A_1930_295#_M1001_d N_A_1735_329#_M1001_g N_VGND_M1043_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.09555 PD=1.36 PS=0.875 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75004.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_1735_329#_M1015_g N_Q_N_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1030 N_VGND_M1030_d N_A_1735_329#_M1030_g N_Q_N_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.24375 AS=0.104 PD=2.05 PS=0.97 NRD=20.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1033 N_VGND_M1033_d N_A_1735_329#_M1033_g N_A_2739_47#_M1033_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0889065 AS=0.1302 PD=0.804673 PS=1.46 NRD=5.712 NRS=12.852
+ M=1 R=2.8 SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 N_Q_M1006_d N_A_2739_47#_M1006_g N_VGND_M1033_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.137593 PD=0.97 PS=1.24533 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75000.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1034 N_Q_M1006_d N_A_2739_47#_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=8.304 NRS=8.304 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_SCD_M1007_g N_A_27_369#_M1007_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1036 A_211_369# N_SCE_M1036_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0736 AS=0.0928 PD=0.87 PS=0.93 NRD=18.4589 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1040 N_A_199_47#_M1040_d N_D_M1040_g A_211_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.0736 PD=0.93 PS=0.87 NRD=1.5366 NRS=18.4589 M=1 R=3.55556
+ SA=90001.1 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1022 N_A_27_369#_M1022_d N_A_349_21#_M1022_g N_A_199_47#_M1040_d VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1
+ R=3.55556 SA=90001.5 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1011 N_VPWR_M1011_d N_SCE_M1011_g N_A_349_21#_M1011_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.1728 PD=1.82 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1044 N_VPWR_M1044_d N_CLK_M1044_g N_A_693_369#_M1044_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1027 N_A_877_369#_M1027_d N_A_693_369#_M1027_g N_VPWR_M1044_d VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1
+ R=3.55556 SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1003 N_A_1075_413#_M1003_d N_A_877_369#_M1003_g N_A_199_47#_M1003_s VPB
+ PHIGHVT L=0.18 W=0.42 AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443
+ NRS=2.3443 M=1 R=2.33333 SA=90000.2 SB=90005.4 A=0.0756 P=1.2 MULT=1
MM1041 A_1169_413# N_A_693_369#_M1041_g N_A_1075_413#_M1003_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0798 AS=0.0609 PD=0.8 PS=0.71 NRD=63.3158 NRS=2.3443 M=1 R=2.33333
+ SA=90000.6 SB=90004.9 A=0.0756 P=1.2 MULT=1
MM1042 N_VPWR_M1042_d N_A_1219_21#_M1042_g A_1169_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0966 AS=0.0798 PD=0.88 PS=0.8 NRD=30.4759 NRS=63.3158 M=1 R=2.33333
+ SA=90001.2 SB=90004.4 A=0.0756 P=1.2 MULT=1
MM1008 N_A_1219_21#_M1008_d N_A_1075_413#_M1008_g N_VPWR_M1042_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.08505 AS=0.0966 PD=0.825 PS=0.88 NRD=11.7215 NRS=53.9386
+ M=1 R=2.33333 SA=90001.8 SB=90003.7 A=0.0756 P=1.2 MULT=1
MM1023 N_VPWR_M1023_d N_SET_B_M1023_g N_A_1219_21#_M1008_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0994 AS=0.08505 PD=0.86 PS=0.825 NRD=23.443 NRS=46.886 M=1
+ R=2.33333 SA=90002.4 SB=90003.1 A=0.0756 P=1.2 MULT=1
MM1035 A_1652_329# N_A_1075_413#_M1035_g N_VPWR_M1023_d VPB PHIGHVT L=0.18
+ W=0.84 AD=0.0987 AS=0.1988 PD=1.075 PS=1.72 NRD=14.6568 NRS=28.1316 M=1
+ R=4.66667 SA=90001.6 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1012 N_A_1735_329#_M1012_d N_A_693_369#_M1012_g A_1652_329# VPB PHIGHVT L=0.18
+ W=0.84 AD=0.2114 AS=0.0987 PD=1.78 PS=1.075 NRD=35.1645 NRS=14.6568 M=1
+ R=4.66667 SA=90002 SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1009 A_1870_413# N_A_877_369#_M1009_g N_A_1735_329#_M1012_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0651 AS=0.1057 PD=0.73 PS=0.89 NRD=46.886 NRS=30.4759 M=1
+ R=2.33333 SA=90004.2 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1020 N_VPWR_M1020_d N_A_1930_295#_M1020_g A_1870_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.11865 AS=0.0651 PD=0.985 PS=0.73 NRD=107.877 NRS=46.886 M=1
+ R=2.33333 SA=90004.6 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1013 N_A_1735_329#_M1013_d N_SET_B_M1013_g N_VPWR_M1020_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.11865 PD=1.38 PS=0.985 NRD=2.3443 NRS=25.7873 M=1
+ R=2.33333 SA=90005.4 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1002 N_A_1930_295#_M1002_d N_A_1735_329#_M1002_g N_VPWR_M1002_s VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1019 N_VPWR_M1019_d N_A_1735_329#_M1019_g N_Q_N_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1037 N_VPWR_M1037_d N_A_1735_329#_M1037_g N_Q_N_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.335 AS=0.145 PD=2.67 PS=1.29 NRD=13.7703 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_A_1735_329#_M1016_g N_A_2739_47#_M1016_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.122693 AS=0.1728 PD=1.04976 PS=1.82 NRD=16.9223 NRS=1.5366
+ M=1 R=3.55556 SA=90000.2 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1014 N_VPWR_M1016_d N_A_2739_47#_M1014_g N_Q_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.191707 AS=0.145 PD=1.64024 PS=1.29 NRD=1.9503 NRS=0.9653 M=1 R=5.55556
+ SA=90000.5 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1026 N_VPWR_M1026_d N_A_2739_47#_M1026_g N_Q_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.32 AS=0.145 PD=2.64 PS=1.29 NRD=10.8153 NRS=0.9653 M=1 R=5.55556 SA=90001
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX46_noxref VNB VPB NWDIODE A=25.7121 P=35.25
c_133 VNB 0 1.07953e-19 $X=0.15 $Y=-0.085
c_293 VPB 0 1.93782e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__sdfsbp_2.pxi.spice"
*
.ends
*
*
