* File: sky130_fd_sc_hdll__muxb4to1_4.pxi.spice
* Created: Wed Sep  2 08:35:52 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[0] N_D[0]_M1003_g N_D[0]_M1024_g
+ N_D[0]_M1057_g N_D[0]_M1041_g N_D[0]_M1055_g N_D[0]_M1073_g N_D[0]_M1078_g
+ N_D[0]_M1071_g D[0] N_D[0]_c_494_n N_D[0]_c_495_n N_D[0]_c_496_n
+ N_D[0]_c_497_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[0]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_559_265# N_A_559_265#_M1046_d
+ N_A_559_265#_M1004_s N_A_559_265#_c_576_n N_A_559_265#_M1042_g
+ N_A_559_265#_c_577_n N_A_559_265#_c_578_n N_A_559_265#_c_579_n
+ N_A_559_265#_M1056_g N_A_559_265#_c_580_n N_A_559_265#_c_581_n
+ N_A_559_265#_M1063_g N_A_559_265#_c_582_n N_A_559_265#_c_583_n
+ N_A_559_265#_M1072_g N_A_559_265#_c_584_n N_A_559_265#_c_585_n
+ N_A_559_265#_c_569_n N_A_559_265#_c_570_n N_A_559_265#_c_571_n
+ N_A_559_265#_c_572_n N_A_559_265#_c_588_n N_A_559_265#_c_573_n
+ N_A_559_265#_c_574_n N_A_559_265#_c_590_n N_A_559_265#_c_575_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_559_265#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[0] N_S[0]_c_686_n N_S[0]_M1015_g
+ N_S[0]_c_687_n N_S[0]_c_688_n N_S[0]_c_689_n N_S[0]_M1023_g N_S[0]_c_690_n
+ N_S[0]_c_691_n N_S[0]_M1028_g N_S[0]_c_692_n N_S[0]_c_693_n N_S[0]_M1037_g
+ N_S[0]_c_694_n N_S[0]_c_695_n N_S[0]_c_696_n N_S[0]_c_697_n N_S[0]_c_698_n
+ N_S[0]_c_709_n N_S[0]_M1004_g N_S[0]_c_699_n N_S[0]_M1046_g N_S[0]_c_700_n
+ N_S[0]_c_701_n N_S[0]_M1053_g N_S[0]_c_702_n N_S[0]_M1018_g N_S[0]_c_703_n
+ N_S[0]_c_704_n N_S[0]_c_705_n N_S[0]_c_706_n S[0]
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[0]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[1] N_S[1]_c_801_n N_S[1]_c_802_n
+ N_S[1]_M1036_g N_S[1]_c_803_n N_S[1]_M1061_g N_S[1]_c_804_n N_S[1]_c_805_n
+ N_S[1]_M1069_g N_S[1]_c_806_n N_S[1]_c_826_n N_S[1]_M1050_g N_S[1]_c_807_n
+ N_S[1]_c_808_n N_S[1]_c_809_n N_S[1]_c_810_n N_S[1]_c_811_n N_S[1]_M1007_g
+ N_S[1]_c_812_n N_S[1]_c_813_n N_S[1]_M1016_g N_S[1]_c_814_n N_S[1]_c_815_n
+ N_S[1]_M1026_g N_S[1]_c_816_n N_S[1]_c_817_n N_S[1]_M1033_g N_S[1]_c_818_n
+ N_S[1]_c_819_n N_S[1]_c_820_n N_S[1]_c_821_n S[1] N_S[1]_c_822_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[1]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_1430_325# N_A_1430_325#_M1061_s
+ N_A_1430_325#_M1036_s N_A_1430_325#_c_926_n N_A_1430_325#_M1000_g
+ N_A_1430_325#_c_927_n N_A_1430_325#_c_919_n N_A_1430_325#_c_929_n
+ N_A_1430_325#_M1014_g N_A_1430_325#_c_930_n N_A_1430_325#_c_931_n
+ N_A_1430_325#_M1043_g N_A_1430_325#_c_932_n N_A_1430_325#_c_933_n
+ N_A_1430_325#_M1066_g N_A_1430_325#_c_934_n N_A_1430_325#_c_935_n
+ N_A_1430_325#_c_936_n N_A_1430_325#_c_920_n N_A_1430_325#_c_921_n
+ N_A_1430_325#_c_922_n N_A_1430_325#_c_938_n N_A_1430_325#_c_923_n
+ N_A_1430_325#_c_924_n N_A_1430_325#_c_925_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_1430_325#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[1] N_D[1]_M1001_g N_D[1]_M1017_g
+ N_D[1]_M1029_g N_D[1]_M1006_g N_D[1]_M1038_g N_D[1]_M1049_g N_D[1]_M1079_g
+ N_D[1]_M1065_g D[1] N_D[1]_c_1043_n N_D[1]_c_1044_n N_D[1]_c_1045_n
+ N_D[1]_c_1046_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[1]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[2] N_D[2]_M1005_g N_D[2]_M1002_g
+ N_D[2]_M1021_g N_D[2]_M1019_g N_D[2]_M1047_g N_D[2]_M1034_g N_D[2]_M1052_g
+ N_D[2]_M1074_g D[2] N_D[2]_c_1129_n N_D[2]_c_1130_n N_D[2]_c_1131_n
+ N_D[2]_c_1132_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[2]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_3135_265# N_A_3135_265#_M1058_s
+ N_A_3135_265#_M1020_d N_A_3135_265#_c_1216_n N_A_3135_265#_M1025_g
+ N_A_3135_265#_c_1217_n N_A_3135_265#_c_1218_n N_A_3135_265#_c_1219_n
+ N_A_3135_265#_M1044_g N_A_3135_265#_c_1220_n N_A_3135_265#_c_1221_n
+ N_A_3135_265#_M1051_g N_A_3135_265#_c_1222_n N_A_3135_265#_c_1223_n
+ N_A_3135_265#_M1064_g N_A_3135_265#_c_1224_n N_A_3135_265#_c_1225_n
+ N_A_3135_265#_c_1209_n N_A_3135_265#_c_1210_n N_A_3135_265#_c_1211_n
+ N_A_3135_265#_c_1212_n N_A_3135_265#_c_1228_n N_A_3135_265#_c_1213_n
+ N_A_3135_265#_c_1214_n N_A_3135_265#_c_1230_n N_A_3135_265#_c_1215_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_3135_265#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[2] N_S[2]_c_1328_n N_S[2]_M1008_g
+ N_S[2]_c_1329_n N_S[2]_c_1330_n N_S[2]_c_1331_n N_S[2]_M1009_g N_S[2]_c_1332_n
+ N_S[2]_c_1333_n N_S[2]_M1030_g N_S[2]_c_1334_n N_S[2]_c_1335_n N_S[2]_M1077_g
+ N_S[2]_c_1336_n N_S[2]_c_1337_n N_S[2]_c_1338_n N_S[2]_c_1339_n
+ N_S[2]_c_1340_n N_S[2]_c_1351_n N_S[2]_M1020_g N_S[2]_c_1341_n N_S[2]_M1058_g
+ N_S[2]_c_1342_n N_S[2]_c_1343_n N_S[2]_M1062_g N_S[2]_c_1344_n N_S[2]_M1076_g
+ N_S[2]_c_1345_n N_S[2]_c_1346_n N_S[2]_c_1347_n N_S[2]_c_1348_n S[2]
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[2]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[3] N_S[3]_c_1443_n N_S[3]_c_1444_n
+ N_S[3]_M1045_g N_S[3]_c_1445_n N_S[3]_M1059_g N_S[3]_c_1446_n N_S[3]_c_1447_n
+ N_S[3]_M1075_g N_S[3]_c_1448_n N_S[3]_c_1468_n N_S[3]_M1067_g N_S[3]_c_1449_n
+ N_S[3]_c_1450_n N_S[3]_c_1451_n N_S[3]_c_1452_n N_S[3]_c_1453_n N_S[3]_M1011_g
+ N_S[3]_c_1454_n N_S[3]_c_1455_n N_S[3]_M1012_g N_S[3]_c_1456_n N_S[3]_c_1457_n
+ N_S[3]_M1022_g N_S[3]_c_1458_n N_S[3]_c_1459_n N_S[3]_M1031_g N_S[3]_c_1460_n
+ N_S[3]_c_1461_n N_S[3]_c_1462_n N_S[3]_c_1463_n S[3] N_S[3]_c_1464_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[3]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_4006_325# N_A_4006_325#_M1059_s
+ N_A_4006_325#_M1045_d N_A_4006_325#_c_1568_n N_A_4006_325#_M1039_g
+ N_A_4006_325#_c_1569_n N_A_4006_325#_c_1561_n N_A_4006_325#_c_1571_n
+ N_A_4006_325#_M1048_g N_A_4006_325#_c_1572_n N_A_4006_325#_c_1573_n
+ N_A_4006_325#_M1060_g N_A_4006_325#_c_1574_n N_A_4006_325#_c_1575_n
+ N_A_4006_325#_M1068_g N_A_4006_325#_c_1576_n N_A_4006_325#_c_1577_n
+ N_A_4006_325#_c_1578_n N_A_4006_325#_c_1562_n N_A_4006_325#_c_1563_n
+ N_A_4006_325#_c_1564_n N_A_4006_325#_c_1580_n N_A_4006_325#_c_1565_n
+ N_A_4006_325#_c_1566_n N_A_4006_325#_c_1567_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_4006_325#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[3] N_D[3]_M1010_g N_D[3]_M1013_g
+ N_D[3]_M1032_g N_D[3]_M1027_g N_D[3]_M1035_g N_D[3]_M1040_g N_D[3]_M1054_g
+ N_D[3]_M1070_g D[3] N_D[3]_c_1683_n N_D[3]_c_1684_n N_D[3]_c_1685_n
+ N_D[3]_c_1686_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[3]
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%VPWR N_VPWR_M1003_d N_VPWR_M1041_d
+ N_VPWR_M1071_d N_VPWR_M1004_d N_VPWR_M1018_d N_VPWR_M1036_d N_VPWR_M1050_d
+ N_VPWR_M1001_s N_VPWR_M1006_s N_VPWR_M1065_s N_VPWR_M1005_s N_VPWR_M1019_s
+ N_VPWR_M1074_s N_VPWR_M1020_s N_VPWR_M1076_s N_VPWR_M1045_s N_VPWR_M1067_s
+ N_VPWR_M1010_d N_VPWR_M1027_d N_VPWR_M1070_d N_VPWR_c_1757_n N_VPWR_c_1758_n
+ N_VPWR_c_1759_n N_VPWR_c_1760_n N_VPWR_c_1761_n N_VPWR_c_1762_n
+ N_VPWR_c_1763_n N_VPWR_c_1764_n N_VPWR_c_1765_n N_VPWR_c_1766_n
+ N_VPWR_c_1767_n N_VPWR_c_1768_n N_VPWR_c_1769_n N_VPWR_c_1770_n
+ N_VPWR_c_1771_n N_VPWR_c_1772_n N_VPWR_c_1773_n N_VPWR_c_1774_n
+ N_VPWR_c_1775_n N_VPWR_c_1776_n N_VPWR_c_1777_n N_VPWR_c_1778_n
+ N_VPWR_c_1779_n N_VPWR_c_1780_n N_VPWR_c_1781_n N_VPWR_c_1782_n
+ N_VPWR_c_1783_n N_VPWR_c_1784_n N_VPWR_c_1785_n N_VPWR_c_1786_n
+ N_VPWR_c_1787_n N_VPWR_c_1788_n N_VPWR_c_1789_n N_VPWR_c_1790_n
+ N_VPWR_c_1791_n N_VPWR_c_1792_n N_VPWR_c_1793_n N_VPWR_c_1794_n
+ N_VPWR_c_1795_n N_VPWR_c_1796_n N_VPWR_c_1797_n N_VPWR_c_1798_n
+ N_VPWR_c_1799_n VPWR VPWR VPWR VPWR N_VPWR_c_1801_n N_VPWR_c_1802_n
+ N_VPWR_c_1803_n N_VPWR_c_1804_n N_VPWR_c_1805_n N_VPWR_c_1806_n
+ N_VPWR_c_1807_n N_VPWR_c_1808_n N_VPWR_c_1809_n N_VPWR_c_1810_n
+ N_VPWR_c_1811_n N_VPWR_c_1812_n N_VPWR_c_1813_n N_VPWR_c_1814_n
+ N_VPWR_c_1815_n N_VPWR_c_1816_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%VPWR
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_117_297# N_A_117_297#_M1003_s
+ N_A_117_297#_M1055_s N_A_117_297#_M1042_d N_A_117_297#_M1056_d
+ N_A_117_297#_M1072_d N_A_117_297#_c_2110_n N_A_117_297#_c_2114_n
+ N_A_117_297#_c_2117_n N_A_117_297#_c_2121_n N_A_117_297#_c_2102_n
+ N_A_117_297#_c_2103_n N_A_117_297#_c_2104_n N_A_117_297#_c_2105_n
+ N_A_117_297#_c_2106_n N_A_117_297#_c_2107_n N_A_117_297#_c_2108_n
+ N_A_117_297#_c_2126_n N_A_117_297#_c_2109_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_117_297#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%Z N_Z_M1015_s N_Z_M1028_s N_Z_M1007_d
+ N_Z_M1026_d N_Z_M1008_d N_Z_M1030_d N_Z_M1011_d N_Z_M1022_d N_Z_M1042_s
+ N_Z_M1063_s N_Z_M1000_d N_Z_M1043_d N_Z_M1025_s N_Z_M1051_s N_Z_M1039_s
+ N_Z_M1060_s N_Z_c_2191_n N_Z_c_2192_n N_Z_c_2193_n N_Z_c_2194_n N_Z_c_2195_n
+ N_Z_c_2196_n N_Z_c_2197_n N_Z_c_2198_n N_Z_c_2199_n N_Z_c_2200_n N_Z_c_2201_n
+ N_Z_c_2202_n N_Z_c_2203_n N_Z_c_2204_n N_Z_c_2205_n N_Z_c_2206_n N_Z_c_2207_n
+ N_Z_c_2208_n N_Z_c_2209_n N_Z_c_2210_n N_Z_c_2211_n N_Z_c_2212_n N_Z_c_2213_n
+ N_Z_c_2214_n N_Z_c_2219_n N_Z_c_2421_n N_Z_c_2220_n N_Z_c_2435_n N_Z_c_2221_n
+ N_Z_c_2445_n N_Z_c_2298_n N_Z_c_2447_n N_Z_c_2398_n N_Z_c_2449_n Z Z Z Z Z
+ N_Z_c_2239_n N_Z_c_2245_n N_Z_c_2300_n N_Z_c_2307_n N_Z_c_2340_n N_Z_c_2346_n
+ N_Z_c_2400_n N_Z_c_2407_n N_Z_c_2454_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%Z
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_1643_311# N_A_1643_311#_M1000_s
+ N_A_1643_311#_M1014_s N_A_1643_311#_M1066_s N_A_1643_311#_M1001_d
+ N_A_1643_311#_M1038_d N_A_1643_311#_c_2607_n N_A_1643_311#_c_2608_n
+ N_A_1643_311#_c_2609_n N_A_1643_311#_c_2610_n N_A_1643_311#_c_2611_n
+ N_A_1643_311#_c_2612_n N_A_1643_311#_c_2613_n N_A_1643_311#_c_2614_n
+ N_A_1643_311#_c_2633_n N_A_1643_311#_c_2636_n N_A_1643_311#_c_2640_n
+ N_A_1643_311#_c_2644_n N_A_1643_311#_c_2615_n N_A_1643_311#_c_2647_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_1643_311#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_2693_297# N_A_2693_297#_M1005_d
+ N_A_2693_297#_M1047_d N_A_2693_297#_M1025_d N_A_2693_297#_M1044_d
+ N_A_2693_297#_M1064_d N_A_2693_297#_c_2720_n N_A_2693_297#_c_2724_n
+ N_A_2693_297#_c_2727_n N_A_2693_297#_c_2731_n N_A_2693_297#_c_2712_n
+ N_A_2693_297#_c_2713_n N_A_2693_297#_c_2714_n N_A_2693_297#_c_2715_n
+ N_A_2693_297#_c_2716_n N_A_2693_297#_c_2717_n N_A_2693_297#_c_2718_n
+ N_A_2693_297#_c_2736_n N_A_2693_297#_c_2719_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_2693_297#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_4219_311# N_A_4219_311#_M1039_d
+ N_A_4219_311#_M1048_d N_A_4219_311#_M1068_d N_A_4219_311#_M1010_s
+ N_A_4219_311#_M1035_s N_A_4219_311#_c_2814_n N_A_4219_311#_c_2815_n
+ N_A_4219_311#_c_2816_n N_A_4219_311#_c_2817_n N_A_4219_311#_c_2818_n
+ N_A_4219_311#_c_2819_n N_A_4219_311#_c_2820_n N_A_4219_311#_c_2821_n
+ N_A_4219_311#_c_2839_n N_A_4219_311#_c_2842_n N_A_4219_311#_c_2846_n
+ N_A_4219_311#_c_2850_n N_A_4219_311#_c_2822_n N_A_4219_311#_c_2853_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_4219_311#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%VGND N_VGND_M1024_d N_VGND_M1057_d
+ N_VGND_M1078_d N_VGND_M1046_s N_VGND_M1053_s N_VGND_M1061_d N_VGND_M1069_d
+ N_VGND_M1017_d N_VGND_M1029_d N_VGND_M1079_d N_VGND_M1002_s N_VGND_M1021_s
+ N_VGND_M1052_s N_VGND_M1058_d N_VGND_M1062_d N_VGND_M1059_d N_VGND_M1075_d
+ N_VGND_M1013_d N_VGND_M1032_d N_VGND_M1054_d N_VGND_c_2906_n N_VGND_c_2907_n
+ N_VGND_c_2908_n N_VGND_c_2909_n N_VGND_c_2910_n N_VGND_c_2911_n
+ N_VGND_c_2912_n N_VGND_c_2913_n N_VGND_c_2914_n N_VGND_c_2915_n
+ N_VGND_c_2916_n N_VGND_c_2917_n N_VGND_c_2918_n N_VGND_c_2919_n
+ N_VGND_c_2920_n N_VGND_c_2921_n N_VGND_c_2922_n N_VGND_c_2923_n
+ N_VGND_c_2924_n N_VGND_c_2925_n N_VGND_c_2926_n N_VGND_c_2927_n
+ N_VGND_c_2928_n N_VGND_c_2929_n N_VGND_c_2930_n N_VGND_c_2931_n
+ N_VGND_c_2932_n N_VGND_c_2933_n N_VGND_c_2934_n N_VGND_c_2935_n
+ N_VGND_c_2936_n N_VGND_c_2937_n N_VGND_c_2938_n N_VGND_c_2939_n
+ N_VGND_c_2940_n N_VGND_c_2941_n N_VGND_c_2942_n N_VGND_c_2943_n
+ N_VGND_c_2944_n N_VGND_c_2945_n N_VGND_c_2946_n N_VGND_c_2947_n
+ N_VGND_c_2948_n N_VGND_c_2949_n N_VGND_c_2950_n VGND VGND VGND VGND
+ N_VGND_c_2952_n N_VGND_c_2953_n N_VGND_c_2954_n N_VGND_c_2955_n
+ N_VGND_c_2956_n N_VGND_c_2957_n N_VGND_c_2958_n N_VGND_c_2959_n
+ N_VGND_c_2960_n N_VGND_c_2961_n N_VGND_c_2962_n N_VGND_c_2963_n
+ N_VGND_c_2964_n N_VGND_c_2965_n PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%VGND
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_119_47# N_A_119_47#_M1024_s
+ N_A_119_47#_M1073_s N_A_119_47#_M1015_d N_A_119_47#_M1023_d
+ N_A_119_47#_M1037_d N_A_119_47#_c_3254_n N_A_119_47#_c_3257_n
+ N_A_119_47#_c_3246_n N_A_119_47#_c_3265_n N_A_119_47#_c_3247_n
+ N_A_119_47#_c_3248_n N_A_119_47#_c_3249_n N_A_119_47#_c_3250_n
+ N_A_119_47#_c_3274_n N_A_119_47#_c_3251_n N_A_119_47#_c_3252_n
+ N_A_119_47#_c_3253_n N_A_119_47#_c_3287_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_119_47#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_1693_66# N_A_1693_66#_M1007_s
+ N_A_1693_66#_M1016_s N_A_1693_66#_M1033_s N_A_1693_66#_M1017_s
+ N_A_1693_66#_M1049_s N_A_1693_66#_c_3329_n N_A_1693_66#_c_3330_n
+ N_A_1693_66#_c_3331_n N_A_1693_66#_c_3351_n N_A_1693_66#_c_3332_n
+ N_A_1693_66#_c_3333_n N_A_1693_66#_c_3334_n N_A_1693_66#_c_3335_n
+ N_A_1693_66#_c_3354_n N_A_1693_66#_c_3336_n N_A_1693_66#_c_3363_n
+ N_A_1693_66#_c_3348_n N_A_1693_66#_c_3337_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_1693_66#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_2695_47# N_A_2695_47#_M1002_d
+ N_A_2695_47#_M1034_d N_A_2695_47#_M1008_s N_A_2695_47#_M1009_s
+ N_A_2695_47#_M1077_s N_A_2695_47#_c_3421_n N_A_2695_47#_c_3424_n
+ N_A_2695_47#_c_3413_n N_A_2695_47#_c_3432_n N_A_2695_47#_c_3414_n
+ N_A_2695_47#_c_3415_n N_A_2695_47#_c_3416_n N_A_2695_47#_c_3417_n
+ N_A_2695_47#_c_3441_n N_A_2695_47#_c_3418_n N_A_2695_47#_c_3419_n
+ N_A_2695_47#_c_3420_n N_A_2695_47#_c_3454_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_2695_47#
x_PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_4269_66# N_A_4269_66#_M1011_s
+ N_A_4269_66#_M1012_s N_A_4269_66#_M1031_s N_A_4269_66#_M1013_s
+ N_A_4269_66#_M1040_s N_A_4269_66#_c_3496_n N_A_4269_66#_c_3497_n
+ N_A_4269_66#_c_3498_n N_A_4269_66#_c_3518_n N_A_4269_66#_c_3499_n
+ N_A_4269_66#_c_3500_n N_A_4269_66#_c_3501_n N_A_4269_66#_c_3502_n
+ N_A_4269_66#_c_3521_n N_A_4269_66#_c_3503_n N_A_4269_66#_c_3530_n
+ N_A_4269_66#_c_3515_n N_A_4269_66#_c_3504_n
+ PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_4269_66#
cc_1 VNB N_D[0]_M1003_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_2 VNB N_D[0]_M1024_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_3 VNB N_D[0]_M1057_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_4 VNB N_D[0]_M1041_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_5 VNB N_D[0]_M1055_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_6 VNB N_D[0]_M1073_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_7 VNB N_D[0]_M1078_g 0.024303f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_8 VNB N_D[0]_M1071_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_9 VNB N_D[0]_c_494_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.16
cc_10 VNB N_D[0]_c_495_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.16
cc_11 VNB N_D[0]_c_496_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_12 VNB N_D[0]_c_497_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_13 VNB N_A_559_265#_c_569_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_14 VNB N_A_559_265#_c_570_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_559_265#_c_571_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_16 VNB N_A_559_265#_c_572_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_17 VNB N_A_559_265#_c_573_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.16
cc_18 VNB N_A_559_265#_c_574_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.16
cc_19 VNB N_A_559_265#_c_575_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_20 VNB N_S[0]_c_686_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_21 VNB N_S[0]_c_687_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_S[0]_c_688_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_23 VNB N_S[0]_c_689_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_24 VNB N_S[0]_c_690_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_25 VNB N_S[0]_c_691_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_26 VNB N_S[0]_c_692_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_27 VNB N_S[0]_c_693_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_S[0]_c_694_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_29 VNB N_S[0]_c_695_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_30 VNB N_S[0]_c_696_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_31 VNB N_S[0]_c_697_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_S[0]_c_698_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_33 VNB N_S[0]_c_699_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_34 VNB N_S[0]_c_700_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_35 VNB N_S[0]_c_701_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.16
cc_36 VNB N_S[0]_c_702_n 0.065295f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_37 VNB N_S[0]_c_703_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_S[0]_c_704_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_39 VNB N_S[0]_c_705_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_40 VNB N_S[0]_c_706_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_41 VNB S[0] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_42 VNB N_S[1]_c_801_n 0.032202f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_43 VNB N_S[1]_c_802_n 0.0330319f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_44 VNB N_S[1]_c_803_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_45 VNB N_S[1]_c_804_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_46 VNB N_S[1]_c_805_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_47 VNB N_S[1]_c_806_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_48 VNB N_S[1]_c_807_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_49 VNB N_S[1]_c_808_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_50 VNB N_S[1]_c_809_n 0.046608f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_51 VNB N_S[1]_c_810_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_S[1]_c_811_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.025
cc_53 VNB N_S[1]_c_812_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_S[1]_c_813_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_55 VNB N_S[1]_c_814_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_56 VNB N_S[1]_c_815_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.16
cc_57 VNB N_S[1]_c_816_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_58 VNB N_S[1]_c_817_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_59 VNB N_S[1]_c_818_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_60 VNB N_S[1]_c_819_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_61 VNB N_S[1]_c_820_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_62 VNB N_S[1]_c_821_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_63 VNB N_S[1]_c_822_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_64 VNB N_A_1430_325#_c_919_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_65 VNB N_A_1430_325#_c_920_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_66 VNB N_A_1430_325#_c_921_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.16
cc_67 VNB N_A_1430_325#_c_922_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_68 VNB N_A_1430_325#_c_923_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.16
cc_69 VNB N_A_1430_325#_c_924_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_70 VNB N_A_1430_325#_c_925_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_71 VNB N_D[1]_M1001_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_72 VNB N_D[1]_M1017_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_73 VNB N_D[1]_M1029_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_74 VNB N_D[1]_M1006_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_75 VNB N_D[1]_M1038_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_76 VNB N_D[1]_M1049_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_77 VNB N_D[1]_M1079_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_78 VNB N_D[1]_M1065_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_79 VNB N_D[1]_c_1043_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.16
cc_80 VNB N_D[1]_c_1044_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.16
cc_81 VNB N_D[1]_c_1045_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_82 VNB N_D[1]_c_1046_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_D[2]_M1005_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_84 VNB N_D[2]_M1002_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_85 VNB N_D[2]_M1021_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_86 VNB N_D[2]_M1019_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_87 VNB N_D[2]_M1047_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_88 VNB N_D[2]_M1034_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_89 VNB N_D[2]_M1052_g 0.024303f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_90 VNB N_D[2]_M1074_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_91 VNB N_D[2]_c_1129_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.16
cc_92 VNB N_D[2]_c_1130_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.16
cc_93 VNB N_D[2]_c_1131_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_94 VNB N_D[2]_c_1132_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_95 VNB N_A_3135_265#_c_1209_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_96 VNB N_A_3135_265#_c_1210_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_3135_265#_c_1211_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_98 VNB N_A_3135_265#_c_1212_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=1.16
cc_99 VNB N_A_3135_265#_c_1213_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.16
cc_100 VNB N_A_3135_265#_c_1214_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=1.46
+ $Y2=1.16
cc_101 VNB N_A_3135_265#_c_1215_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_102 VNB N_S[2]_c_1328_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_103 VNB N_S[2]_c_1329_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_S[2]_c_1330_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_105 VNB N_S[2]_c_1331_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_106 VNB N_S[2]_c_1332_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_107 VNB N_S[2]_c_1333_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_108 VNB N_S[2]_c_1334_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_109 VNB N_S[2]_c_1335_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_S[2]_c_1336_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_111 VNB N_S[2]_c_1337_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_112 VNB N_S[2]_c_1338_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_113 VNB N_S[2]_c_1339_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_S[2]_c_1340_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_115 VNB N_S[2]_c_1341_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_116 VNB N_S[2]_c_1342_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_117 VNB N_S[2]_c_1343_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.16
cc_118 VNB N_S[2]_c_1344_n 0.065295f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_119 VNB N_S[2]_c_1345_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_S[2]_c_1346_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_121 VNB N_S[2]_c_1347_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_122 VNB N_S[2]_c_1348_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_123 VNB S[2] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_124 VNB N_S[3]_c_1443_n 0.032202f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.295
cc_125 VNB N_S[3]_c_1444_n 0.0330319f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_126 VNB N_S[3]_c_1445_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_127 VNB N_S[3]_c_1446_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.025
cc_128 VNB N_S[3]_c_1447_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_129 VNB N_S[3]_c_1448_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_130 VNB N_S[3]_c_1449_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_131 VNB N_S[3]_c_1450_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_132 VNB N_S[3]_c_1451_n 0.046608f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_133 VNB N_S[3]_c_1452_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_S[3]_c_1453_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.025
cc_135 VNB N_S[3]_c_1454_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_S[3]_c_1455_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_137 VNB N_S[3]_c_1456_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_138 VNB N_S[3]_c_1457_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.16
cc_139 VNB N_S[3]_c_1458_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_140 VNB N_S[3]_c_1459_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_141 VNB N_S[3]_c_1460_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_142 VNB N_S[3]_c_1461_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_143 VNB N_S[3]_c_1462_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_144 VNB N_S[3]_c_1463_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_145 VNB N_S[3]_c_1464_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_146 VNB N_A_4006_325#_c_1561_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_147 VNB N_A_4006_325#_c_1562_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=0.605
+ $Y2=1.105
cc_148 VNB N_A_4006_325#_c_1563_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=1.055
+ $Y2=1.16
cc_149 VNB N_A_4006_325#_c_1564_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_150 VNB N_A_4006_325#_c_1565_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.16
cc_151 VNB N_A_4006_325#_c_1566_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=1.62
+ $Y2=1.16
cc_152 VNB N_A_4006_325#_c_1567_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_153 VNB N_D[3]_M1010_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_154 VNB N_D[3]_M1013_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_155 VNB N_D[3]_M1032_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_156 VNB N_D[3]_M1027_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_157 VNB N_D[3]_M1035_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_158 VNB N_D[3]_M1040_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_159 VNB N_D[3]_M1054_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_160 VNB N_D[3]_M1070_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_161 VNB N_D[3]_c_1683_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.16
cc_162 VNB N_D[3]_c_1684_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.16
cc_163 VNB N_D[3]_c_1685_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_164 VNB N_D[3]_c_1686_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_165 VNB VPWR 1.06677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_166 VNB N_Z_c_2191_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_167 VNB N_Z_c_2192_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_168 VNB N_Z_c_2193_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.19
cc_169 VNB N_Z_c_2194_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.19
cc_170 VNB N_Z_c_2195_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_171 VNB N_Z_c_2196_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_172 VNB N_Z_c_2197_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_173 VNB N_Z_c_2198_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_174 VNB N_Z_c_2199_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_175 VNB N_Z_c_2200_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_176 VNB N_Z_c_2201_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_177 VNB N_Z_c_2202_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_178 VNB N_Z_c_2203_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_179 VNB N_Z_c_2204_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_180 VNB N_Z_c_2205_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_181 VNB N_Z_c_2206_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_182 VNB N_Z_c_2207_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_183 VNB N_Z_c_2208_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_184 VNB N_Z_c_2209_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_185 VNB N_Z_c_2210_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_186 VNB N_Z_c_2211_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_187 VNB N_Z_c_2212_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_188 VNB N_Z_c_2213_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_189 VNB N_Z_c_2214_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_190 VNB N_VGND_c_2906_n 0.0116316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_191 VNB N_VGND_c_2907_n 0.0086067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_192 VNB N_VGND_c_2908_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_193 VNB N_VGND_c_2909_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_194 VNB N_VGND_c_2910_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_195 VNB N_VGND_c_2911_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_196 VNB N_VGND_c_2912_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_197 VNB N_VGND_c_2913_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_198 VNB N_VGND_c_2914_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_199 VNB N_VGND_c_2915_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_200 VNB N_VGND_c_2916_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_201 VNB N_VGND_c_2917_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_202 VNB N_VGND_c_2918_n 0.00916474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_203 VNB N_VGND_c_2919_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_204 VNB N_VGND_c_2920_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_205 VNB N_VGND_c_2921_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_206 VNB N_VGND_c_2922_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_207 VNB N_VGND_c_2923_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_208 VNB N_VGND_c_2924_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_209 VNB N_VGND_c_2925_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_210 VNB N_VGND_c_2926_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_211 VNB N_VGND_c_2927_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_212 VNB N_VGND_c_2928_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_213 VNB N_VGND_c_2929_n 0.0116316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_214 VNB N_VGND_c_2930_n 0.0086067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_215 VNB N_VGND_c_2931_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_216 VNB N_VGND_c_2932_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_217 VNB N_VGND_c_2933_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_218 VNB N_VGND_c_2934_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_219 VNB N_VGND_c_2935_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_220 VNB N_VGND_c_2936_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_221 VNB N_VGND_c_2937_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_222 VNB N_VGND_c_2938_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_223 VNB N_VGND_c_2939_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_224 VNB N_VGND_c_2940_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_225 VNB N_VGND_c_2941_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_226 VNB N_VGND_c_2942_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_227 VNB N_VGND_c_2943_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_228 VNB N_VGND_c_2944_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_229 VNB N_VGND_c_2945_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_230 VNB N_VGND_c_2946_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_231 VNB N_VGND_c_2947_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_232 VNB N_VGND_c_2948_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_233 VNB N_VGND_c_2949_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_234 VNB N_VGND_c_2950_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_235 VNB VGND 1.19676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_236 VNB N_VGND_c_2952_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_237 VNB N_VGND_c_2953_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_238 VNB N_VGND_c_2954_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_239 VNB N_VGND_c_2955_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_240 VNB N_VGND_c_2956_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_241 VNB N_VGND_c_2957_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_242 VNB N_VGND_c_2958_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_243 VNB N_VGND_c_2959_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_244 VNB N_VGND_c_2960_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_245 VNB N_VGND_c_2961_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_246 VNB N_VGND_c_2962_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_247 VNB N_VGND_c_2963_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_248 VNB N_VGND_c_2964_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_249 VNB N_VGND_c_2965_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_250 VNB N_A_119_47#_c_3246_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.025
cc_251 VNB N_A_119_47#_c_3247_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_252 VNB N_A_119_47#_c_3248_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=1.905
+ $Y2=1.985
cc_253 VNB N_A_119_47#_c_3249_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_254 VNB N_A_119_47#_c_3250_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=0.605
+ $Y2=1.105
cc_255 VNB N_A_119_47#_c_3251_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_256 VNB N_A_119_47#_c_3252_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_257 VNB N_A_119_47#_c_3253_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_258 VNB N_A_1693_66#_c_3329_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=1.435
+ $Y2=1.985
cc_259 VNB N_A_1693_66#_c_3330_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_260 VNB N_A_1693_66#_c_3331_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=1.46
+ $Y2=1.025
cc_261 VNB N_A_1693_66#_c_3332_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_262 VNB N_A_1693_66#_c_3333_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=1.905
+ $Y2=1.985
cc_263 VNB N_A_1693_66#_c_3334_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_264 VNB N_A_1693_66#_c_3335_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=0.605
+ $Y2=1.105
cc_265 VNB N_A_1693_66#_c_3336_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_266 VNB N_A_1693_66#_c_3337_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_267 VNB N_A_2695_47#_c_3413_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.46
+ $Y2=1.025
cc_268 VNB N_A_2695_47#_c_3414_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_269 VNB N_A_2695_47#_c_3415_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=1.905
+ $Y2=1.985
cc_270 VNB N_A_2695_47#_c_3416_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_271 VNB N_A_2695_47#_c_3417_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=0.605
+ $Y2=1.105
cc_272 VNB N_A_2695_47#_c_3418_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_273 VNB N_A_2695_47#_c_3419_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_274 VNB N_A_2695_47#_c_3420_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_275 VNB N_A_4269_66#_c_3496_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=1.435
+ $Y2=1.985
cc_276 VNB N_A_4269_66#_c_3497_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_277 VNB N_A_4269_66#_c_3498_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=1.46
+ $Y2=1.025
cc_278 VNB N_A_4269_66#_c_3499_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_279 VNB N_A_4269_66#_c_3500_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=1.905
+ $Y2=1.985
cc_280 VNB N_A_4269_66#_c_3501_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_281 VNB N_A_4269_66#_c_3502_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=0.605
+ $Y2=1.105
cc_282 VNB N_A_4269_66#_c_3503_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_283 VNB N_A_4269_66#_c_3504_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_284 VPB N_D[0]_M1003_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_285 VPB N_D[0]_M1041_g 0.0219201f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_286 VPB N_D[0]_M1055_g 0.0219201f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_287 VPB N_D[0]_M1071_g 0.0300864f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_288 VPB N_D[0]_c_496_n 0.00910964f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_289 VPB N_A_559_265#_c_576_n 0.0263825f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_290 VPB N_A_559_265#_c_577_n 0.0145708f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_291 VPB N_A_559_265#_c_578_n 0.0168203f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_292 VPB N_A_559_265#_c_579_n 0.0213854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_293 VPB N_A_559_265#_c_580_n 0.013221f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_294 VPB N_A_559_265#_c_581_n 0.0213854f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.295
cc_295 VPB N_A_559_265#_c_582_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_296 VPB N_A_559_265#_c_583_n 0.027976f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_297 VPB N_A_559_265#_c_584_n 0.00747525f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.025
cc_298 VPB N_A_559_265#_c_585_n 0.00800249f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_299 VPB N_A_559_265#_c_569_n 0.00733901f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_300 VPB N_A_559_265#_c_570_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_301 VPB N_A_559_265#_c_588_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_302 VPB N_A_559_265#_c_574_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.16
cc_303 VPB N_A_559_265#_c_590_n 0.00195069f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_304 VPB N_A_559_265#_c_575_n 0.0215674f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_305 VPB N_S[0]_c_698_n 0.00781808f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_306 VPB N_S[0]_c_709_n 0.0302591f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_307 VPB N_S[0]_c_702_n 0.0568258f $X=-0.19 $Y=1.305 $X2=1.28 $Y2=1.16
cc_308 VPB S[0] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_309 VPB N_S[1]_c_801_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.295
cc_310 VPB N_S[1]_c_802_n 0.0435876f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_311 VPB N_S[1]_c_806_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_312 VPB N_S[1]_c_826_n 0.0302591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_313 VPB N_S[1]_c_822_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_314 VPB N_A_1430_325#_c_926_n 0.027976f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_315 VPB N_A_1430_325#_c_927_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_316 VPB N_A_1430_325#_c_919_n 0.0215674f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_317 VPB N_A_1430_325#_c_929_n 0.0213854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_318 VPB N_A_1430_325#_c_930_n 0.013221f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_319 VPB N_A_1430_325#_c_931_n 0.0213854f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.295
cc_320 VPB N_A_1430_325#_c_932_n 0.0312612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_321 VPB N_A_1430_325#_c_933_n 0.0263825f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_322 VPB N_A_1430_325#_c_934_n 0.00800249f $X=-0.19 $Y=1.305 $X2=1.88
+ $Y2=1.025
cc_323 VPB N_A_1430_325#_c_935_n 0.00747525f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_324 VPB N_A_1430_325#_c_936_n 0.00751381f $X=-0.19 $Y=1.305 $X2=1.905
+ $Y2=1.295
cc_325 VPB N_A_1430_325#_c_922_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_326 VPB N_A_1430_325#_c_938_n 0.00195069f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.16
cc_327 VPB N_A_1430_325#_c_924_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_328 VPB N_A_1430_325#_c_925_n 0.0150864f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_329 VPB N_D[1]_M1001_g 0.0300864f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_330 VPB N_D[1]_M1006_g 0.0219201f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_331 VPB N_D[1]_M1038_g 0.0219201f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_332 VPB N_D[1]_M1065_g 0.0296461f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_333 VPB N_D[1]_c_1045_n 0.0083121f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_334 VPB N_D[2]_M1005_g 0.0296461f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_335 VPB N_D[2]_M1019_g 0.0219201f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_336 VPB N_D[2]_M1047_g 0.0219201f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_337 VPB N_D[2]_M1074_g 0.0300864f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_338 VPB N_D[2]_c_1131_n 0.0083121f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_339 VPB N_A_3135_265#_c_1216_n 0.0263825f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_340 VPB N_A_3135_265#_c_1217_n 0.0145708f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_341 VPB N_A_3135_265#_c_1218_n 0.0166904f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_342 VPB N_A_3135_265#_c_1219_n 0.0213854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_343 VPB N_A_3135_265#_c_1220_n 0.013221f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_344 VPB N_A_3135_265#_c_1221_n 0.0213854f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.295
cc_345 VPB N_A_3135_265#_c_1222_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_346 VPB N_A_3135_265#_c_1223_n 0.027976f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_347 VPB N_A_3135_265#_c_1224_n 0.00747525f $X=-0.19 $Y=1.305 $X2=1.88
+ $Y2=1.025
cc_348 VPB N_A_3135_265#_c_1225_n 0.00800249f $X=-0.19 $Y=1.305 $X2=1.88
+ $Y2=0.56
cc_349 VPB N_A_3135_265#_c_1209_n 0.00733901f $X=-0.19 $Y=1.305 $X2=1.88
+ $Y2=0.56
cc_350 VPB N_A_3135_265#_c_1210_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_351 VPB N_A_3135_265#_c_1228_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.16
cc_352 VPB N_A_3135_265#_c_1214_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=1.46
+ $Y2=1.16
cc_353 VPB N_A_3135_265#_c_1230_n 0.00195069f $X=-0.19 $Y=1.305 $X2=1.62
+ $Y2=1.16
cc_354 VPB N_A_3135_265#_c_1215_n 0.0215674f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_355 VPB N_S[2]_c_1340_n 0.00781808f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_356 VPB N_S[2]_c_1351_n 0.0302591f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_357 VPB N_S[2]_c_1344_n 0.0568258f $X=-0.19 $Y=1.305 $X2=1.28 $Y2=1.16
cc_358 VPB S[2] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_359 VPB N_S[3]_c_1443_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.295
cc_360 VPB N_S[3]_c_1444_n 0.0435876f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_361 VPB N_S[3]_c_1448_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_362 VPB N_S[3]_c_1468_n 0.0302591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_363 VPB N_S[3]_c_1464_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_364 VPB N_A_4006_325#_c_1568_n 0.027976f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_365 VPB N_A_4006_325#_c_1569_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_366 VPB N_A_4006_325#_c_1561_n 0.0215674f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_367 VPB N_A_4006_325#_c_1571_n 0.0213854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_368 VPB N_A_4006_325#_c_1572_n 0.013221f $X=-0.19 $Y=1.305 $X2=0.965
+ $Y2=1.985
cc_369 VPB N_A_4006_325#_c_1573_n 0.0213854f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.295
cc_370 VPB N_A_4006_325#_c_1574_n 0.0313911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_371 VPB N_A_4006_325#_c_1575_n 0.0263825f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_372 VPB N_A_4006_325#_c_1576_n 0.00800249f $X=-0.19 $Y=1.305 $X2=1.88
+ $Y2=1.025
cc_373 VPB N_A_4006_325#_c_1577_n 0.00747525f $X=-0.19 $Y=1.305 $X2=1.88
+ $Y2=0.56
cc_374 VPB N_A_4006_325#_c_1578_n 0.00751381f $X=-0.19 $Y=1.305 $X2=1.905
+ $Y2=1.295
cc_375 VPB N_A_4006_325#_c_1564_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.16
cc_376 VPB N_A_4006_325#_c_1580_n 0.00195069f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.16
cc_377 VPB N_A_4006_325#_c_1566_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=1.62
+ $Y2=1.16
cc_378 VPB N_A_4006_325#_c_1567_n 0.0150864f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_379 VPB N_D[3]_M1010_g 0.0300864f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_380 VPB N_D[3]_M1027_g 0.0219201f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_381 VPB N_D[3]_M1035_g 0.0219201f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_382 VPB N_D[3]_M1070_g 0.0296461f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_383 VPB N_D[3]_c_1685_n 0.00910964f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_384 VPB N_VPWR_c_1757_n 0.0113525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_385 VPB N_VPWR_c_1758_n 0.0413001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_386 VPB N_VPWR_c_1759_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_387 VPB N_VPWR_c_1760_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_388 VPB N_VPWR_c_1761_n 0.0103001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_389 VPB N_VPWR_c_1762_n 0.0169817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_390 VPB N_VPWR_c_1763_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_391 VPB N_VPWR_c_1764_n 0.013938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_392 VPB N_VPWR_c_1765_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_393 VPB N_VPWR_c_1766_n 0.0169817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_394 VPB N_VPWR_c_1767_n 0.00986069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_395 VPB N_VPWR_c_1768_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_396 VPB N_VPWR_c_1769_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_397 VPB N_VPWR_c_1770_n 0.00789186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_398 VPB N_VPWR_c_1771_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_399 VPB N_VPWR_c_1772_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_400 VPB N_VPWR_c_1773_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_401 VPB N_VPWR_c_1774_n 0.00986069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_402 VPB N_VPWR_c_1775_n 0.0169817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_403 VPB N_VPWR_c_1776_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_404 VPB N_VPWR_c_1777_n 0.013938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_405 VPB N_VPWR_c_1778_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_406 VPB N_VPWR_c_1779_n 0.0169817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_407 VPB N_VPWR_c_1780_n 0.0103001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_408 VPB N_VPWR_c_1781_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_409 VPB N_VPWR_c_1782_n 0.0113525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_410 VPB N_VPWR_c_1783_n 0.0413001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_411 VPB N_VPWR_c_1784_n 0.0637101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_412 VPB N_VPWR_c_1785_n 0.00526366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_413 VPB N_VPWR_c_1786_n 0.0187412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_414 VPB N_VPWR_c_1787_n 0.00574121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_415 VPB N_VPWR_c_1788_n 0.0187412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_416 VPB N_VPWR_c_1789_n 0.00526366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_417 VPB N_VPWR_c_1790_n 0.0637101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_418 VPB N_VPWR_c_1791_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_419 VPB N_VPWR_c_1792_n 0.0637101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_420 VPB N_VPWR_c_1793_n 0.00526366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_421 VPB N_VPWR_c_1794_n 0.0187412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_422 VPB N_VPWR_c_1795_n 0.00574121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_423 VPB N_VPWR_c_1796_n 0.0187412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_424 VPB N_VPWR_c_1797_n 0.00526366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_425 VPB N_VPWR_c_1798_n 0.0637101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_426 VPB N_VPWR_c_1799_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_427 VPB VPWR 0.140555f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_428 VPB N_VPWR_c_1801_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_429 VPB N_VPWR_c_1802_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_430 VPB N_VPWR_c_1803_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_431 VPB N_VPWR_c_1804_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_432 VPB N_VPWR_c_1805_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_433 VPB N_VPWR_c_1806_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_434 VPB N_VPWR_c_1807_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_435 VPB N_VPWR_c_1808_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_436 VPB N_VPWR_c_1809_n 0.00574121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_437 VPB N_VPWR_c_1810_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_438 VPB N_VPWR_c_1811_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_439 VPB N_VPWR_c_1812_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_440 VPB N_VPWR_c_1813_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_441 VPB N_VPWR_c_1814_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_442 VPB N_VPWR_c_1815_n 0.00574121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_443 VPB N_VPWR_c_1816_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_444 VPB N_A_117_297#_c_2102_n 0.0199901f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_445 VPB N_A_117_297#_c_2103_n 0.00635149f $X=-0.19 $Y=1.305 $X2=1.905
+ $Y2=1.985
cc_446 VPB N_A_117_297#_c_2104_n 0.00219354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_447 VPB N_A_117_297#_c_2105_n 0.00409031f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=1.105
cc_448 VPB N_A_117_297#_c_2106_n 0.00229202f $X=-0.19 $Y=1.305 $X2=1.055
+ $Y2=1.16
cc_449 VPB N_A_117_297#_c_2107_n 0.00637482f $X=-0.19 $Y=1.305 $X2=1.28 $Y2=1.16
cc_450 VPB N_A_117_297#_c_2108_n 0.00712701f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_451 VPB N_A_117_297#_c_2109_n 0.00196597f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.16
cc_452 VPB N_Z_c_2204_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_453 VPB N_Z_c_2207_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_454 VPB N_Z_c_2210_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_455 VPB N_Z_c_2213_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_456 VPB N_Z_c_2219_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_457 VPB N_Z_c_2220_n 0.0210274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_458 VPB N_Z_c_2221_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_459 VPB N_A_1643_311#_c_2607_n 0.00712701f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.985
cc_460 VPB N_A_1643_311#_c_2608_n 0.00219354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_461 VPB N_A_1643_311#_c_2609_n 0.00418127f $X=-0.19 $Y=1.305 $X2=1.46
+ $Y2=1.025
cc_462 VPB N_A_1643_311#_c_2610_n 0.00229202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_463 VPB N_A_1643_311#_c_2611_n 0.00628386f $X=-0.19 $Y=1.305 $X2=1.88
+ $Y2=0.56
cc_464 VPB N_A_1643_311#_c_2612_n 0.00591976f $X=-0.19 $Y=1.305 $X2=1.905
+ $Y2=1.985
cc_465 VPB N_A_1643_311#_c_2613_n 0.0075016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_466 VPB N_A_1643_311#_c_2614_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=1.105
cc_467 VPB N_A_1643_311#_c_2615_n 0.00196597f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.16
cc_468 VPB N_A_2693_297#_c_2712_n 0.0147622f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_469 VPB N_A_2693_297#_c_2713_n 0.00591976f $X=-0.19 $Y=1.305 $X2=1.905
+ $Y2=1.985
cc_470 VPB N_A_2693_297#_c_2714_n 0.00219354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_471 VPB N_A_2693_297#_c_2715_n 0.00409031f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=1.105
cc_472 VPB N_A_2693_297#_c_2716_n 0.00229202f $X=-0.19 $Y=1.305 $X2=1.055
+ $Y2=1.16
cc_473 VPB N_A_2693_297#_c_2717_n 0.00637482f $X=-0.19 $Y=1.305 $X2=1.28
+ $Y2=1.16
cc_474 VPB N_A_2693_297#_c_2718_n 0.00712701f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=1.16
cc_475 VPB N_A_2693_297#_c_2719_n 0.00196597f $X=-0.19 $Y=1.305 $X2=1.46
+ $Y2=1.16
cc_476 VPB N_A_4219_311#_c_2814_n 0.00712701f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.985
cc_477 VPB N_A_4219_311#_c_2815_n 0.00219354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_478 VPB N_A_4219_311#_c_2816_n 0.00418127f $X=-0.19 $Y=1.305 $X2=1.46
+ $Y2=1.025
cc_479 VPB N_A_4219_311#_c_2817_n 0.00229202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_480 VPB N_A_4219_311#_c_2818_n 0.00628386f $X=-0.19 $Y=1.305 $X2=1.88
+ $Y2=0.56
cc_481 VPB N_A_4219_311#_c_2819_n 0.00635149f $X=-0.19 $Y=1.305 $X2=1.905
+ $Y2=1.985
cc_482 VPB N_A_4219_311#_c_2820_n 0.0127295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_483 VPB N_A_4219_311#_c_2821_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=1.105
cc_484 VPB N_A_4219_311#_c_2822_n 0.00196597f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.16
cc_485 N_D[0]_M1003_g N_VPWR_c_1758_n 0.00354866f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_486 N_D[0]_M1041_g N_VPWR_c_1759_n 0.00173895f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_487 N_D[0]_M1055_g N_VPWR_c_1759_n 0.00173895f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_488 N_D[0]_M1055_g N_VPWR_c_1760_n 0.00673617f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_489 N_D[0]_M1071_g N_VPWR_c_1760_n 0.00673617f $X=1.905 $Y=1.985 $X2=0 $Y2=0
cc_490 N_D[0]_M1071_g N_VPWR_c_1761_n 0.00354866f $X=1.905 $Y=1.985 $X2=0 $Y2=0
cc_491 N_D[0]_M1003_g VPWR 0.0126298f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_492 N_D[0]_M1041_g VPWR 0.0117184f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_493 N_D[0]_M1055_g VPWR 0.0117184f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_494 N_D[0]_M1071_g VPWR 0.0130007f $X=1.905 $Y=1.985 $X2=0 $Y2=0
cc_495 N_D[0]_M1003_g N_VPWR_c_1801_n 0.00673617f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_496 N_D[0]_M1041_g N_VPWR_c_1801_n 0.00673617f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_497 N_D[0]_M1003_g N_A_117_297#_c_2110_n 0.00215964f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_498 N_D[0]_M1041_g N_A_117_297#_c_2110_n 5.79575e-19 $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_D[0]_c_495_n N_A_117_297#_c_2110_n 8.03631e-19 $X=1.055 $Y=1.16 $X2=0
+ $Y2=0
cc_500 N_D[0]_c_496_n N_A_117_297#_c_2110_n 0.022724f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_501 N_D[0]_M1003_g N_A_117_297#_c_2114_n 0.00897418f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_502 N_D[0]_M1041_g N_A_117_297#_c_2114_n 0.0100233f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_503 N_D[0]_M1055_g N_A_117_297#_c_2114_n 5.91934e-19 $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_504 N_D[0]_M1041_g N_A_117_297#_c_2117_n 0.0137916f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_505 N_D[0]_M1055_g N_A_117_297#_c_2117_n 0.0137916f $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_506 N_D[0]_c_494_n N_A_117_297#_c_2117_n 7.15862e-19 $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_507 N_D[0]_c_496_n N_A_117_297#_c_2117_n 0.0405252f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_508 N_D[0]_M1041_g N_A_117_297#_c_2121_n 5.91934e-19 $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_509 N_D[0]_M1055_g N_A_117_297#_c_2121_n 0.0100233f $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_510 N_D[0]_M1071_g N_A_117_297#_c_2121_n 0.010906f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_511 N_D[0]_M1071_g N_A_117_297#_c_2102_n 0.017872f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_512 N_D[0]_M1071_g N_A_117_297#_c_2103_n 0.00330737f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_513 N_D[0]_M1055_g N_A_117_297#_c_2126_n 5.79575e-19 $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_514 N_D[0]_M1071_g N_A_117_297#_c_2126_n 8.61029e-19 $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_515 N_D[0]_c_496_n N_A_117_297#_c_2126_n 0.0199757f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_516 N_D[0]_c_497_n N_A_117_297#_c_2126_n 8.03631e-19 $X=1.905 $Y=1.16 $X2=0
+ $Y2=0
cc_517 N_D[0]_M1024_g N_VGND_c_2907_n 0.00345859f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_518 N_D[0]_M1024_g N_VGND_c_2908_n 2.64031e-19 $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_519 N_D[0]_M1057_g N_VGND_c_2908_n 0.00166854f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_520 N_D[0]_M1073_g N_VGND_c_2908_n 0.0019152f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_521 N_D[0]_M1073_g N_VGND_c_2909_n 0.00430643f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_522 N_D[0]_M1078_g N_VGND_c_2909_n 0.00422241f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_523 N_D[0]_M1073_g N_VGND_c_2910_n 2.6376e-19 $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_524 N_D[0]_M1078_g N_VGND_c_2910_n 0.00321269f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_525 N_D[0]_M1024_g VGND 0.0107845f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_526 N_D[0]_M1057_g VGND 0.00593887f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_527 N_D[0]_M1073_g VGND 0.00624811f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_528 N_D[0]_M1078_g VGND 0.00702263f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_529 N_D[0]_M1024_g N_VGND_c_2952_n 0.00551064f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_530 N_D[0]_M1057_g N_VGND_c_2952_n 0.00422241f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_531 N_D[0]_M1024_g N_A_119_47#_c_3254_n 0.00529286f $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_532 N_D[0]_M1057_g N_A_119_47#_c_3254_n 0.00661134f $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_533 N_D[0]_M1073_g N_A_119_47#_c_3254_n 5.22365e-19 $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_534 N_D[0]_M1057_g N_A_119_47#_c_3257_n 0.00899636f $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_535 N_D[0]_M1073_g N_A_119_47#_c_3257_n 0.00900364f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_536 N_D[0]_c_494_n N_A_119_47#_c_3257_n 0.00463549f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_537 N_D[0]_c_496_n N_A_119_47#_c_3257_n 0.0394855f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_538 N_D[0]_M1024_g N_A_119_47#_c_3246_n 0.00228093f $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_539 N_D[0]_M1057_g N_A_119_47#_c_3246_n 8.68782e-19 $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_540 N_D[0]_c_495_n N_A_119_47#_c_3246_n 0.00208088f $X=1.055 $Y=1.16 $X2=0
+ $Y2=0
cc_541 N_D[0]_c_496_n N_A_119_47#_c_3246_n 0.021403f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_542 N_D[0]_M1057_g N_A_119_47#_c_3265_n 5.22365e-19 $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_543 N_D[0]_M1073_g N_A_119_47#_c_3265_n 0.00661764f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_544 N_D[0]_M1078_g N_A_119_47#_c_3265_n 0.00699463f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_545 N_D[0]_M1078_g N_A_119_47#_c_3247_n 0.0121912f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_546 N_D[0]_M1078_g N_A_119_47#_c_3248_n 0.00261078f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_547 N_D[0]_M1073_g N_A_119_47#_c_3253_n 8.68782e-19 $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_548 N_D[0]_M1078_g N_A_119_47#_c_3253_n 0.00128201f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_549 N_D[0]_c_496_n N_A_119_47#_c_3253_n 0.018367f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_550 N_D[0]_c_497_n N_A_119_47#_c_3253_n 0.00208088f $X=1.905 $Y=1.16 $X2=0
+ $Y2=0
cc_551 N_A_559_265#_c_578_n N_S[0]_c_686_n 0.00507426f $X=2.985 $Y=1.4 $X2=-0.19
+ $Y2=-0.24
cc_552 N_A_559_265#_c_577_n N_S[0]_c_689_n 0.00509391f $X=3.275 $Y=1.4 $X2=0
+ $Y2=0
cc_553 N_A_559_265#_c_580_n N_S[0]_c_691_n 0.00509204f $X=3.745 $Y=1.4 $X2=0
+ $Y2=0
cc_554 N_A_559_265#_c_582_n N_S[0]_c_693_n 0.00507688f $X=4.215 $Y=1.4 $X2=0
+ $Y2=0
cc_555 N_A_559_265#_c_571_n N_S[0]_c_695_n 6.53442e-19 $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_556 N_A_559_265#_c_569_n N_S[0]_c_697_n 0.0103812f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_557 N_A_559_265#_c_570_n N_S[0]_c_697_n 0.0179529f $X=4.875 $Y=1.23 $X2=0
+ $Y2=0
cc_558 N_A_559_265#_c_569_n N_S[0]_c_698_n 0.0206368f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_559 N_A_559_265#_c_570_n N_S[0]_c_698_n 0.0175393f $X=4.875 $Y=1.23 $X2=0
+ $Y2=0
cc_560 N_A_559_265#_c_572_n N_S[0]_c_698_n 0.0085951f $X=5.505 $Y=1.065 $X2=0
+ $Y2=0
cc_561 N_A_559_265#_c_574_n N_S[0]_c_698_n 0.00322131f $X=5.505 $Y=1.23 $X2=0
+ $Y2=0
cc_562 N_A_559_265#_c_590_n N_S[0]_c_698_n 0.00255921f $X=5.585 $Y=1.605 $X2=0
+ $Y2=0
cc_563 N_A_559_265#_c_575_n N_S[0]_c_698_n 0.00262132f $X=4.625 $Y=1.23 $X2=0
+ $Y2=0
cc_564 N_A_559_265#_c_588_n N_S[0]_c_709_n 0.0118819f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_565 N_A_559_265#_c_590_n N_S[0]_c_709_n 0.00762115f $X=5.585 $Y=1.605 $X2=0
+ $Y2=0
cc_566 N_A_559_265#_c_571_n N_S[0]_c_699_n 0.00603996f $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_567 N_A_559_265#_c_573_n N_S[0]_c_699_n 9.67113e-19 $X=5.545 $Y=0.825 $X2=0
+ $Y2=0
cc_568 N_A_559_265#_c_572_n N_S[0]_c_700_n 0.00429801f $X=5.505 $Y=1.065 $X2=0
+ $Y2=0
cc_569 N_A_559_265#_c_573_n N_S[0]_c_700_n 0.0111895f $X=5.545 $Y=0.825 $X2=0
+ $Y2=0
cc_570 N_A_559_265#_c_571_n N_S[0]_c_701_n 0.00207203f $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_571 N_A_559_265#_c_572_n N_S[0]_c_702_n 0.00289358f $X=5.505 $Y=1.065 $X2=0
+ $Y2=0
cc_572 N_A_559_265#_c_588_n N_S[0]_c_702_n 0.0128955f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_573 N_A_559_265#_c_574_n N_S[0]_c_702_n 0.00416423f $X=5.505 $Y=1.23 $X2=0
+ $Y2=0
cc_574 N_A_559_265#_c_590_n N_S[0]_c_702_n 0.00454075f $X=5.585 $Y=1.605 $X2=0
+ $Y2=0
cc_575 N_A_559_265#_c_572_n N_S[0]_c_706_n 0.00268644f $X=5.505 $Y=1.065 $X2=0
+ $Y2=0
cc_576 N_A_559_265#_c_573_n N_S[0]_c_706_n 0.00426435f $X=5.545 $Y=0.825 $X2=0
+ $Y2=0
cc_577 N_A_559_265#_c_572_n S[0] 0.00541767f $X=5.505 $Y=1.065 $X2=0 $Y2=0
cc_578 N_A_559_265#_c_574_n S[0] 0.0228692f $X=5.505 $Y=1.23 $X2=0 $Y2=0
cc_579 N_A_559_265#_c_576_n N_VPWR_c_1761_n 0.00287722f $X=2.895 $Y=1.475 $X2=0
+ $Y2=0
cc_580 N_A_559_265#_c_583_n N_VPWR_c_1762_n 0.00279288f $X=4.305 $Y=1.475 $X2=0
+ $Y2=0
cc_581 N_A_559_265#_c_569_n N_VPWR_c_1762_n 0.0193185f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_582 N_A_559_265#_c_570_n N_VPWR_c_1762_n 6.4101e-19 $X=4.875 $Y=1.23 $X2=0
+ $Y2=0
cc_583 N_A_559_265#_c_588_n N_VPWR_c_1762_n 0.0316788f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_584 N_A_559_265#_c_588_n N_VPWR_c_1763_n 0.0356181f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_585 N_A_559_265#_c_576_n N_VPWR_c_1784_n 0.00429453f $X=2.895 $Y=1.475 $X2=0
+ $Y2=0
cc_586 N_A_559_265#_c_579_n N_VPWR_c_1784_n 0.00429453f $X=3.365 $Y=1.475 $X2=0
+ $Y2=0
cc_587 N_A_559_265#_c_581_n N_VPWR_c_1784_n 0.00429453f $X=3.835 $Y=1.475 $X2=0
+ $Y2=0
cc_588 N_A_559_265#_c_583_n N_VPWR_c_1784_n 0.00429453f $X=4.305 $Y=1.475 $X2=0
+ $Y2=0
cc_589 N_A_559_265#_c_588_n N_VPWR_c_1786_n 0.0233824f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_590 N_A_559_265#_c_576_n VPWR 0.00743756f $X=2.895 $Y=1.475 $X2=0 $Y2=0
cc_591 N_A_559_265#_c_579_n VPWR 0.0060424f $X=3.365 $Y=1.475 $X2=0 $Y2=0
cc_592 N_A_559_265#_c_581_n VPWR 0.0060424f $X=3.835 $Y=1.475 $X2=0 $Y2=0
cc_593 N_A_559_265#_c_583_n VPWR 0.00737407f $X=4.305 $Y=1.475 $X2=0 $Y2=0
cc_594 N_A_559_265#_c_588_n VPWR 0.00593513f $X=5.585 $Y=1.77 $X2=0 $Y2=0
cc_595 N_A_559_265#_c_576_n N_A_117_297#_c_2102_n 0.00151141f $X=2.895 $Y=1.475
+ $X2=0 $Y2=0
cc_596 N_A_559_265#_c_576_n N_A_117_297#_c_2104_n 0.0155783f $X=2.895 $Y=1.475
+ $X2=0 $Y2=0
cc_597 N_A_559_265#_c_579_n N_A_117_297#_c_2104_n 0.010844f $X=3.365 $Y=1.475
+ $X2=0 $Y2=0
cc_598 N_A_559_265#_c_579_n N_A_117_297#_c_2106_n 0.00102951f $X=3.365 $Y=1.475
+ $X2=0 $Y2=0
cc_599 N_A_559_265#_c_580_n N_A_117_297#_c_2106_n 0.00251792f $X=3.745 $Y=1.4
+ $X2=0 $Y2=0
cc_600 N_A_559_265#_c_581_n N_A_117_297#_c_2106_n 0.00102951f $X=3.835 $Y=1.475
+ $X2=0 $Y2=0
cc_601 N_A_559_265#_c_581_n N_A_117_297#_c_2107_n 0.010844f $X=3.835 $Y=1.475
+ $X2=0 $Y2=0
cc_602 N_A_559_265#_c_583_n N_A_117_297#_c_2107_n 0.0115457f $X=4.305 $Y=1.475
+ $X2=0 $Y2=0
cc_603 N_A_559_265#_c_583_n N_A_117_297#_c_2108_n 0.00246857f $X=4.305 $Y=1.475
+ $X2=0 $Y2=0
cc_604 N_A_559_265#_c_569_n N_A_117_297#_c_2108_n 0.0218124f $X=5.42 $Y=1.23
+ $X2=0 $Y2=0
cc_605 N_A_559_265#_c_570_n N_A_117_297#_c_2108_n 5.74251e-19 $X=4.875 $Y=1.23
+ $X2=0 $Y2=0
cc_606 N_A_559_265#_c_575_n N_A_117_297#_c_2108_n 0.00561627f $X=4.625 $Y=1.23
+ $X2=0 $Y2=0
cc_607 N_A_559_265#_c_580_n N_Z_c_2192_n 0.00762343f $X=3.745 $Y=1.4 $X2=0 $Y2=0
cc_608 N_A_559_265#_c_584_n N_Z_c_2192_n 0.00704092f $X=3.365 $Y=1.4 $X2=0 $Y2=0
cc_609 N_A_559_265#_c_578_n N_Z_c_2203_n 0.00248496f $X=2.985 $Y=1.4 $X2=0 $Y2=0
cc_610 N_A_559_265#_c_577_n N_Z_c_2204_n 0.00678861f $X=3.275 $Y=1.4 $X2=0 $Y2=0
cc_611 N_A_559_265#_c_578_n N_Z_c_2204_n 0.00239476f $X=2.985 $Y=1.4 $X2=0 $Y2=0
cc_612 N_A_559_265#_c_584_n N_Z_c_2204_n 2.98555e-19 $X=3.365 $Y=1.4 $X2=0 $Y2=0
cc_613 N_A_559_265#_c_580_n N_Z_c_2205_n 0.00145542f $X=3.745 $Y=1.4 $X2=0 $Y2=0
cc_614 N_A_559_265#_c_582_n N_Z_c_2205_n 0.00597584f $X=4.215 $Y=1.4 $X2=0 $Y2=0
cc_615 N_A_559_265#_c_585_n N_Z_c_2205_n 0.00909323f $X=3.835 $Y=1.4 $X2=0 $Y2=0
cc_616 N_A_559_265#_c_569_n N_Z_c_2205_n 0.0266078f $X=5.42 $Y=1.23 $X2=0 $Y2=0
cc_617 N_A_559_265#_c_575_n N_Z_c_2205_n 0.00747617f $X=4.625 $Y=1.23 $X2=0
+ $Y2=0
cc_618 N_A_559_265#_c_583_n N_Z_c_2219_n 0.0080184f $X=4.305 $Y=1.475 $X2=0
+ $Y2=0
cc_619 N_A_559_265#_c_569_n N_Z_c_2219_n 0.0186685f $X=5.42 $Y=1.23 $X2=0 $Y2=0
cc_620 N_A_559_265#_c_588_n N_Z_c_2219_n 0.0329704f $X=5.585 $Y=1.77 $X2=0 $Y2=0
cc_621 N_A_559_265#_c_575_n N_Z_c_2219_n 2.19754e-19 $X=4.625 $Y=1.23 $X2=0
+ $Y2=0
cc_622 N_A_559_265#_c_579_n Z 0.00378723f $X=3.365 $Y=1.475 $X2=0 $Y2=0
cc_623 N_A_559_265#_c_581_n Z 0.00378512f $X=3.835 $Y=1.475 $X2=0 $Y2=0
cc_624 N_A_559_265#_c_576_n N_Z_c_2239_n 0.00899738f $X=2.895 $Y=1.475 $X2=0
+ $Y2=0
cc_625 N_A_559_265#_c_577_n N_Z_c_2239_n 0.00554725f $X=3.275 $Y=1.4 $X2=0 $Y2=0
cc_626 N_A_559_265#_c_578_n N_Z_c_2239_n 0.00474497f $X=2.985 $Y=1.4 $X2=0 $Y2=0
cc_627 N_A_559_265#_c_579_n N_Z_c_2239_n 0.00814309f $X=3.365 $Y=1.475 $X2=0
+ $Y2=0
cc_628 N_A_559_265#_c_581_n N_Z_c_2239_n 3.67612e-19 $X=3.835 $Y=1.475 $X2=0
+ $Y2=0
cc_629 N_A_559_265#_c_584_n N_Z_c_2239_n 0.00313387f $X=3.365 $Y=1.4 $X2=0 $Y2=0
cc_630 N_A_559_265#_c_579_n N_Z_c_2245_n 3.67612e-19 $X=3.365 $Y=1.475 $X2=0
+ $Y2=0
cc_631 N_A_559_265#_c_581_n N_Z_c_2245_n 0.00814309f $X=3.835 $Y=1.475 $X2=0
+ $Y2=0
cc_632 N_A_559_265#_c_582_n N_Z_c_2245_n 0.00554725f $X=4.215 $Y=1.4 $X2=0 $Y2=0
cc_633 N_A_559_265#_c_583_n N_Z_c_2245_n 0.0107691f $X=4.305 $Y=1.475 $X2=0
+ $Y2=0
cc_634 N_A_559_265#_c_585_n N_Z_c_2245_n 0.00313387f $X=3.835 $Y=1.4 $X2=0 $Y2=0
cc_635 N_A_559_265#_c_569_n N_Z_c_2245_n 0.00227722f $X=5.42 $Y=1.23 $X2=0 $Y2=0
cc_636 N_A_559_265#_c_575_n N_Z_c_2245_n 0.00415799f $X=4.625 $Y=1.23 $X2=0
+ $Y2=0
cc_637 N_A_559_265#_c_569_n N_VGND_c_2911_n 0.0123065f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_638 N_A_559_265#_c_570_n N_VGND_c_2911_n 2.04129e-19 $X=4.875 $Y=1.23 $X2=0
+ $Y2=0
cc_639 N_A_559_265#_c_571_n N_VGND_c_2933_n 0.0129994f $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_640 N_A_559_265#_M1046_d VGND 0.00394793f $X=5.45 $Y=0.235 $X2=0 $Y2=0
cc_641 N_A_559_265#_c_571_n VGND 0.00927134f $X=5.585 $Y=0.445 $X2=0 $Y2=0
cc_642 N_A_559_265#_c_584_n N_A_119_47#_c_3274_n 7.0477e-19 $X=3.365 $Y=1.4
+ $X2=0 $Y2=0
cc_643 N_A_559_265#_c_569_n N_A_119_47#_c_3252_n 0.0028695f $X=5.42 $Y=1.23
+ $X2=0 $Y2=0
cc_644 N_A_559_265#_c_575_n N_A_119_47#_c_3252_n 0.00589316f $X=4.625 $Y=1.23
+ $X2=0 $Y2=0
cc_645 N_S[0]_c_702_n N_S[1]_c_801_n 0.0215827f $X=5.82 $Y=1.55 $X2=-0.19
+ $Y2=-0.24
cc_646 S[0] N_S[1]_c_801_n 0.00113563f $X=6.125 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_647 N_S[0]_c_702_n N_S[1]_c_822_n 0.00113563f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_648 S[0] N_S[1]_c_822_n 0.0301108f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_649 N_S[0]_c_709_n N_VPWR_c_1762_n 0.00950399f $X=5.35 $Y=1.55 $X2=0 $Y2=0
cc_650 N_S[0]_c_702_n N_VPWR_c_1763_n 0.016386f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_651 S[0] N_VPWR_c_1763_n 0.0157609f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_652 N_S[0]_c_709_n N_VPWR_c_1786_n 0.00673617f $X=5.35 $Y=1.55 $X2=0 $Y2=0
cc_653 N_S[0]_c_702_n N_VPWR_c_1786_n 0.00673617f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_654 N_S[0]_c_709_n VPWR 0.00852996f $X=5.35 $Y=1.55 $X2=0 $Y2=0
cc_655 N_S[0]_c_702_n VPWR 0.00846723f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_656 N_S[0]_c_686_n N_A_117_297#_c_2102_n 0.00168571f $X=2.82 $Y=0.255 $X2=0
+ $Y2=0
cc_657 N_S[0]_c_709_n N_A_117_297#_c_2108_n 0.00209354f $X=5.35 $Y=1.55 $X2=0
+ $Y2=0
cc_658 N_S[0]_c_686_n N_Z_c_2191_n 0.002324f $X=2.82 $Y=0.255 $X2=0 $Y2=0
cc_659 N_S[0]_c_689_n N_Z_c_2191_n 0.00283489f $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_660 N_S[0]_c_689_n N_Z_c_2192_n 3.10191e-19 $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_661 N_S[0]_c_691_n N_Z_c_2192_n 0.00190704f $X=3.66 $Y=0.255 $X2=0 $Y2=0
cc_662 N_S[0]_c_689_n N_Z_c_2193_n 6.35774e-19 $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_663 N_S[0]_c_691_n N_Z_c_2193_n 0.0077801f $X=3.66 $Y=0.255 $X2=0 $Y2=0
cc_664 N_S[0]_c_693_n N_Z_c_2193_n 0.0134253f $X=4.08 $Y=0.255 $X2=0 $Y2=0
cc_665 N_S[0]_c_686_n N_Z_c_2203_n 0.00443615f $X=2.82 $Y=0.255 $X2=0 $Y2=0
cc_666 N_S[0]_c_689_n N_Z_c_2203_n 0.00462308f $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_667 N_S[0]_c_691_n N_Z_c_2203_n 6.35664e-19 $X=3.66 $Y=0.255 $X2=0 $Y2=0
cc_668 N_S[0]_c_689_n N_Z_c_2204_n 0.00180363f $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_669 N_S[0]_c_693_n N_Z_c_2205_n 0.00216436f $X=4.08 $Y=0.255 $X2=0 $Y2=0
cc_670 N_S[0]_c_709_n N_Z_c_2219_n 0.00478771f $X=5.35 $Y=1.55 $X2=0 $Y2=0
cc_671 N_S[0]_c_702_n N_Z_c_2219_n 0.00760321f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_672 S[0] N_Z_c_2219_n 0.010609f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_673 N_S[0]_c_686_n N_VGND_c_2910_n 5.5039e-19 $X=2.82 $Y=0.255 $X2=0 $Y2=0
cc_674 N_S[0]_c_688_n N_VGND_c_2910_n 0.0028166f $X=2.895 $Y=0.18 $X2=0 $Y2=0
cc_675 N_S[0]_c_694_n N_VGND_c_2911_n 0.00862298f $X=4.765 $Y=0.18 $X2=0 $Y2=0
cc_676 N_S[0]_c_696_n N_VGND_c_2911_n 0.00525833f $X=5.25 $Y=0.81 $X2=0 $Y2=0
cc_677 N_S[0]_c_699_n N_VGND_c_2911_n 0.00173127f $X=5.375 $Y=0.735 $X2=0 $Y2=0
cc_678 N_S[0]_c_701_n N_VGND_c_2912_n 0.00374526f $X=5.795 $Y=0.735 $X2=0 $Y2=0
cc_679 N_S[0]_c_702_n N_VGND_c_2912_n 0.00578076f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_680 S[0] N_VGND_c_2912_n 0.0116413f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_681 N_S[0]_c_688_n N_VGND_c_2931_n 0.0559651f $X=2.895 $Y=0.18 $X2=0 $Y2=0
cc_682 N_S[0]_c_699_n N_VGND_c_2933_n 0.00542362f $X=5.375 $Y=0.735 $X2=0 $Y2=0
cc_683 N_S[0]_c_700_n N_VGND_c_2933_n 2.16067e-19 $X=5.72 $Y=0.81 $X2=0 $Y2=0
cc_684 N_S[0]_c_701_n N_VGND_c_2933_n 0.00585385f $X=5.795 $Y=0.735 $X2=0 $Y2=0
cc_685 N_S[0]_c_687_n VGND 0.00642387f $X=3.165 $Y=0.18 $X2=0 $Y2=0
cc_686 N_S[0]_c_688_n VGND 0.00591981f $X=2.895 $Y=0.18 $X2=0 $Y2=0
cc_687 N_S[0]_c_690_n VGND 0.0064237f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_688 N_S[0]_c_692_n VGND 0.00642387f $X=4.005 $Y=0.18 $X2=0 $Y2=0
cc_689 N_S[0]_c_694_n VGND 0.0345801f $X=4.765 $Y=0.18 $X2=0 $Y2=0
cc_690 N_S[0]_c_699_n VGND 0.00990284f $X=5.375 $Y=0.735 $X2=0 $Y2=0
cc_691 N_S[0]_c_701_n VGND 0.0119653f $X=5.795 $Y=0.735 $X2=0 $Y2=0
cc_692 N_S[0]_c_703_n VGND 0.00366655f $X=3.24 $Y=0.18 $X2=0 $Y2=0
cc_693 N_S[0]_c_704_n VGND 0.00366655f $X=3.66 $Y=0.18 $X2=0 $Y2=0
cc_694 N_S[0]_c_705_n VGND 0.00366655f $X=4.08 $Y=0.18 $X2=0 $Y2=0
cc_695 N_S[0]_c_686_n N_A_119_47#_c_3247_n 0.00206084f $X=2.82 $Y=0.255 $X2=0
+ $Y2=0
cc_696 N_S[0]_c_686_n N_A_119_47#_c_3249_n 0.0139014f $X=2.82 $Y=0.255 $X2=0
+ $Y2=0
cc_697 N_S[0]_c_687_n N_A_119_47#_c_3249_n 0.00211351f $X=3.165 $Y=0.18 $X2=0
+ $Y2=0
cc_698 N_S[0]_c_689_n N_A_119_47#_c_3249_n 0.0106826f $X=3.24 $Y=0.255 $X2=0
+ $Y2=0
cc_699 N_S[0]_c_691_n N_A_119_47#_c_3251_n 0.0106844f $X=3.66 $Y=0.255 $X2=0
+ $Y2=0
cc_700 N_S[0]_c_692_n N_A_119_47#_c_3251_n 0.00211351f $X=4.005 $Y=0.18 $X2=0
+ $Y2=0
cc_701 N_S[0]_c_693_n N_A_119_47#_c_3251_n 0.0112916f $X=4.08 $Y=0.255 $X2=0
+ $Y2=0
cc_702 N_S[0]_c_694_n N_A_119_47#_c_3251_n 0.00685838f $X=4.765 $Y=0.18 $X2=0
+ $Y2=0
cc_703 N_S[0]_c_695_n N_A_119_47#_c_3251_n 0.00189496f $X=4.84 $Y=0.735 $X2=0
+ $Y2=0
cc_704 N_S[0]_c_695_n N_A_119_47#_c_3252_n 0.00529837f $X=4.84 $Y=0.735 $X2=0
+ $Y2=0
cc_705 N_S[0]_c_690_n N_A_119_47#_c_3287_n 0.0034777f $X=3.585 $Y=0.18 $X2=0
+ $Y2=0
cc_706 N_S[1]_c_811_n N_A_1430_325#_c_927_n 0.00507688f $X=8.8 $Y=0.255 $X2=0
+ $Y2=0
cc_707 N_S[1]_c_806_n N_A_1430_325#_c_919_n 0.00262132f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_708 N_S[1]_c_813_n N_A_1430_325#_c_930_n 0.00509204f $X=9.22 $Y=0.255 $X2=0
+ $Y2=0
cc_709 N_S[1]_c_817_n N_A_1430_325#_c_932_n 0.00507426f $X=10.06 $Y=0.255 $X2=0
+ $Y2=0
cc_710 N_S[1]_c_815_n N_A_1430_325#_c_935_n 0.00509391f $X=9.64 $Y=0.255 $X2=0
+ $Y2=0
cc_711 N_S[1]_c_802_n N_A_1430_325#_c_936_n 0.0128955f $X=7.06 $Y=1.55 $X2=0
+ $Y2=0
cc_712 N_S[1]_c_826_n N_A_1430_325#_c_936_n 0.0118819f $X=7.53 $Y=1.55 $X2=0
+ $Y2=0
cc_713 N_S[1]_c_803_n N_A_1430_325#_c_920_n 0.00207203f $X=7.085 $Y=0.735 $X2=0
+ $Y2=0
cc_714 N_S[1]_c_805_n N_A_1430_325#_c_920_n 0.00603996f $X=7.505 $Y=0.735 $X2=0
+ $Y2=0
cc_715 N_S[1]_c_808_n N_A_1430_325#_c_920_n 6.53442e-19 $X=8.04 $Y=0.735 $X2=0
+ $Y2=0
cc_716 N_S[1]_c_802_n N_A_1430_325#_c_921_n 0.00289358f $X=7.06 $Y=1.55 $X2=0
+ $Y2=0
cc_717 N_S[1]_c_804_n N_A_1430_325#_c_921_n 0.00429801f $X=7.43 $Y=0.81 $X2=0
+ $Y2=0
cc_718 N_S[1]_c_806_n N_A_1430_325#_c_921_n 0.0085951f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_719 N_S[1]_c_818_n N_A_1430_325#_c_921_n 0.00268644f $X=7.53 $Y=0.81 $X2=0
+ $Y2=0
cc_720 N_S[1]_c_822_n N_A_1430_325#_c_921_n 0.00541767f $X=7.02 $Y=1.16 $X2=0
+ $Y2=0
cc_721 N_S[1]_c_806_n N_A_1430_325#_c_922_n 0.0206368f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_722 N_S[1]_c_807_n N_A_1430_325#_c_922_n 0.0103812f $X=7.965 $Y=0.81 $X2=0
+ $Y2=0
cc_723 N_S[1]_c_802_n N_A_1430_325#_c_938_n 0.00454075f $X=7.06 $Y=1.55 $X2=0
+ $Y2=0
cc_724 N_S[1]_c_806_n N_A_1430_325#_c_938_n 0.00255921f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_725 N_S[1]_c_826_n N_A_1430_325#_c_938_n 0.00762115f $X=7.53 $Y=1.55 $X2=0
+ $Y2=0
cc_726 N_S[1]_c_804_n N_A_1430_325#_c_923_n 0.0111895f $X=7.43 $Y=0.81 $X2=0
+ $Y2=0
cc_727 N_S[1]_c_805_n N_A_1430_325#_c_923_n 9.67113e-19 $X=7.505 $Y=0.735 $X2=0
+ $Y2=0
cc_728 N_S[1]_c_818_n N_A_1430_325#_c_923_n 0.00426435f $X=7.53 $Y=0.81 $X2=0
+ $Y2=0
cc_729 N_S[1]_c_802_n N_A_1430_325#_c_924_n 0.00416423f $X=7.06 $Y=1.55 $X2=0
+ $Y2=0
cc_730 N_S[1]_c_806_n N_A_1430_325#_c_924_n 0.00322131f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_731 N_S[1]_c_822_n N_A_1430_325#_c_924_n 0.0228692f $X=7.02 $Y=1.16 $X2=0
+ $Y2=0
cc_732 N_S[1]_c_806_n N_A_1430_325#_c_925_n 0.0175393f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_733 N_S[1]_c_807_n N_A_1430_325#_c_925_n 0.0179529f $X=7.965 $Y=0.81 $X2=0
+ $Y2=0
cc_734 N_S[1]_c_801_n N_VPWR_c_1765_n 0.00652399f $X=6.96 $Y=1.16 $X2=0 $Y2=0
cc_735 N_S[1]_c_802_n N_VPWR_c_1765_n 0.00986205f $X=7.06 $Y=1.55 $X2=0 $Y2=0
cc_736 N_S[1]_c_822_n N_VPWR_c_1765_n 0.0157609f $X=7.02 $Y=1.16 $X2=0 $Y2=0
cc_737 N_S[1]_c_826_n N_VPWR_c_1766_n 0.00950399f $X=7.53 $Y=1.55 $X2=0 $Y2=0
cc_738 N_S[1]_c_802_n N_VPWR_c_1788_n 0.00673617f $X=7.06 $Y=1.55 $X2=0 $Y2=0
cc_739 N_S[1]_c_826_n N_VPWR_c_1788_n 0.00673617f $X=7.53 $Y=1.55 $X2=0 $Y2=0
cc_740 N_S[1]_c_802_n VPWR 0.00846723f $X=7.06 $Y=1.55 $X2=0 $Y2=0
cc_741 N_S[1]_c_826_n VPWR 0.00852996f $X=7.53 $Y=1.55 $X2=0 $Y2=0
cc_742 N_S[1]_c_811_n N_Z_c_2194_n 0.0134253f $X=8.8 $Y=0.255 $X2=0 $Y2=0
cc_743 N_S[1]_c_813_n N_Z_c_2194_n 0.0077801f $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_744 N_S[1]_c_815_n N_Z_c_2194_n 6.35774e-19 $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_745 N_S[1]_c_813_n N_Z_c_2195_n 0.00190704f $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_746 N_S[1]_c_815_n N_Z_c_2195_n 3.10191e-19 $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_747 N_S[1]_c_815_n N_Z_c_2196_n 0.00283489f $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_748 N_S[1]_c_817_n N_Z_c_2196_n 0.002324f $X=10.06 $Y=0.255 $X2=0 $Y2=0
cc_749 N_S[1]_c_811_n N_Z_c_2206_n 0.00216436f $X=8.8 $Y=0.255 $X2=0 $Y2=0
cc_750 N_S[1]_c_815_n N_Z_c_2207_n 0.00180363f $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_751 N_S[1]_c_813_n N_Z_c_2208_n 6.35664e-19 $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_752 N_S[1]_c_815_n N_Z_c_2208_n 0.00462308f $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_753 N_S[1]_c_817_n N_Z_c_2208_n 0.00443615f $X=10.06 $Y=0.255 $X2=0 $Y2=0
cc_754 N_S[1]_c_801_n N_Z_c_2219_n 0.00234109f $X=6.96 $Y=1.16 $X2=0 $Y2=0
cc_755 N_S[1]_c_802_n N_Z_c_2219_n 0.0052507f $X=7.06 $Y=1.55 $X2=0 $Y2=0
cc_756 N_S[1]_c_826_n N_Z_c_2219_n 0.00478771f $X=7.53 $Y=1.55 $X2=0 $Y2=0
cc_757 N_S[1]_c_822_n N_Z_c_2219_n 0.0105931f $X=7.02 $Y=1.16 $X2=0 $Y2=0
cc_758 N_S[1]_c_826_n N_A_1643_311#_c_2607_n 0.00209354f $X=7.53 $Y=1.55 $X2=0
+ $Y2=0
cc_759 N_S[1]_c_817_n N_A_1643_311#_c_2614_n 0.00168571f $X=10.06 $Y=0.255 $X2=0
+ $Y2=0
cc_760 N_S[1]_c_801_n N_VGND_c_2913_n 0.00576464f $X=6.96 $Y=1.16 $X2=0 $Y2=0
cc_761 N_S[1]_c_803_n N_VGND_c_2913_n 0.00374526f $X=7.085 $Y=0.735 $X2=0 $Y2=0
cc_762 N_S[1]_c_822_n N_VGND_c_2913_n 0.0116218f $X=7.02 $Y=1.16 $X2=0 $Y2=0
cc_763 N_S[1]_c_805_n N_VGND_c_2914_n 0.00173127f $X=7.505 $Y=0.735 $X2=0 $Y2=0
cc_764 N_S[1]_c_807_n N_VGND_c_2914_n 0.00525833f $X=7.965 $Y=0.81 $X2=0 $Y2=0
cc_765 N_S[1]_c_810_n N_VGND_c_2914_n 0.00862298f $X=8.115 $Y=0.18 $X2=0 $Y2=0
cc_766 N_S[1]_c_816_n N_VGND_c_2915_n 0.0028166f $X=9.985 $Y=0.18 $X2=0 $Y2=0
cc_767 N_S[1]_c_817_n N_VGND_c_2915_n 5.5039e-19 $X=10.06 $Y=0.255 $X2=0 $Y2=0
cc_768 N_S[1]_c_803_n N_VGND_c_2937_n 0.00585385f $X=7.085 $Y=0.735 $X2=0 $Y2=0
cc_769 N_S[1]_c_804_n N_VGND_c_2937_n 2.16067e-19 $X=7.43 $Y=0.81 $X2=0 $Y2=0
cc_770 N_S[1]_c_805_n N_VGND_c_2937_n 0.00542362f $X=7.505 $Y=0.735 $X2=0 $Y2=0
cc_771 N_S[1]_c_810_n N_VGND_c_2939_n 0.0559651f $X=8.115 $Y=0.18 $X2=0 $Y2=0
cc_772 N_S[1]_c_803_n VGND 0.0119653f $X=7.085 $Y=0.735 $X2=0 $Y2=0
cc_773 N_S[1]_c_805_n VGND 0.00990284f $X=7.505 $Y=0.735 $X2=0 $Y2=0
cc_774 N_S[1]_c_809_n VGND 0.0244174f $X=8.725 $Y=0.18 $X2=0 $Y2=0
cc_775 N_S[1]_c_810_n VGND 0.0101627f $X=8.115 $Y=0.18 $X2=0 $Y2=0
cc_776 N_S[1]_c_812_n VGND 0.00642387f $X=9.145 $Y=0.18 $X2=0 $Y2=0
cc_777 N_S[1]_c_814_n VGND 0.0064237f $X=9.565 $Y=0.18 $X2=0 $Y2=0
cc_778 N_S[1]_c_816_n VGND 0.0123437f $X=9.985 $Y=0.18 $X2=0 $Y2=0
cc_779 N_S[1]_c_819_n VGND 0.00366655f $X=8.8 $Y=0.18 $X2=0 $Y2=0
cc_780 N_S[1]_c_820_n VGND 0.00366655f $X=9.22 $Y=0.18 $X2=0 $Y2=0
cc_781 N_S[1]_c_821_n VGND 0.00366655f $X=9.64 $Y=0.18 $X2=0 $Y2=0
cc_782 N_S[1]_c_808_n N_A_1693_66#_c_3329_n 0.00529837f $X=8.04 $Y=0.735 $X2=0
+ $Y2=0
cc_783 N_S[1]_c_811_n N_A_1693_66#_c_3330_n 0.0112916f $X=8.8 $Y=0.255 $X2=0
+ $Y2=0
cc_784 N_S[1]_c_812_n N_A_1693_66#_c_3330_n 0.00211351f $X=9.145 $Y=0.18 $X2=0
+ $Y2=0
cc_785 N_S[1]_c_813_n N_A_1693_66#_c_3330_n 0.0106844f $X=9.22 $Y=0.255 $X2=0
+ $Y2=0
cc_786 N_S[1]_c_808_n N_A_1693_66#_c_3331_n 0.00189496f $X=8.04 $Y=0.735 $X2=0
+ $Y2=0
cc_787 N_S[1]_c_809_n N_A_1693_66#_c_3331_n 0.00685838f $X=8.725 $Y=0.18 $X2=0
+ $Y2=0
cc_788 N_S[1]_c_815_n N_A_1693_66#_c_3332_n 0.0106826f $X=9.64 $Y=0.255 $X2=0
+ $Y2=0
cc_789 N_S[1]_c_816_n N_A_1693_66#_c_3332_n 0.00211351f $X=9.985 $Y=0.18 $X2=0
+ $Y2=0
cc_790 N_S[1]_c_817_n N_A_1693_66#_c_3332_n 0.0139014f $X=10.06 $Y=0.255 $X2=0
+ $Y2=0
cc_791 N_S[1]_c_817_n N_A_1693_66#_c_3335_n 0.00206084f $X=10.06 $Y=0.255 $X2=0
+ $Y2=0
cc_792 N_S[1]_c_814_n N_A_1693_66#_c_3348_n 0.0034777f $X=9.565 $Y=0.18 $X2=0
+ $Y2=0
cc_793 N_A_1430_325#_c_936_n N_VPWR_c_1765_n 0.0356181f $X=7.295 $Y=1.77 $X2=0
+ $Y2=0
cc_794 N_A_1430_325#_c_926_n N_VPWR_c_1766_n 0.00279288f $X=8.575 $Y=1.475 $X2=0
+ $Y2=0
cc_795 N_A_1430_325#_c_936_n N_VPWR_c_1766_n 0.0316788f $X=7.295 $Y=1.77 $X2=0
+ $Y2=0
cc_796 N_A_1430_325#_c_922_n N_VPWR_c_1766_n 0.0193185f $X=8.345 $Y=1.23 $X2=0
+ $Y2=0
cc_797 N_A_1430_325#_c_925_n N_VPWR_c_1766_n 6.4101e-19 $X=8.255 $Y=1.23 $X2=0
+ $Y2=0
cc_798 N_A_1430_325#_c_933_n N_VPWR_c_1767_n 0.00287722f $X=9.985 $Y=1.475 $X2=0
+ $Y2=0
cc_799 N_A_1430_325#_c_936_n N_VPWR_c_1788_n 0.0233824f $X=7.295 $Y=1.77 $X2=0
+ $Y2=0
cc_800 N_A_1430_325#_c_926_n N_VPWR_c_1790_n 0.00429453f $X=8.575 $Y=1.475 $X2=0
+ $Y2=0
cc_801 N_A_1430_325#_c_929_n N_VPWR_c_1790_n 0.00429453f $X=9.045 $Y=1.475 $X2=0
+ $Y2=0
cc_802 N_A_1430_325#_c_931_n N_VPWR_c_1790_n 0.00429453f $X=9.515 $Y=1.475 $X2=0
+ $Y2=0
cc_803 N_A_1430_325#_c_933_n N_VPWR_c_1790_n 0.00429453f $X=9.985 $Y=1.475 $X2=0
+ $Y2=0
cc_804 N_A_1430_325#_c_926_n VPWR 0.00737407f $X=8.575 $Y=1.475 $X2=0 $Y2=0
cc_805 N_A_1430_325#_c_929_n VPWR 0.0060424f $X=9.045 $Y=1.475 $X2=0 $Y2=0
cc_806 N_A_1430_325#_c_931_n VPWR 0.0060424f $X=9.515 $Y=1.475 $X2=0 $Y2=0
cc_807 N_A_1430_325#_c_933_n VPWR 0.00737407f $X=9.985 $Y=1.475 $X2=0 $Y2=0
cc_808 N_A_1430_325#_c_936_n VPWR 0.00593513f $X=7.295 $Y=1.77 $X2=0 $Y2=0
cc_809 N_A_1430_325#_c_930_n N_Z_c_2195_n 0.00762343f $X=9.425 $Y=1.4 $X2=0
+ $Y2=0
cc_810 N_A_1430_325#_c_935_n N_Z_c_2195_n 0.00704092f $X=9.515 $Y=1.4 $X2=0
+ $Y2=0
cc_811 N_A_1430_325#_c_927_n N_Z_c_2206_n 0.00597584f $X=8.955 $Y=1.4 $X2=0
+ $Y2=0
cc_812 N_A_1430_325#_c_919_n N_Z_c_2206_n 0.00747617f $X=8.665 $Y=1.4 $X2=0
+ $Y2=0
cc_813 N_A_1430_325#_c_930_n N_Z_c_2206_n 0.00145542f $X=9.425 $Y=1.4 $X2=0
+ $Y2=0
cc_814 N_A_1430_325#_c_934_n N_Z_c_2206_n 0.00909323f $X=9.045 $Y=1.4 $X2=0
+ $Y2=0
cc_815 N_A_1430_325#_c_922_n N_Z_c_2206_n 0.0266078f $X=8.345 $Y=1.23 $X2=0
+ $Y2=0
cc_816 N_A_1430_325#_c_932_n N_Z_c_2207_n 0.00918337f $X=9.895 $Y=1.4 $X2=0
+ $Y2=0
cc_817 N_A_1430_325#_c_935_n N_Z_c_2207_n 2.98555e-19 $X=9.515 $Y=1.4 $X2=0
+ $Y2=0
cc_818 N_A_1430_325#_c_932_n N_Z_c_2208_n 0.00248496f $X=9.895 $Y=1.4 $X2=0
+ $Y2=0
cc_819 N_A_1430_325#_c_926_n N_Z_c_2219_n 0.0080184f $X=8.575 $Y=1.475 $X2=0
+ $Y2=0
cc_820 N_A_1430_325#_c_919_n N_Z_c_2219_n 2.19754e-19 $X=8.665 $Y=1.4 $X2=0
+ $Y2=0
cc_821 N_A_1430_325#_c_936_n N_Z_c_2219_n 0.0329704f $X=7.295 $Y=1.77 $X2=0
+ $Y2=0
cc_822 N_A_1430_325#_c_922_n N_Z_c_2219_n 0.0186685f $X=8.345 $Y=1.23 $X2=0
+ $Y2=0
cc_823 N_A_1430_325#_c_933_n N_Z_c_2220_n 0.00841093f $X=9.985 $Y=1.475 $X2=0
+ $Y2=0
cc_824 N_A_1430_325#_c_929_n N_Z_c_2298_n 0.00378512f $X=9.045 $Y=1.475 $X2=0
+ $Y2=0
cc_825 N_A_1430_325#_c_931_n N_Z_c_2298_n 0.00378723f $X=9.515 $Y=1.475 $X2=0
+ $Y2=0
cc_826 N_A_1430_325#_c_926_n N_Z_c_2300_n 0.0107691f $X=8.575 $Y=1.475 $X2=0
+ $Y2=0
cc_827 N_A_1430_325#_c_927_n N_Z_c_2300_n 0.00554725f $X=8.955 $Y=1.4 $X2=0
+ $Y2=0
cc_828 N_A_1430_325#_c_919_n N_Z_c_2300_n 0.00415799f $X=8.665 $Y=1.4 $X2=0
+ $Y2=0
cc_829 N_A_1430_325#_c_929_n N_Z_c_2300_n 0.00814309f $X=9.045 $Y=1.475 $X2=0
+ $Y2=0
cc_830 N_A_1430_325#_c_931_n N_Z_c_2300_n 3.67612e-19 $X=9.515 $Y=1.475 $X2=0
+ $Y2=0
cc_831 N_A_1430_325#_c_934_n N_Z_c_2300_n 0.00313387f $X=9.045 $Y=1.4 $X2=0
+ $Y2=0
cc_832 N_A_1430_325#_c_922_n N_Z_c_2300_n 0.00227722f $X=8.345 $Y=1.23 $X2=0
+ $Y2=0
cc_833 N_A_1430_325#_c_929_n N_Z_c_2307_n 3.67612e-19 $X=9.045 $Y=1.475 $X2=0
+ $Y2=0
cc_834 N_A_1430_325#_c_931_n N_Z_c_2307_n 0.00814309f $X=9.515 $Y=1.475 $X2=0
+ $Y2=0
cc_835 N_A_1430_325#_c_932_n N_Z_c_2307_n 0.0102922f $X=9.895 $Y=1.4 $X2=0 $Y2=0
cc_836 N_A_1430_325#_c_933_n N_Z_c_2307_n 0.00850547f $X=9.985 $Y=1.475 $X2=0
+ $Y2=0
cc_837 N_A_1430_325#_c_935_n N_Z_c_2307_n 0.00313387f $X=9.515 $Y=1.4 $X2=0
+ $Y2=0
cc_838 N_A_1430_325#_c_926_n N_A_1643_311#_c_2607_n 0.00246857f $X=8.575
+ $Y=1.475 $X2=0 $Y2=0
cc_839 N_A_1430_325#_c_919_n N_A_1643_311#_c_2607_n 0.00561627f $X=8.665 $Y=1.4
+ $X2=0 $Y2=0
cc_840 N_A_1430_325#_c_922_n N_A_1643_311#_c_2607_n 0.0218124f $X=8.345 $Y=1.23
+ $X2=0 $Y2=0
cc_841 N_A_1430_325#_c_925_n N_A_1643_311#_c_2607_n 5.74251e-19 $X=8.255 $Y=1.23
+ $X2=0 $Y2=0
cc_842 N_A_1430_325#_c_926_n N_A_1643_311#_c_2608_n 0.0115457f $X=8.575 $Y=1.475
+ $X2=0 $Y2=0
cc_843 N_A_1430_325#_c_929_n N_A_1643_311#_c_2608_n 0.010844f $X=9.045 $Y=1.475
+ $X2=0 $Y2=0
cc_844 N_A_1430_325#_c_929_n N_A_1643_311#_c_2610_n 0.00102951f $X=9.045
+ $Y=1.475 $X2=0 $Y2=0
cc_845 N_A_1430_325#_c_930_n N_A_1643_311#_c_2610_n 0.00251792f $X=9.425 $Y=1.4
+ $X2=0 $Y2=0
cc_846 N_A_1430_325#_c_931_n N_A_1643_311#_c_2610_n 0.00102951f $X=9.515
+ $Y=1.475 $X2=0 $Y2=0
cc_847 N_A_1430_325#_c_931_n N_A_1643_311#_c_2611_n 0.010844f $X=9.515 $Y=1.475
+ $X2=0 $Y2=0
cc_848 N_A_1430_325#_c_933_n N_A_1643_311#_c_2611_n 0.0115457f $X=9.985 $Y=1.475
+ $X2=0 $Y2=0
cc_849 N_A_1430_325#_c_933_n N_A_1643_311#_c_2612_n 0.00301583f $X=9.985
+ $Y=1.475 $X2=0 $Y2=0
cc_850 N_A_1430_325#_c_933_n N_A_1643_311#_c_2614_n 0.00151141f $X=9.985
+ $Y=1.475 $X2=0 $Y2=0
cc_851 N_A_1430_325#_c_922_n N_VGND_c_2914_n 0.0123065f $X=8.345 $Y=1.23 $X2=0
+ $Y2=0
cc_852 N_A_1430_325#_c_925_n N_VGND_c_2914_n 2.04129e-19 $X=8.255 $Y=1.23 $X2=0
+ $Y2=0
cc_853 N_A_1430_325#_c_920_n N_VGND_c_2937_n 0.0129994f $X=7.295 $Y=0.445 $X2=0
+ $Y2=0
cc_854 N_A_1430_325#_M1061_s VGND 0.00394793f $X=7.16 $Y=0.235 $X2=0 $Y2=0
cc_855 N_A_1430_325#_c_920_n VGND 0.00927134f $X=7.295 $Y=0.445 $X2=0 $Y2=0
cc_856 N_A_1430_325#_c_919_n N_A_1693_66#_c_3329_n 0.00600378f $X=8.665 $Y=1.4
+ $X2=0 $Y2=0
cc_857 N_A_1430_325#_c_922_n N_A_1693_66#_c_3329_n 0.0028695f $X=8.345 $Y=1.23
+ $X2=0 $Y2=0
cc_858 N_A_1430_325#_c_930_n N_A_1693_66#_c_3351_n 7.0477e-19 $X=9.425 $Y=1.4
+ $X2=0 $Y2=0
cc_859 N_D[1]_M1001_g N_VPWR_c_1767_n 0.00369766f $X=10.975 $Y=1.985 $X2=0 $Y2=0
cc_860 N_D[1]_M1006_g N_VPWR_c_1768_n 0.00188795f $X=11.445 $Y=1.985 $X2=0 $Y2=0
cc_861 N_D[1]_M1038_g N_VPWR_c_1768_n 0.00188795f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_862 N_D[1]_M1065_g N_VPWR_c_1769_n 0.00374733f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_863 N_D[1]_M1001_g VPWR 0.00832888f $X=10.975 $Y=1.985 $X2=0 $Y2=0
cc_864 N_D[1]_M1006_g VPWR 0.00704653f $X=11.445 $Y=1.985 $X2=0 $Y2=0
cc_865 N_D[1]_M1038_g VPWR 0.00704653f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_866 N_D[1]_M1065_g VPWR 0.00832888f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_867 N_D[1]_M1001_g N_VPWR_c_1802_n 0.00673617f $X=10.975 $Y=1.985 $X2=0 $Y2=0
cc_868 N_D[1]_M1006_g N_VPWR_c_1802_n 0.00673617f $X=11.445 $Y=1.985 $X2=0 $Y2=0
cc_869 N_D[1]_M1038_g N_VPWR_c_1803_n 0.00673617f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_870 N_D[1]_M1065_g N_VPWR_c_1803_n 0.00673617f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_871 N_D[1]_M1001_g N_Z_c_2220_n 0.0041057f $X=10.975 $Y=1.985 $X2=0 $Y2=0
cc_872 N_D[1]_M1006_g N_Z_c_2220_n 0.00405638f $X=11.445 $Y=1.985 $X2=0 $Y2=0
cc_873 N_D[1]_M1038_g N_Z_c_2220_n 0.00405638f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_874 N_D[1]_M1065_g N_Z_c_2220_n 0.00470782f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_875 N_D[1]_c_1045_n N_Z_c_2220_n 0.00846955f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_876 N_D[1]_M1001_g N_A_1643_311#_c_2612_n 0.00314224f $X=10.975 $Y=1.985
+ $X2=0 $Y2=0
cc_877 N_D[1]_M1001_g N_A_1643_311#_c_2613_n 0.013247f $X=10.975 $Y=1.985 $X2=0
+ $Y2=0
cc_878 N_D[1]_M1001_g N_A_1643_311#_c_2633_n 0.0102796f $X=10.975 $Y=1.985 $X2=0
+ $Y2=0
cc_879 N_D[1]_M1006_g N_A_1643_311#_c_2633_n 0.00954371f $X=11.445 $Y=1.985
+ $X2=0 $Y2=0
cc_880 N_D[1]_M1038_g N_A_1643_311#_c_2633_n 6.58815e-19 $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_881 N_D[1]_M1006_g N_A_1643_311#_c_2636_n 0.00916655f $X=11.445 $Y=1.985
+ $X2=0 $Y2=0
cc_882 N_D[1]_M1038_g N_A_1643_311#_c_2636_n 0.00916655f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_883 N_D[1]_c_1043_n N_A_1643_311#_c_2636_n 7.15862e-19 $X=11.825 $Y=1.16
+ $X2=0 $Y2=0
cc_884 N_D[1]_c_1045_n N_A_1643_311#_c_2636_n 0.0387168f $X=12.28 $Y=1.16 $X2=0
+ $Y2=0
cc_885 N_D[1]_M1038_g N_A_1643_311#_c_2640_n 5.79575e-19 $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_886 N_D[1]_M1065_g N_A_1643_311#_c_2640_n 0.00215964f $X=12.385 $Y=1.985
+ $X2=0 $Y2=0
cc_887 N_D[1]_c_1045_n N_A_1643_311#_c_2640_n 0.0217153f $X=12.28 $Y=1.16 $X2=0
+ $Y2=0
cc_888 N_D[1]_c_1046_n N_A_1643_311#_c_2640_n 8.03631e-19 $X=12.385 $Y=1.16
+ $X2=0 $Y2=0
cc_889 N_D[1]_M1006_g N_A_1643_311#_c_2644_n 6.58815e-19 $X=11.445 $Y=1.985
+ $X2=0 $Y2=0
cc_890 N_D[1]_M1038_g N_A_1643_311#_c_2644_n 0.00954371f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_891 N_D[1]_M1065_g N_A_1643_311#_c_2644_n 0.00848227f $X=12.385 $Y=1.985
+ $X2=0 $Y2=0
cc_892 N_D[1]_M1001_g N_A_1643_311#_c_2647_n 8.61029e-19 $X=10.975 $Y=1.985
+ $X2=0 $Y2=0
cc_893 N_D[1]_M1006_g N_A_1643_311#_c_2647_n 5.79575e-19 $X=11.445 $Y=1.985
+ $X2=0 $Y2=0
cc_894 N_D[1]_c_1044_n N_A_1643_311#_c_2647_n 8.03631e-19 $X=11.535 $Y=1.16
+ $X2=0 $Y2=0
cc_895 N_D[1]_c_1045_n N_A_1643_311#_c_2647_n 0.0191156f $X=12.28 $Y=1.16 $X2=0
+ $Y2=0
cc_896 N_D[1]_M1017_g N_VGND_c_2915_n 0.00321269f $X=11 $Y=0.56 $X2=0 $Y2=0
cc_897 N_D[1]_M1029_g N_VGND_c_2915_n 2.6376e-19 $X=11.42 $Y=0.56 $X2=0 $Y2=0
cc_898 N_D[1]_M1029_g N_VGND_c_2916_n 0.0019152f $X=11.42 $Y=0.56 $X2=0 $Y2=0
cc_899 N_D[1]_M1049_g N_VGND_c_2916_n 0.00166854f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_900 N_D[1]_M1079_g N_VGND_c_2916_n 2.64031e-19 $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_901 N_D[1]_M1079_g N_VGND_c_2917_n 0.00345859f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_902 N_D[1]_M1017_g VGND 0.00702263f $X=11 $Y=0.56 $X2=0 $Y2=0
cc_903 N_D[1]_M1029_g VGND 0.00624811f $X=11.42 $Y=0.56 $X2=0 $Y2=0
cc_904 N_D[1]_M1049_g VGND 0.00593887f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_905 N_D[1]_M1079_g VGND 0.0111368f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_906 N_D[1]_M1017_g N_VGND_c_2953_n 0.00422241f $X=11 $Y=0.56 $X2=0 $Y2=0
cc_907 N_D[1]_M1029_g N_VGND_c_2953_n 0.00430643f $X=11.42 $Y=0.56 $X2=0 $Y2=0
cc_908 N_D[1]_M1049_g N_VGND_c_2954_n 0.00422241f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_909 N_D[1]_M1079_g N_VGND_c_2954_n 0.00551064f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_910 N_D[1]_M1017_g N_A_1693_66#_c_3333_n 0.00261078f $X=11 $Y=0.56 $X2=0
+ $Y2=0
cc_911 N_D[1]_M1017_g N_A_1693_66#_c_3334_n 0.0121912f $X=11 $Y=0.56 $X2=0 $Y2=0
cc_912 N_D[1]_M1017_g N_A_1693_66#_c_3354_n 0.00699463f $X=11 $Y=0.56 $X2=0
+ $Y2=0
cc_913 N_D[1]_M1029_g N_A_1693_66#_c_3354_n 0.00661764f $X=11.42 $Y=0.56 $X2=0
+ $Y2=0
cc_914 N_D[1]_M1049_g N_A_1693_66#_c_3354_n 5.22365e-19 $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_915 N_D[1]_M1029_g N_A_1693_66#_c_3336_n 0.00900364f $X=11.42 $Y=0.56 $X2=0
+ $Y2=0
cc_916 N_D[1]_M1049_g N_A_1693_66#_c_3336_n 0.00986515f $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_917 N_D[1]_M1079_g N_A_1693_66#_c_3336_n 0.00228093f $X=12.36 $Y=0.56 $X2=0
+ $Y2=0
cc_918 N_D[1]_c_1043_n N_A_1693_66#_c_3336_n 0.00463549f $X=11.825 $Y=1.16 $X2=0
+ $Y2=0
cc_919 N_D[1]_c_1045_n N_A_1693_66#_c_3336_n 0.0608884f $X=12.28 $Y=1.16 $X2=0
+ $Y2=0
cc_920 N_D[1]_c_1046_n N_A_1693_66#_c_3336_n 0.00208088f $X=12.385 $Y=1.16 $X2=0
+ $Y2=0
cc_921 N_D[1]_M1029_g N_A_1693_66#_c_3363_n 5.22365e-19 $X=11.42 $Y=0.56 $X2=0
+ $Y2=0
cc_922 N_D[1]_M1049_g N_A_1693_66#_c_3363_n 0.00661134f $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_923 N_D[1]_M1079_g N_A_1693_66#_c_3363_n 0.00529286f $X=12.36 $Y=0.56 $X2=0
+ $Y2=0
cc_924 N_D[1]_M1017_g N_A_1693_66#_c_3337_n 0.00128201f $X=11 $Y=0.56 $X2=0
+ $Y2=0
cc_925 N_D[1]_M1029_g N_A_1693_66#_c_3337_n 8.68782e-19 $X=11.42 $Y=0.56 $X2=0
+ $Y2=0
cc_926 N_D[1]_c_1044_n N_A_1693_66#_c_3337_n 0.00208088f $X=11.535 $Y=1.16 $X2=0
+ $Y2=0
cc_927 N_D[1]_c_1045_n N_A_1693_66#_c_3337_n 0.018367f $X=12.28 $Y=1.16 $X2=0
+ $Y2=0
cc_928 N_D[2]_M1005_g N_VPWR_c_1771_n 0.00374733f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_929 N_D[2]_M1019_g N_VPWR_c_1772_n 0.00188795f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_930 N_D[2]_M1047_g N_VPWR_c_1772_n 0.00188795f $X=14.315 $Y=1.985 $X2=0 $Y2=0
cc_931 N_D[2]_M1047_g N_VPWR_c_1773_n 0.00673617f $X=14.315 $Y=1.985 $X2=0 $Y2=0
cc_932 N_D[2]_M1074_g N_VPWR_c_1773_n 0.00673617f $X=14.785 $Y=1.985 $X2=0 $Y2=0
cc_933 N_D[2]_M1074_g N_VPWR_c_1774_n 0.00369766f $X=14.785 $Y=1.985 $X2=0 $Y2=0
cc_934 N_D[2]_M1005_g VPWR 0.00832888f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_935 N_D[2]_M1019_g VPWR 0.00704653f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_936 N_D[2]_M1047_g VPWR 0.00704653f $X=14.315 $Y=1.985 $X2=0 $Y2=0
cc_937 N_D[2]_M1074_g VPWR 0.00832888f $X=14.785 $Y=1.985 $X2=0 $Y2=0
cc_938 N_D[2]_M1005_g N_VPWR_c_1804_n 0.00673617f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_939 N_D[2]_M1019_g N_VPWR_c_1804_n 0.00673617f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_940 N_D[2]_M1005_g N_Z_c_2220_n 0.00470782f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_941 N_D[2]_M1019_g N_Z_c_2220_n 0.00405638f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_942 N_D[2]_M1047_g N_Z_c_2220_n 0.00405638f $X=14.315 $Y=1.985 $X2=0 $Y2=0
cc_943 N_D[2]_M1074_g N_Z_c_2220_n 0.0041057f $X=14.785 $Y=1.985 $X2=0 $Y2=0
cc_944 N_D[2]_c_1131_n N_Z_c_2220_n 0.00846955f $X=14.5 $Y=1.16 $X2=0 $Y2=0
cc_945 N_D[2]_M1005_g N_A_2693_297#_c_2720_n 0.00215964f $X=13.375 $Y=1.985
+ $X2=0 $Y2=0
cc_946 N_D[2]_M1019_g N_A_2693_297#_c_2720_n 5.79575e-19 $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_947 N_D[2]_c_1130_n N_A_2693_297#_c_2720_n 8.03631e-19 $X=13.935 $Y=1.16
+ $X2=0 $Y2=0
cc_948 N_D[2]_c_1131_n N_A_2693_297#_c_2720_n 0.0217153f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_949 N_D[2]_M1005_g N_A_2693_297#_c_2724_n 0.00848227f $X=13.375 $Y=1.985
+ $X2=0 $Y2=0
cc_950 N_D[2]_M1019_g N_A_2693_297#_c_2724_n 0.00954371f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_951 N_D[2]_M1047_g N_A_2693_297#_c_2724_n 6.58815e-19 $X=14.315 $Y=1.985
+ $X2=0 $Y2=0
cc_952 N_D[2]_M1019_g N_A_2693_297#_c_2727_n 0.00916655f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_953 N_D[2]_M1047_g N_A_2693_297#_c_2727_n 0.00916655f $X=14.315 $Y=1.985
+ $X2=0 $Y2=0
cc_954 N_D[2]_c_1129_n N_A_2693_297#_c_2727_n 7.15862e-19 $X=14.225 $Y=1.16
+ $X2=0 $Y2=0
cc_955 N_D[2]_c_1131_n N_A_2693_297#_c_2727_n 0.0387168f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_956 N_D[2]_M1019_g N_A_2693_297#_c_2731_n 6.58815e-19 $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_957 N_D[2]_M1047_g N_A_2693_297#_c_2731_n 0.00954371f $X=14.315 $Y=1.985
+ $X2=0 $Y2=0
cc_958 N_D[2]_M1074_g N_A_2693_297#_c_2731_n 0.0102796f $X=14.785 $Y=1.985 $X2=0
+ $Y2=0
cc_959 N_D[2]_M1074_g N_A_2693_297#_c_2712_n 0.013247f $X=14.785 $Y=1.985 $X2=0
+ $Y2=0
cc_960 N_D[2]_M1074_g N_A_2693_297#_c_2713_n 0.00314224f $X=14.785 $Y=1.985
+ $X2=0 $Y2=0
cc_961 N_D[2]_M1047_g N_A_2693_297#_c_2736_n 5.79575e-19 $X=14.315 $Y=1.985
+ $X2=0 $Y2=0
cc_962 N_D[2]_M1074_g N_A_2693_297#_c_2736_n 8.61029e-19 $X=14.785 $Y=1.985
+ $X2=0 $Y2=0
cc_963 N_D[2]_c_1131_n N_A_2693_297#_c_2736_n 0.0191156f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_964 N_D[2]_c_1132_n N_A_2693_297#_c_2736_n 8.03631e-19 $X=14.785 $Y=1.16
+ $X2=0 $Y2=0
cc_965 N_D[2]_M1002_g N_VGND_c_2919_n 0.00345859f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_966 N_D[2]_M1002_g N_VGND_c_2920_n 2.64031e-19 $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_967 N_D[2]_M1021_g N_VGND_c_2920_n 0.00166854f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_968 N_D[2]_M1034_g N_VGND_c_2920_n 0.0019152f $X=14.34 $Y=0.56 $X2=0 $Y2=0
cc_969 N_D[2]_M1034_g N_VGND_c_2921_n 0.00430643f $X=14.34 $Y=0.56 $X2=0 $Y2=0
cc_970 N_D[2]_M1052_g N_VGND_c_2921_n 0.00422241f $X=14.76 $Y=0.56 $X2=0 $Y2=0
cc_971 N_D[2]_M1034_g N_VGND_c_2922_n 2.6376e-19 $X=14.34 $Y=0.56 $X2=0 $Y2=0
cc_972 N_D[2]_M1052_g N_VGND_c_2922_n 0.00321269f $X=14.76 $Y=0.56 $X2=0 $Y2=0
cc_973 N_D[2]_M1002_g VGND 0.0111368f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_974 N_D[2]_M1021_g VGND 0.00593887f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_975 N_D[2]_M1034_g VGND 0.00624811f $X=14.34 $Y=0.56 $X2=0 $Y2=0
cc_976 N_D[2]_M1052_g VGND 0.00702263f $X=14.76 $Y=0.56 $X2=0 $Y2=0
cc_977 N_D[2]_M1002_g N_VGND_c_2955_n 0.00551064f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_978 N_D[2]_M1021_g N_VGND_c_2955_n 0.00422241f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_979 N_D[2]_M1002_g N_A_2695_47#_c_3421_n 0.00529286f $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_980 N_D[2]_M1021_g N_A_2695_47#_c_3421_n 0.00661134f $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_981 N_D[2]_M1034_g N_A_2695_47#_c_3421_n 5.22365e-19 $X=14.34 $Y=0.56 $X2=0
+ $Y2=0
cc_982 N_D[2]_M1021_g N_A_2695_47#_c_3424_n 0.00899636f $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_983 N_D[2]_M1034_g N_A_2695_47#_c_3424_n 0.00900364f $X=14.34 $Y=0.56 $X2=0
+ $Y2=0
cc_984 N_D[2]_c_1129_n N_A_2695_47#_c_3424_n 0.00463549f $X=14.225 $Y=1.16 $X2=0
+ $Y2=0
cc_985 N_D[2]_c_1131_n N_A_2695_47#_c_3424_n 0.0394855f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_986 N_D[2]_M1002_g N_A_2695_47#_c_3413_n 0.00228093f $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_987 N_D[2]_M1021_g N_A_2695_47#_c_3413_n 8.68782e-19 $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_988 N_D[2]_c_1130_n N_A_2695_47#_c_3413_n 0.00208088f $X=13.935 $Y=1.16 $X2=0
+ $Y2=0
cc_989 N_D[2]_c_1131_n N_A_2695_47#_c_3413_n 0.021403f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_990 N_D[2]_M1021_g N_A_2695_47#_c_3432_n 5.22365e-19 $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_991 N_D[2]_M1034_g N_A_2695_47#_c_3432_n 0.00661764f $X=14.34 $Y=0.56 $X2=0
+ $Y2=0
cc_992 N_D[2]_M1052_g N_A_2695_47#_c_3432_n 0.00699463f $X=14.76 $Y=0.56 $X2=0
+ $Y2=0
cc_993 N_D[2]_M1052_g N_A_2695_47#_c_3414_n 0.0121912f $X=14.76 $Y=0.56 $X2=0
+ $Y2=0
cc_994 N_D[2]_M1052_g N_A_2695_47#_c_3415_n 0.00261078f $X=14.76 $Y=0.56 $X2=0
+ $Y2=0
cc_995 N_D[2]_M1034_g N_A_2695_47#_c_3420_n 8.68782e-19 $X=14.34 $Y=0.56 $X2=0
+ $Y2=0
cc_996 N_D[2]_M1052_g N_A_2695_47#_c_3420_n 0.00128201f $X=14.76 $Y=0.56 $X2=0
+ $Y2=0
cc_997 N_D[2]_c_1131_n N_A_2695_47#_c_3420_n 0.018367f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_998 N_D[2]_c_1132_n N_A_2695_47#_c_3420_n 0.00208088f $X=14.785 $Y=1.16 $X2=0
+ $Y2=0
cc_999 N_A_3135_265#_c_1218_n N_S[2]_c_1328_n 0.00507426f $X=15.865 $Y=1.4
+ $X2=-0.19 $Y2=-0.24
cc_1000 N_A_3135_265#_c_1217_n N_S[2]_c_1331_n 0.00509391f $X=16.155 $Y=1.4
+ $X2=0 $Y2=0
cc_1001 N_A_3135_265#_c_1220_n N_S[2]_c_1333_n 0.00509204f $X=16.625 $Y=1.4
+ $X2=0 $Y2=0
cc_1002 N_A_3135_265#_c_1222_n N_S[2]_c_1335_n 0.00507688f $X=17.095 $Y=1.4
+ $X2=0 $Y2=0
cc_1003 N_A_3135_265#_c_1211_n N_S[2]_c_1337_n 6.53442e-19 $X=18.465 $Y=0.445
+ $X2=0 $Y2=0
cc_1004 N_A_3135_265#_c_1209_n N_S[2]_c_1339_n 0.0103812f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_1005 N_A_3135_265#_c_1210_n N_S[2]_c_1339_n 0.0179529f $X=17.755 $Y=1.23
+ $X2=0 $Y2=0
cc_1006 N_A_3135_265#_c_1209_n N_S[2]_c_1340_n 0.0206368f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_1007 N_A_3135_265#_c_1210_n N_S[2]_c_1340_n 0.0175393f $X=17.755 $Y=1.23
+ $X2=0 $Y2=0
cc_1008 N_A_3135_265#_c_1212_n N_S[2]_c_1340_n 0.0085951f $X=18.385 $Y=1.065
+ $X2=0 $Y2=0
cc_1009 N_A_3135_265#_c_1214_n N_S[2]_c_1340_n 0.00322131f $X=18.385 $Y=1.23
+ $X2=0 $Y2=0
cc_1010 N_A_3135_265#_c_1230_n N_S[2]_c_1340_n 0.00255921f $X=18.465 $Y=1.605
+ $X2=0 $Y2=0
cc_1011 N_A_3135_265#_c_1215_n N_S[2]_c_1340_n 0.00262132f $X=17.505 $Y=1.23
+ $X2=0 $Y2=0
cc_1012 N_A_3135_265#_c_1228_n N_S[2]_c_1351_n 0.0118819f $X=18.465 $Y=1.77
+ $X2=0 $Y2=0
cc_1013 N_A_3135_265#_c_1230_n N_S[2]_c_1351_n 0.00762115f $X=18.465 $Y=1.605
+ $X2=0 $Y2=0
cc_1014 N_A_3135_265#_c_1211_n N_S[2]_c_1341_n 0.00603996f $X=18.465 $Y=0.445
+ $X2=0 $Y2=0
cc_1015 N_A_3135_265#_c_1213_n N_S[2]_c_1341_n 9.67113e-19 $X=18.425 $Y=0.825
+ $X2=0 $Y2=0
cc_1016 N_A_3135_265#_c_1212_n N_S[2]_c_1342_n 0.00429801f $X=18.385 $Y=1.065
+ $X2=0 $Y2=0
cc_1017 N_A_3135_265#_c_1213_n N_S[2]_c_1342_n 0.0111895f $X=18.425 $Y=0.825
+ $X2=0 $Y2=0
cc_1018 N_A_3135_265#_c_1211_n N_S[2]_c_1343_n 0.00207203f $X=18.465 $Y=0.445
+ $X2=0 $Y2=0
cc_1019 N_A_3135_265#_c_1212_n N_S[2]_c_1344_n 0.00289358f $X=18.385 $Y=1.065
+ $X2=0 $Y2=0
cc_1020 N_A_3135_265#_c_1228_n N_S[2]_c_1344_n 0.0128955f $X=18.465 $Y=1.77
+ $X2=0 $Y2=0
cc_1021 N_A_3135_265#_c_1214_n N_S[2]_c_1344_n 0.00416423f $X=18.385 $Y=1.23
+ $X2=0 $Y2=0
cc_1022 N_A_3135_265#_c_1230_n N_S[2]_c_1344_n 0.00454075f $X=18.465 $Y=1.605
+ $X2=0 $Y2=0
cc_1023 N_A_3135_265#_c_1212_n N_S[2]_c_1348_n 0.00268644f $X=18.385 $Y=1.065
+ $X2=0 $Y2=0
cc_1024 N_A_3135_265#_c_1213_n N_S[2]_c_1348_n 0.00426435f $X=18.425 $Y=0.825
+ $X2=0 $Y2=0
cc_1025 N_A_3135_265#_c_1212_n S[2] 0.00541767f $X=18.385 $Y=1.065 $X2=0 $Y2=0
cc_1026 N_A_3135_265#_c_1214_n S[2] 0.0228692f $X=18.385 $Y=1.23 $X2=0 $Y2=0
cc_1027 N_A_3135_265#_c_1216_n N_VPWR_c_1774_n 0.00287722f $X=15.775 $Y=1.475
+ $X2=0 $Y2=0
cc_1028 N_A_3135_265#_c_1223_n N_VPWR_c_1775_n 0.00279288f $X=17.185 $Y=1.475
+ $X2=0 $Y2=0
cc_1029 N_A_3135_265#_c_1209_n N_VPWR_c_1775_n 0.0193185f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_1030 N_A_3135_265#_c_1210_n N_VPWR_c_1775_n 6.4101e-19 $X=17.755 $Y=1.23
+ $X2=0 $Y2=0
cc_1031 N_A_3135_265#_c_1228_n N_VPWR_c_1775_n 0.0316788f $X=18.465 $Y=1.77
+ $X2=0 $Y2=0
cc_1032 N_A_3135_265#_c_1228_n N_VPWR_c_1776_n 0.0356181f $X=18.465 $Y=1.77
+ $X2=0 $Y2=0
cc_1033 N_A_3135_265#_c_1216_n N_VPWR_c_1792_n 0.00429453f $X=15.775 $Y=1.475
+ $X2=0 $Y2=0
cc_1034 N_A_3135_265#_c_1219_n N_VPWR_c_1792_n 0.00429453f $X=16.245 $Y=1.475
+ $X2=0 $Y2=0
cc_1035 N_A_3135_265#_c_1221_n N_VPWR_c_1792_n 0.00429453f $X=16.715 $Y=1.475
+ $X2=0 $Y2=0
cc_1036 N_A_3135_265#_c_1223_n N_VPWR_c_1792_n 0.00429453f $X=17.185 $Y=1.475
+ $X2=0 $Y2=0
cc_1037 N_A_3135_265#_c_1228_n N_VPWR_c_1794_n 0.0233824f $X=18.465 $Y=1.77
+ $X2=0 $Y2=0
cc_1038 N_A_3135_265#_c_1216_n VPWR 0.00737407f $X=15.775 $Y=1.475 $X2=0 $Y2=0
cc_1039 N_A_3135_265#_c_1219_n VPWR 0.0060424f $X=16.245 $Y=1.475 $X2=0 $Y2=0
cc_1040 N_A_3135_265#_c_1221_n VPWR 0.0060424f $X=16.715 $Y=1.475 $X2=0 $Y2=0
cc_1041 N_A_3135_265#_c_1223_n VPWR 0.00737407f $X=17.185 $Y=1.475 $X2=0 $Y2=0
cc_1042 N_A_3135_265#_c_1228_n VPWR 0.00593513f $X=18.465 $Y=1.77 $X2=0 $Y2=0
cc_1043 N_A_3135_265#_c_1220_n N_Z_c_2198_n 0.00762343f $X=16.625 $Y=1.4 $X2=0
+ $Y2=0
cc_1044 N_A_3135_265#_c_1224_n N_Z_c_2198_n 0.00704092f $X=16.245 $Y=1.4 $X2=0
+ $Y2=0
cc_1045 N_A_3135_265#_c_1218_n N_Z_c_2209_n 0.00248496f $X=15.865 $Y=1.4 $X2=0
+ $Y2=0
cc_1046 N_A_3135_265#_c_1217_n N_Z_c_2210_n 0.00678861f $X=16.155 $Y=1.4 $X2=0
+ $Y2=0
cc_1047 N_A_3135_265#_c_1218_n N_Z_c_2210_n 0.00239476f $X=15.865 $Y=1.4 $X2=0
+ $Y2=0
cc_1048 N_A_3135_265#_c_1224_n N_Z_c_2210_n 2.98555e-19 $X=16.245 $Y=1.4 $X2=0
+ $Y2=0
cc_1049 N_A_3135_265#_c_1220_n N_Z_c_2211_n 0.00145542f $X=16.625 $Y=1.4 $X2=0
+ $Y2=0
cc_1050 N_A_3135_265#_c_1222_n N_Z_c_2211_n 0.00597584f $X=17.095 $Y=1.4 $X2=0
+ $Y2=0
cc_1051 N_A_3135_265#_c_1225_n N_Z_c_2211_n 0.00909323f $X=16.715 $Y=1.4 $X2=0
+ $Y2=0
cc_1052 N_A_3135_265#_c_1209_n N_Z_c_2211_n 0.0266078f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_1053 N_A_3135_265#_c_1215_n N_Z_c_2211_n 0.00747617f $X=17.505 $Y=1.23 $X2=0
+ $Y2=0
cc_1054 N_A_3135_265#_c_1216_n N_Z_c_2220_n 0.00841093f $X=15.775 $Y=1.475 $X2=0
+ $Y2=0
cc_1055 N_A_3135_265#_c_1223_n N_Z_c_2221_n 0.0080184f $X=17.185 $Y=1.475 $X2=0
+ $Y2=0
cc_1056 N_A_3135_265#_c_1209_n N_Z_c_2221_n 0.0186685f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_1057 N_A_3135_265#_c_1228_n N_Z_c_2221_n 0.0329704f $X=18.465 $Y=1.77 $X2=0
+ $Y2=0
cc_1058 N_A_3135_265#_c_1215_n N_Z_c_2221_n 2.19754e-19 $X=17.505 $Y=1.23 $X2=0
+ $Y2=0
cc_1059 N_A_3135_265#_c_1219_n Z 0.00378723f $X=16.245 $Y=1.475 $X2=0 $Y2=0
cc_1060 N_A_3135_265#_c_1221_n Z 0.00378512f $X=16.715 $Y=1.475 $X2=0 $Y2=0
cc_1061 N_A_3135_265#_c_1216_n N_Z_c_2340_n 0.00850547f $X=15.775 $Y=1.475 $X2=0
+ $Y2=0
cc_1062 N_A_3135_265#_c_1217_n N_Z_c_2340_n 0.00554725f $X=16.155 $Y=1.4 $X2=0
+ $Y2=0
cc_1063 N_A_3135_265#_c_1218_n N_Z_c_2340_n 0.00474497f $X=15.865 $Y=1.4 $X2=0
+ $Y2=0
cc_1064 N_A_3135_265#_c_1219_n N_Z_c_2340_n 0.00814309f $X=16.245 $Y=1.475 $X2=0
+ $Y2=0
cc_1065 N_A_3135_265#_c_1221_n N_Z_c_2340_n 3.67612e-19 $X=16.715 $Y=1.475 $X2=0
+ $Y2=0
cc_1066 N_A_3135_265#_c_1224_n N_Z_c_2340_n 0.00313387f $X=16.245 $Y=1.4 $X2=0
+ $Y2=0
cc_1067 N_A_3135_265#_c_1219_n N_Z_c_2346_n 3.67612e-19 $X=16.245 $Y=1.475 $X2=0
+ $Y2=0
cc_1068 N_A_3135_265#_c_1221_n N_Z_c_2346_n 0.00814309f $X=16.715 $Y=1.475 $X2=0
+ $Y2=0
cc_1069 N_A_3135_265#_c_1222_n N_Z_c_2346_n 0.00554725f $X=17.095 $Y=1.4 $X2=0
+ $Y2=0
cc_1070 N_A_3135_265#_c_1223_n N_Z_c_2346_n 0.0107691f $X=17.185 $Y=1.475 $X2=0
+ $Y2=0
cc_1071 N_A_3135_265#_c_1225_n N_Z_c_2346_n 0.00313387f $X=16.715 $Y=1.4 $X2=0
+ $Y2=0
cc_1072 N_A_3135_265#_c_1209_n N_Z_c_2346_n 0.00227722f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_1073 N_A_3135_265#_c_1215_n N_Z_c_2346_n 0.00415799f $X=17.505 $Y=1.23 $X2=0
+ $Y2=0
cc_1074 N_A_3135_265#_c_1216_n N_A_2693_297#_c_2712_n 0.00151141f $X=15.775
+ $Y=1.475 $X2=0 $Y2=0
cc_1075 N_A_3135_265#_c_1216_n N_A_2693_297#_c_2713_n 0.00301583f $X=15.775
+ $Y=1.475 $X2=0 $Y2=0
cc_1076 N_A_3135_265#_c_1216_n N_A_2693_297#_c_2714_n 0.0115457f $X=15.775
+ $Y=1.475 $X2=0 $Y2=0
cc_1077 N_A_3135_265#_c_1219_n N_A_2693_297#_c_2714_n 0.010844f $X=16.245
+ $Y=1.475 $X2=0 $Y2=0
cc_1078 N_A_3135_265#_c_1219_n N_A_2693_297#_c_2716_n 0.00102951f $X=16.245
+ $Y=1.475 $X2=0 $Y2=0
cc_1079 N_A_3135_265#_c_1220_n N_A_2693_297#_c_2716_n 0.00251792f $X=16.625
+ $Y=1.4 $X2=0 $Y2=0
cc_1080 N_A_3135_265#_c_1221_n N_A_2693_297#_c_2716_n 0.00102951f $X=16.715
+ $Y=1.475 $X2=0 $Y2=0
cc_1081 N_A_3135_265#_c_1221_n N_A_2693_297#_c_2717_n 0.010844f $X=16.715
+ $Y=1.475 $X2=0 $Y2=0
cc_1082 N_A_3135_265#_c_1223_n N_A_2693_297#_c_2717_n 0.0115457f $X=17.185
+ $Y=1.475 $X2=0 $Y2=0
cc_1083 N_A_3135_265#_c_1223_n N_A_2693_297#_c_2718_n 0.00246857f $X=17.185
+ $Y=1.475 $X2=0 $Y2=0
cc_1084 N_A_3135_265#_c_1209_n N_A_2693_297#_c_2718_n 0.0218124f $X=18.3 $Y=1.23
+ $X2=0 $Y2=0
cc_1085 N_A_3135_265#_c_1210_n N_A_2693_297#_c_2718_n 5.74251e-19 $X=17.755
+ $Y=1.23 $X2=0 $Y2=0
cc_1086 N_A_3135_265#_c_1215_n N_A_2693_297#_c_2718_n 0.00561627f $X=17.505
+ $Y=1.23 $X2=0 $Y2=0
cc_1087 N_A_3135_265#_c_1209_n N_VGND_c_2923_n 0.0123065f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_1088 N_A_3135_265#_c_1210_n N_VGND_c_2923_n 2.04129e-19 $X=17.755 $Y=1.23
+ $X2=0 $Y2=0
cc_1089 N_A_3135_265#_c_1211_n N_VGND_c_2943_n 0.0129994f $X=18.465 $Y=0.445
+ $X2=0 $Y2=0
cc_1090 N_A_3135_265#_M1058_s VGND 0.00394793f $X=18.33 $Y=0.235 $X2=0 $Y2=0
cc_1091 N_A_3135_265#_c_1211_n VGND 0.00927134f $X=18.465 $Y=0.445 $X2=0 $Y2=0
cc_1092 N_A_3135_265#_c_1224_n N_A_2695_47#_c_3441_n 7.0477e-19 $X=16.245 $Y=1.4
+ $X2=0 $Y2=0
cc_1093 N_A_3135_265#_c_1209_n N_A_2695_47#_c_3419_n 0.0028695f $X=18.3 $Y=1.23
+ $X2=0 $Y2=0
cc_1094 N_A_3135_265#_c_1215_n N_A_2695_47#_c_3419_n 0.00589316f $X=17.505
+ $Y=1.23 $X2=0 $Y2=0
cc_1095 N_S[2]_c_1344_n N_S[3]_c_1443_n 0.0215827f $X=18.7 $Y=1.55 $X2=-0.19
+ $Y2=-0.24
cc_1096 S[2] N_S[3]_c_1443_n 0.00113563f $X=19.005 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_1097 N_S[2]_c_1344_n N_S[3]_c_1464_n 0.00113563f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_1098 S[2] N_S[3]_c_1464_n 0.0301108f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1099 N_S[2]_c_1351_n N_VPWR_c_1775_n 0.00950399f $X=18.23 $Y=1.55 $X2=0 $Y2=0
cc_1100 N_S[2]_c_1344_n N_VPWR_c_1776_n 0.016386f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_1101 S[2] N_VPWR_c_1776_n 0.0157609f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1102 N_S[2]_c_1351_n N_VPWR_c_1794_n 0.00673617f $X=18.23 $Y=1.55 $X2=0 $Y2=0
cc_1103 N_S[2]_c_1344_n N_VPWR_c_1794_n 0.00673617f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_1104 N_S[2]_c_1351_n VPWR 0.00852996f $X=18.23 $Y=1.55 $X2=0 $Y2=0
cc_1105 N_S[2]_c_1344_n VPWR 0.00846723f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_1106 N_S[2]_c_1328_n N_Z_c_2197_n 0.002324f $X=15.7 $Y=0.255 $X2=0 $Y2=0
cc_1107 N_S[2]_c_1331_n N_Z_c_2197_n 0.00283489f $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_1108 N_S[2]_c_1331_n N_Z_c_2198_n 3.10191e-19 $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_1109 N_S[2]_c_1333_n N_Z_c_2198_n 0.00190704f $X=16.54 $Y=0.255 $X2=0 $Y2=0
cc_1110 N_S[2]_c_1331_n N_Z_c_2199_n 6.35774e-19 $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_1111 N_S[2]_c_1333_n N_Z_c_2199_n 0.0077801f $X=16.54 $Y=0.255 $X2=0 $Y2=0
cc_1112 N_S[2]_c_1335_n N_Z_c_2199_n 0.0134253f $X=16.96 $Y=0.255 $X2=0 $Y2=0
cc_1113 N_S[2]_c_1328_n N_Z_c_2209_n 0.00443615f $X=15.7 $Y=0.255 $X2=0 $Y2=0
cc_1114 N_S[2]_c_1331_n N_Z_c_2209_n 0.00462308f $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_1115 N_S[2]_c_1333_n N_Z_c_2209_n 6.35664e-19 $X=16.54 $Y=0.255 $X2=0 $Y2=0
cc_1116 N_S[2]_c_1331_n N_Z_c_2210_n 0.00180363f $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_1117 N_S[2]_c_1335_n N_Z_c_2211_n 0.00216436f $X=16.96 $Y=0.255 $X2=0 $Y2=0
cc_1118 N_S[2]_c_1351_n N_Z_c_2221_n 0.00478771f $X=18.23 $Y=1.55 $X2=0 $Y2=0
cc_1119 N_S[2]_c_1344_n N_Z_c_2221_n 0.00760321f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_1120 S[2] N_Z_c_2221_n 0.010609f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1121 N_S[2]_c_1328_n N_A_2693_297#_c_2712_n 0.00168571f $X=15.7 $Y=0.255
+ $X2=0 $Y2=0
cc_1122 N_S[2]_c_1351_n N_A_2693_297#_c_2718_n 0.00209354f $X=18.23 $Y=1.55
+ $X2=0 $Y2=0
cc_1123 N_S[2]_c_1328_n N_VGND_c_2922_n 5.5039e-19 $X=15.7 $Y=0.255 $X2=0 $Y2=0
cc_1124 N_S[2]_c_1330_n N_VGND_c_2922_n 0.0028166f $X=15.775 $Y=0.18 $X2=0 $Y2=0
cc_1125 N_S[2]_c_1336_n N_VGND_c_2923_n 0.00862298f $X=17.645 $Y=0.18 $X2=0
+ $Y2=0
cc_1126 N_S[2]_c_1338_n N_VGND_c_2923_n 0.00525833f $X=18.13 $Y=0.81 $X2=0 $Y2=0
cc_1127 N_S[2]_c_1341_n N_VGND_c_2923_n 0.00173127f $X=18.255 $Y=0.735 $X2=0
+ $Y2=0
cc_1128 N_S[2]_c_1343_n N_VGND_c_2924_n 0.00374526f $X=18.675 $Y=0.735 $X2=0
+ $Y2=0
cc_1129 N_S[2]_c_1344_n N_VGND_c_2924_n 0.00578076f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_1130 S[2] N_VGND_c_2924_n 0.0116413f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_1131 N_S[2]_c_1330_n N_VGND_c_2941_n 0.0559651f $X=15.775 $Y=0.18 $X2=0 $Y2=0
cc_1132 N_S[2]_c_1341_n N_VGND_c_2943_n 0.00542362f $X=18.255 $Y=0.735 $X2=0
+ $Y2=0
cc_1133 N_S[2]_c_1342_n N_VGND_c_2943_n 2.16067e-19 $X=18.6 $Y=0.81 $X2=0 $Y2=0
cc_1134 N_S[2]_c_1343_n N_VGND_c_2943_n 0.00585385f $X=18.675 $Y=0.735 $X2=0
+ $Y2=0
cc_1135 N_S[2]_c_1329_n VGND 0.00642387f $X=16.045 $Y=0.18 $X2=0 $Y2=0
cc_1136 N_S[2]_c_1330_n VGND 0.00591981f $X=15.775 $Y=0.18 $X2=0 $Y2=0
cc_1137 N_S[2]_c_1332_n VGND 0.0064237f $X=16.465 $Y=0.18 $X2=0 $Y2=0
cc_1138 N_S[2]_c_1334_n VGND 0.00642387f $X=16.885 $Y=0.18 $X2=0 $Y2=0
cc_1139 N_S[2]_c_1336_n VGND 0.0345801f $X=17.645 $Y=0.18 $X2=0 $Y2=0
cc_1140 N_S[2]_c_1341_n VGND 0.00990284f $X=18.255 $Y=0.735 $X2=0 $Y2=0
cc_1141 N_S[2]_c_1343_n VGND 0.0119653f $X=18.675 $Y=0.735 $X2=0 $Y2=0
cc_1142 N_S[2]_c_1345_n VGND 0.00366655f $X=16.12 $Y=0.18 $X2=0 $Y2=0
cc_1143 N_S[2]_c_1346_n VGND 0.00366655f $X=16.54 $Y=0.18 $X2=0 $Y2=0
cc_1144 N_S[2]_c_1347_n VGND 0.00366655f $X=16.96 $Y=0.18 $X2=0 $Y2=0
cc_1145 N_S[2]_c_1328_n N_A_2695_47#_c_3414_n 0.00206084f $X=15.7 $Y=0.255 $X2=0
+ $Y2=0
cc_1146 N_S[2]_c_1328_n N_A_2695_47#_c_3416_n 0.0139014f $X=15.7 $Y=0.255 $X2=0
+ $Y2=0
cc_1147 N_S[2]_c_1329_n N_A_2695_47#_c_3416_n 0.00211351f $X=16.045 $Y=0.18
+ $X2=0 $Y2=0
cc_1148 N_S[2]_c_1331_n N_A_2695_47#_c_3416_n 0.0106826f $X=16.12 $Y=0.255 $X2=0
+ $Y2=0
cc_1149 N_S[2]_c_1333_n N_A_2695_47#_c_3418_n 0.0106844f $X=16.54 $Y=0.255 $X2=0
+ $Y2=0
cc_1150 N_S[2]_c_1334_n N_A_2695_47#_c_3418_n 0.00211351f $X=16.885 $Y=0.18
+ $X2=0 $Y2=0
cc_1151 N_S[2]_c_1335_n N_A_2695_47#_c_3418_n 0.0112916f $X=16.96 $Y=0.255 $X2=0
+ $Y2=0
cc_1152 N_S[2]_c_1336_n N_A_2695_47#_c_3418_n 0.00685838f $X=17.645 $Y=0.18
+ $X2=0 $Y2=0
cc_1153 N_S[2]_c_1337_n N_A_2695_47#_c_3418_n 0.00189496f $X=17.72 $Y=0.735
+ $X2=0 $Y2=0
cc_1154 N_S[2]_c_1337_n N_A_2695_47#_c_3419_n 0.00529837f $X=17.72 $Y=0.735
+ $X2=0 $Y2=0
cc_1155 N_S[2]_c_1332_n N_A_2695_47#_c_3454_n 0.0034777f $X=16.465 $Y=0.18 $X2=0
+ $Y2=0
cc_1156 N_S[3]_c_1453_n N_A_4006_325#_c_1569_n 0.00507688f $X=21.68 $Y=0.255
+ $X2=0 $Y2=0
cc_1157 N_S[3]_c_1448_n N_A_4006_325#_c_1561_n 0.00262132f $X=20.41 $Y=1.45
+ $X2=0 $Y2=0
cc_1158 N_S[3]_c_1455_n N_A_4006_325#_c_1572_n 0.00509204f $X=22.1 $Y=0.255
+ $X2=0 $Y2=0
cc_1159 N_S[3]_c_1459_n N_A_4006_325#_c_1574_n 0.00507426f $X=22.94 $Y=0.255
+ $X2=0 $Y2=0
cc_1160 N_S[3]_c_1457_n N_A_4006_325#_c_1577_n 0.00509391f $X=22.52 $Y=0.255
+ $X2=0 $Y2=0
cc_1161 N_S[3]_c_1444_n N_A_4006_325#_c_1578_n 0.0128955f $X=19.94 $Y=1.55 $X2=0
+ $Y2=0
cc_1162 N_S[3]_c_1468_n N_A_4006_325#_c_1578_n 0.0118819f $X=20.41 $Y=1.55 $X2=0
+ $Y2=0
cc_1163 N_S[3]_c_1445_n N_A_4006_325#_c_1562_n 0.00207203f $X=19.965 $Y=0.735
+ $X2=0 $Y2=0
cc_1164 N_S[3]_c_1447_n N_A_4006_325#_c_1562_n 0.00603996f $X=20.385 $Y=0.735
+ $X2=0 $Y2=0
cc_1165 N_S[3]_c_1450_n N_A_4006_325#_c_1562_n 6.53442e-19 $X=20.92 $Y=0.735
+ $X2=0 $Y2=0
cc_1166 N_S[3]_c_1444_n N_A_4006_325#_c_1563_n 0.00289358f $X=19.94 $Y=1.55
+ $X2=0 $Y2=0
cc_1167 N_S[3]_c_1446_n N_A_4006_325#_c_1563_n 0.00429801f $X=20.31 $Y=0.81
+ $X2=0 $Y2=0
cc_1168 N_S[3]_c_1448_n N_A_4006_325#_c_1563_n 0.0085951f $X=20.41 $Y=1.45 $X2=0
+ $Y2=0
cc_1169 N_S[3]_c_1460_n N_A_4006_325#_c_1563_n 0.00268644f $X=20.41 $Y=0.81
+ $X2=0 $Y2=0
cc_1170 N_S[3]_c_1464_n N_A_4006_325#_c_1563_n 0.00541767f $X=19.9 $Y=1.16 $X2=0
+ $Y2=0
cc_1171 N_S[3]_c_1448_n N_A_4006_325#_c_1564_n 0.0206368f $X=20.41 $Y=1.45 $X2=0
+ $Y2=0
cc_1172 N_S[3]_c_1449_n N_A_4006_325#_c_1564_n 0.0103812f $X=20.845 $Y=0.81
+ $X2=0 $Y2=0
cc_1173 N_S[3]_c_1444_n N_A_4006_325#_c_1580_n 0.00454075f $X=19.94 $Y=1.55
+ $X2=0 $Y2=0
cc_1174 N_S[3]_c_1448_n N_A_4006_325#_c_1580_n 0.00255921f $X=20.41 $Y=1.45
+ $X2=0 $Y2=0
cc_1175 N_S[3]_c_1468_n N_A_4006_325#_c_1580_n 0.00762115f $X=20.41 $Y=1.55
+ $X2=0 $Y2=0
cc_1176 N_S[3]_c_1446_n N_A_4006_325#_c_1565_n 0.0111895f $X=20.31 $Y=0.81 $X2=0
+ $Y2=0
cc_1177 N_S[3]_c_1447_n N_A_4006_325#_c_1565_n 9.67113e-19 $X=20.385 $Y=0.735
+ $X2=0 $Y2=0
cc_1178 N_S[3]_c_1460_n N_A_4006_325#_c_1565_n 0.00426435f $X=20.41 $Y=0.81
+ $X2=0 $Y2=0
cc_1179 N_S[3]_c_1444_n N_A_4006_325#_c_1566_n 0.00416423f $X=19.94 $Y=1.55
+ $X2=0 $Y2=0
cc_1180 N_S[3]_c_1448_n N_A_4006_325#_c_1566_n 0.00322131f $X=20.41 $Y=1.45
+ $X2=0 $Y2=0
cc_1181 N_S[3]_c_1464_n N_A_4006_325#_c_1566_n 0.0228692f $X=19.9 $Y=1.16 $X2=0
+ $Y2=0
cc_1182 N_S[3]_c_1448_n N_A_4006_325#_c_1567_n 0.0175393f $X=20.41 $Y=1.45 $X2=0
+ $Y2=0
cc_1183 N_S[3]_c_1449_n N_A_4006_325#_c_1567_n 0.0179529f $X=20.845 $Y=0.81
+ $X2=0 $Y2=0
cc_1184 N_S[3]_c_1443_n N_VPWR_c_1778_n 0.00652399f $X=19.84 $Y=1.16 $X2=0 $Y2=0
cc_1185 N_S[3]_c_1444_n N_VPWR_c_1778_n 0.00986205f $X=19.94 $Y=1.55 $X2=0 $Y2=0
cc_1186 N_S[3]_c_1464_n N_VPWR_c_1778_n 0.0157609f $X=19.9 $Y=1.16 $X2=0 $Y2=0
cc_1187 N_S[3]_c_1468_n N_VPWR_c_1779_n 0.00950399f $X=20.41 $Y=1.55 $X2=0 $Y2=0
cc_1188 N_S[3]_c_1444_n N_VPWR_c_1796_n 0.00673617f $X=19.94 $Y=1.55 $X2=0 $Y2=0
cc_1189 N_S[3]_c_1468_n N_VPWR_c_1796_n 0.00673617f $X=20.41 $Y=1.55 $X2=0 $Y2=0
cc_1190 N_S[3]_c_1444_n VPWR 0.00846723f $X=19.94 $Y=1.55 $X2=0 $Y2=0
cc_1191 N_S[3]_c_1468_n VPWR 0.00852996f $X=20.41 $Y=1.55 $X2=0 $Y2=0
cc_1192 N_S[3]_c_1453_n N_Z_c_2200_n 0.0134253f $X=21.68 $Y=0.255 $X2=0 $Y2=0
cc_1193 N_S[3]_c_1455_n N_Z_c_2200_n 0.0077801f $X=22.1 $Y=0.255 $X2=0 $Y2=0
cc_1194 N_S[3]_c_1457_n N_Z_c_2200_n 6.35774e-19 $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_1195 N_S[3]_c_1455_n N_Z_c_2201_n 0.00190704f $X=22.1 $Y=0.255 $X2=0 $Y2=0
cc_1196 N_S[3]_c_1457_n N_Z_c_2201_n 3.10191e-19 $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_1197 N_S[3]_c_1457_n N_Z_c_2202_n 0.00283489f $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_1198 N_S[3]_c_1459_n N_Z_c_2202_n 0.002324f $X=22.94 $Y=0.255 $X2=0 $Y2=0
cc_1199 N_S[3]_c_1453_n N_Z_c_2212_n 0.00216436f $X=21.68 $Y=0.255 $X2=0 $Y2=0
cc_1200 N_S[3]_c_1457_n N_Z_c_2213_n 0.00180363f $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_1201 N_S[3]_c_1455_n N_Z_c_2214_n 6.35664e-19 $X=22.1 $Y=0.255 $X2=0 $Y2=0
cc_1202 N_S[3]_c_1457_n N_Z_c_2214_n 0.00462308f $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_1203 N_S[3]_c_1459_n N_Z_c_2214_n 0.00443615f $X=22.94 $Y=0.255 $X2=0 $Y2=0
cc_1204 N_S[3]_c_1443_n N_Z_c_2221_n 0.00234109f $X=19.84 $Y=1.16 $X2=0 $Y2=0
cc_1205 N_S[3]_c_1444_n N_Z_c_2221_n 0.0052507f $X=19.94 $Y=1.55 $X2=0 $Y2=0
cc_1206 N_S[3]_c_1468_n N_Z_c_2221_n 0.00478771f $X=20.41 $Y=1.55 $X2=0 $Y2=0
cc_1207 N_S[3]_c_1464_n N_Z_c_2221_n 0.0105931f $X=19.9 $Y=1.16 $X2=0 $Y2=0
cc_1208 N_S[3]_c_1468_n N_A_4219_311#_c_2814_n 0.00209354f $X=20.41 $Y=1.55
+ $X2=0 $Y2=0
cc_1209 N_S[3]_c_1459_n N_A_4219_311#_c_2821_n 0.00168571f $X=22.94 $Y=0.255
+ $X2=0 $Y2=0
cc_1210 N_S[3]_c_1443_n N_VGND_c_2925_n 0.00576464f $X=19.84 $Y=1.16 $X2=0 $Y2=0
cc_1211 N_S[3]_c_1445_n N_VGND_c_2925_n 0.00374526f $X=19.965 $Y=0.735 $X2=0
+ $Y2=0
cc_1212 N_S[3]_c_1464_n N_VGND_c_2925_n 0.0116218f $X=19.9 $Y=1.16 $X2=0 $Y2=0
cc_1213 N_S[3]_c_1447_n N_VGND_c_2926_n 0.00173127f $X=20.385 $Y=0.735 $X2=0
+ $Y2=0
cc_1214 N_S[3]_c_1449_n N_VGND_c_2926_n 0.00525833f $X=20.845 $Y=0.81 $X2=0
+ $Y2=0
cc_1215 N_S[3]_c_1452_n N_VGND_c_2926_n 0.00862298f $X=20.995 $Y=0.18 $X2=0
+ $Y2=0
cc_1216 N_S[3]_c_1458_n N_VGND_c_2927_n 0.0028166f $X=22.865 $Y=0.18 $X2=0 $Y2=0
cc_1217 N_S[3]_c_1459_n N_VGND_c_2927_n 5.5039e-19 $X=22.94 $Y=0.255 $X2=0 $Y2=0
cc_1218 N_S[3]_c_1445_n N_VGND_c_2947_n 0.00585385f $X=19.965 $Y=0.735 $X2=0
+ $Y2=0
cc_1219 N_S[3]_c_1446_n N_VGND_c_2947_n 2.16067e-19 $X=20.31 $Y=0.81 $X2=0 $Y2=0
cc_1220 N_S[3]_c_1447_n N_VGND_c_2947_n 0.00542362f $X=20.385 $Y=0.735 $X2=0
+ $Y2=0
cc_1221 N_S[3]_c_1452_n N_VGND_c_2949_n 0.0559651f $X=20.995 $Y=0.18 $X2=0 $Y2=0
cc_1222 N_S[3]_c_1445_n VGND 0.0119653f $X=19.965 $Y=0.735 $X2=0 $Y2=0
cc_1223 N_S[3]_c_1447_n VGND 0.00990284f $X=20.385 $Y=0.735 $X2=0 $Y2=0
cc_1224 N_S[3]_c_1451_n VGND 0.0244174f $X=21.605 $Y=0.18 $X2=0 $Y2=0
cc_1225 N_S[3]_c_1452_n VGND 0.0101627f $X=20.995 $Y=0.18 $X2=0 $Y2=0
cc_1226 N_S[3]_c_1454_n VGND 0.00642387f $X=22.025 $Y=0.18 $X2=0 $Y2=0
cc_1227 N_S[3]_c_1456_n VGND 0.0064237f $X=22.445 $Y=0.18 $X2=0 $Y2=0
cc_1228 N_S[3]_c_1458_n VGND 0.0123437f $X=22.865 $Y=0.18 $X2=0 $Y2=0
cc_1229 N_S[3]_c_1461_n VGND 0.00366655f $X=21.68 $Y=0.18 $X2=0 $Y2=0
cc_1230 N_S[3]_c_1462_n VGND 0.00366655f $X=22.1 $Y=0.18 $X2=0 $Y2=0
cc_1231 N_S[3]_c_1463_n VGND 0.00366655f $X=22.52 $Y=0.18 $X2=0 $Y2=0
cc_1232 N_S[3]_c_1450_n N_A_4269_66#_c_3496_n 0.00529837f $X=20.92 $Y=0.735
+ $X2=0 $Y2=0
cc_1233 N_S[3]_c_1453_n N_A_4269_66#_c_3497_n 0.0112916f $X=21.68 $Y=0.255 $X2=0
+ $Y2=0
cc_1234 N_S[3]_c_1454_n N_A_4269_66#_c_3497_n 0.00211351f $X=22.025 $Y=0.18
+ $X2=0 $Y2=0
cc_1235 N_S[3]_c_1455_n N_A_4269_66#_c_3497_n 0.0106844f $X=22.1 $Y=0.255 $X2=0
+ $Y2=0
cc_1236 N_S[3]_c_1450_n N_A_4269_66#_c_3498_n 0.00189496f $X=20.92 $Y=0.735
+ $X2=0 $Y2=0
cc_1237 N_S[3]_c_1451_n N_A_4269_66#_c_3498_n 0.00685838f $X=21.605 $Y=0.18
+ $X2=0 $Y2=0
cc_1238 N_S[3]_c_1457_n N_A_4269_66#_c_3499_n 0.0106826f $X=22.52 $Y=0.255 $X2=0
+ $Y2=0
cc_1239 N_S[3]_c_1458_n N_A_4269_66#_c_3499_n 0.00211351f $X=22.865 $Y=0.18
+ $X2=0 $Y2=0
cc_1240 N_S[3]_c_1459_n N_A_4269_66#_c_3499_n 0.0139014f $X=22.94 $Y=0.255 $X2=0
+ $Y2=0
cc_1241 N_S[3]_c_1459_n N_A_4269_66#_c_3502_n 0.00206084f $X=22.94 $Y=0.255
+ $X2=0 $Y2=0
cc_1242 N_S[3]_c_1456_n N_A_4269_66#_c_3515_n 0.0034777f $X=22.445 $Y=0.18 $X2=0
+ $Y2=0
cc_1243 N_A_4006_325#_c_1578_n N_VPWR_c_1778_n 0.0356181f $X=20.175 $Y=1.77
+ $X2=0 $Y2=0
cc_1244 N_A_4006_325#_c_1568_n N_VPWR_c_1779_n 0.00279288f $X=21.455 $Y=1.475
+ $X2=0 $Y2=0
cc_1245 N_A_4006_325#_c_1578_n N_VPWR_c_1779_n 0.0316788f $X=20.175 $Y=1.77
+ $X2=0 $Y2=0
cc_1246 N_A_4006_325#_c_1564_n N_VPWR_c_1779_n 0.0193185f $X=21.225 $Y=1.23
+ $X2=0 $Y2=0
cc_1247 N_A_4006_325#_c_1567_n N_VPWR_c_1779_n 6.4101e-19 $X=21.135 $Y=1.23
+ $X2=0 $Y2=0
cc_1248 N_A_4006_325#_c_1575_n N_VPWR_c_1780_n 0.00287722f $X=22.865 $Y=1.475
+ $X2=0 $Y2=0
cc_1249 N_A_4006_325#_c_1578_n N_VPWR_c_1796_n 0.0233824f $X=20.175 $Y=1.77
+ $X2=0 $Y2=0
cc_1250 N_A_4006_325#_c_1568_n N_VPWR_c_1798_n 0.00429453f $X=21.455 $Y=1.475
+ $X2=0 $Y2=0
cc_1251 N_A_4006_325#_c_1571_n N_VPWR_c_1798_n 0.00429453f $X=21.925 $Y=1.475
+ $X2=0 $Y2=0
cc_1252 N_A_4006_325#_c_1573_n N_VPWR_c_1798_n 0.00429453f $X=22.395 $Y=1.475
+ $X2=0 $Y2=0
cc_1253 N_A_4006_325#_c_1575_n N_VPWR_c_1798_n 0.00429453f $X=22.865 $Y=1.475
+ $X2=0 $Y2=0
cc_1254 N_A_4006_325#_c_1568_n VPWR 0.00737407f $X=21.455 $Y=1.475 $X2=0 $Y2=0
cc_1255 N_A_4006_325#_c_1571_n VPWR 0.0060424f $X=21.925 $Y=1.475 $X2=0 $Y2=0
cc_1256 N_A_4006_325#_c_1573_n VPWR 0.0060424f $X=22.395 $Y=1.475 $X2=0 $Y2=0
cc_1257 N_A_4006_325#_c_1575_n VPWR 0.00743756f $X=22.865 $Y=1.475 $X2=0 $Y2=0
cc_1258 N_A_4006_325#_c_1578_n VPWR 0.00593513f $X=20.175 $Y=1.77 $X2=0 $Y2=0
cc_1259 N_A_4006_325#_c_1572_n N_Z_c_2201_n 0.00762343f $X=22.305 $Y=1.4 $X2=0
+ $Y2=0
cc_1260 N_A_4006_325#_c_1577_n N_Z_c_2201_n 0.00704092f $X=22.395 $Y=1.4 $X2=0
+ $Y2=0
cc_1261 N_A_4006_325#_c_1569_n N_Z_c_2212_n 0.00597584f $X=21.835 $Y=1.4 $X2=0
+ $Y2=0
cc_1262 N_A_4006_325#_c_1561_n N_Z_c_2212_n 0.00747617f $X=21.545 $Y=1.4 $X2=0
+ $Y2=0
cc_1263 N_A_4006_325#_c_1572_n N_Z_c_2212_n 0.00145542f $X=22.305 $Y=1.4 $X2=0
+ $Y2=0
cc_1264 N_A_4006_325#_c_1576_n N_Z_c_2212_n 0.00909323f $X=21.925 $Y=1.4 $X2=0
+ $Y2=0
cc_1265 N_A_4006_325#_c_1564_n N_Z_c_2212_n 0.0266078f $X=21.225 $Y=1.23 $X2=0
+ $Y2=0
cc_1266 N_A_4006_325#_c_1574_n N_Z_c_2213_n 0.00918337f $X=22.775 $Y=1.4 $X2=0
+ $Y2=0
cc_1267 N_A_4006_325#_c_1577_n N_Z_c_2213_n 2.98555e-19 $X=22.395 $Y=1.4 $X2=0
+ $Y2=0
cc_1268 N_A_4006_325#_c_1574_n N_Z_c_2214_n 0.00248496f $X=22.775 $Y=1.4 $X2=0
+ $Y2=0
cc_1269 N_A_4006_325#_c_1568_n N_Z_c_2221_n 0.0080184f $X=21.455 $Y=1.475 $X2=0
+ $Y2=0
cc_1270 N_A_4006_325#_c_1561_n N_Z_c_2221_n 2.19754e-19 $X=21.545 $Y=1.4 $X2=0
+ $Y2=0
cc_1271 N_A_4006_325#_c_1578_n N_Z_c_2221_n 0.0329704f $X=20.175 $Y=1.77 $X2=0
+ $Y2=0
cc_1272 N_A_4006_325#_c_1564_n N_Z_c_2221_n 0.0186685f $X=21.225 $Y=1.23 $X2=0
+ $Y2=0
cc_1273 N_A_4006_325#_c_1571_n N_Z_c_2398_n 0.00378512f $X=21.925 $Y=1.475 $X2=0
+ $Y2=0
cc_1274 N_A_4006_325#_c_1573_n N_Z_c_2398_n 0.00378723f $X=22.395 $Y=1.475 $X2=0
+ $Y2=0
cc_1275 N_A_4006_325#_c_1568_n N_Z_c_2400_n 0.0107691f $X=21.455 $Y=1.475 $X2=0
+ $Y2=0
cc_1276 N_A_4006_325#_c_1569_n N_Z_c_2400_n 0.00554725f $X=21.835 $Y=1.4 $X2=0
+ $Y2=0
cc_1277 N_A_4006_325#_c_1561_n N_Z_c_2400_n 0.00415799f $X=21.545 $Y=1.4 $X2=0
+ $Y2=0
cc_1278 N_A_4006_325#_c_1571_n N_Z_c_2400_n 0.00814309f $X=21.925 $Y=1.475 $X2=0
+ $Y2=0
cc_1279 N_A_4006_325#_c_1573_n N_Z_c_2400_n 3.67612e-19 $X=22.395 $Y=1.475 $X2=0
+ $Y2=0
cc_1280 N_A_4006_325#_c_1576_n N_Z_c_2400_n 0.00313387f $X=21.925 $Y=1.4 $X2=0
+ $Y2=0
cc_1281 N_A_4006_325#_c_1564_n N_Z_c_2400_n 0.00227722f $X=21.225 $Y=1.23 $X2=0
+ $Y2=0
cc_1282 N_A_4006_325#_c_1571_n N_Z_c_2407_n 3.67612e-19 $X=21.925 $Y=1.475 $X2=0
+ $Y2=0
cc_1283 N_A_4006_325#_c_1573_n N_Z_c_2407_n 0.00814309f $X=22.395 $Y=1.475 $X2=0
+ $Y2=0
cc_1284 N_A_4006_325#_c_1574_n N_Z_c_2407_n 0.0102922f $X=22.775 $Y=1.4 $X2=0
+ $Y2=0
cc_1285 N_A_4006_325#_c_1575_n N_Z_c_2407_n 0.00899738f $X=22.865 $Y=1.475 $X2=0
+ $Y2=0
cc_1286 N_A_4006_325#_c_1577_n N_Z_c_2407_n 0.00313387f $X=22.395 $Y=1.4 $X2=0
+ $Y2=0
cc_1287 N_A_4006_325#_c_1568_n N_A_4219_311#_c_2814_n 0.00246857f $X=21.455
+ $Y=1.475 $X2=0 $Y2=0
cc_1288 N_A_4006_325#_c_1561_n N_A_4219_311#_c_2814_n 0.00561627f $X=21.545
+ $Y=1.4 $X2=0 $Y2=0
cc_1289 N_A_4006_325#_c_1564_n N_A_4219_311#_c_2814_n 0.0218124f $X=21.225
+ $Y=1.23 $X2=0 $Y2=0
cc_1290 N_A_4006_325#_c_1567_n N_A_4219_311#_c_2814_n 5.74251e-19 $X=21.135
+ $Y=1.23 $X2=0 $Y2=0
cc_1291 N_A_4006_325#_c_1568_n N_A_4219_311#_c_2815_n 0.0115457f $X=21.455
+ $Y=1.475 $X2=0 $Y2=0
cc_1292 N_A_4006_325#_c_1571_n N_A_4219_311#_c_2815_n 0.010844f $X=21.925
+ $Y=1.475 $X2=0 $Y2=0
cc_1293 N_A_4006_325#_c_1571_n N_A_4219_311#_c_2817_n 0.00102951f $X=21.925
+ $Y=1.475 $X2=0 $Y2=0
cc_1294 N_A_4006_325#_c_1572_n N_A_4219_311#_c_2817_n 0.00251792f $X=22.305
+ $Y=1.4 $X2=0 $Y2=0
cc_1295 N_A_4006_325#_c_1573_n N_A_4219_311#_c_2817_n 0.00102951f $X=22.395
+ $Y=1.475 $X2=0 $Y2=0
cc_1296 N_A_4006_325#_c_1573_n N_A_4219_311#_c_2818_n 0.010844f $X=22.395
+ $Y=1.475 $X2=0 $Y2=0
cc_1297 N_A_4006_325#_c_1575_n N_A_4219_311#_c_2818_n 0.0155783f $X=22.865
+ $Y=1.475 $X2=0 $Y2=0
cc_1298 N_A_4006_325#_c_1575_n N_A_4219_311#_c_2821_n 0.00151141f $X=22.865
+ $Y=1.475 $X2=0 $Y2=0
cc_1299 N_A_4006_325#_c_1564_n N_VGND_c_2926_n 0.0123065f $X=21.225 $Y=1.23
+ $X2=0 $Y2=0
cc_1300 N_A_4006_325#_c_1567_n N_VGND_c_2926_n 2.04129e-19 $X=21.135 $Y=1.23
+ $X2=0 $Y2=0
cc_1301 N_A_4006_325#_c_1562_n N_VGND_c_2947_n 0.0129994f $X=20.175 $Y=0.445
+ $X2=0 $Y2=0
cc_1302 N_A_4006_325#_M1059_s VGND 0.00394793f $X=20.04 $Y=0.235 $X2=0 $Y2=0
cc_1303 N_A_4006_325#_c_1562_n VGND 0.00927134f $X=20.175 $Y=0.445 $X2=0 $Y2=0
cc_1304 N_A_4006_325#_c_1561_n N_A_4269_66#_c_3496_n 0.00600378f $X=21.545
+ $Y=1.4 $X2=0 $Y2=0
cc_1305 N_A_4006_325#_c_1564_n N_A_4269_66#_c_3496_n 0.0028695f $X=21.225
+ $Y=1.23 $X2=0 $Y2=0
cc_1306 N_A_4006_325#_c_1572_n N_A_4269_66#_c_3518_n 7.0477e-19 $X=22.305 $Y=1.4
+ $X2=0 $Y2=0
cc_1307 N_D[3]_M1010_g N_VPWR_c_1780_n 0.00354866f $X=23.855 $Y=1.985 $X2=0
+ $Y2=0
cc_1308 N_D[3]_M1027_g N_VPWR_c_1781_n 0.00173895f $X=24.325 $Y=1.985 $X2=0
+ $Y2=0
cc_1309 N_D[3]_M1035_g N_VPWR_c_1781_n 0.00173895f $X=24.795 $Y=1.985 $X2=0
+ $Y2=0
cc_1310 N_D[3]_M1070_g N_VPWR_c_1783_n 0.00354866f $X=25.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1311 N_D[3]_M1010_g VPWR 0.0130007f $X=23.855 $Y=1.985 $X2=0 $Y2=0
cc_1312 N_D[3]_M1027_g VPWR 0.0117184f $X=24.325 $Y=1.985 $X2=0 $Y2=0
cc_1313 N_D[3]_M1035_g VPWR 0.0117184f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_1314 N_D[3]_M1070_g VPWR 0.0126298f $X=25.265 $Y=1.985 $X2=0 $Y2=0
cc_1315 N_D[3]_M1010_g N_VPWR_c_1805_n 0.00673617f $X=23.855 $Y=1.985 $X2=0
+ $Y2=0
cc_1316 N_D[3]_M1027_g N_VPWR_c_1805_n 0.00673617f $X=24.325 $Y=1.985 $X2=0
+ $Y2=0
cc_1317 N_D[3]_M1035_g N_VPWR_c_1806_n 0.00673617f $X=24.795 $Y=1.985 $X2=0
+ $Y2=0
cc_1318 N_D[3]_M1070_g N_VPWR_c_1806_n 0.00673617f $X=25.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1319 N_D[3]_M1010_g N_A_4219_311#_c_2819_n 0.00330737f $X=23.855 $Y=1.985
+ $X2=0 $Y2=0
cc_1320 N_D[3]_M1010_g N_A_4219_311#_c_2820_n 0.017872f $X=23.855 $Y=1.985 $X2=0
+ $Y2=0
cc_1321 N_D[3]_M1010_g N_A_4219_311#_c_2839_n 0.010906f $X=23.855 $Y=1.985 $X2=0
+ $Y2=0
cc_1322 N_D[3]_M1027_g N_A_4219_311#_c_2839_n 0.0100233f $X=24.325 $Y=1.985
+ $X2=0 $Y2=0
cc_1323 N_D[3]_M1035_g N_A_4219_311#_c_2839_n 5.91934e-19 $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_1324 N_D[3]_M1027_g N_A_4219_311#_c_2842_n 0.0137916f $X=24.325 $Y=1.985
+ $X2=0 $Y2=0
cc_1325 N_D[3]_M1035_g N_A_4219_311#_c_2842_n 0.0137916f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_1326 N_D[3]_c_1683_n N_A_4219_311#_c_2842_n 7.15862e-19 $X=24.705 $Y=1.16
+ $X2=0 $Y2=0
cc_1327 N_D[3]_c_1685_n N_A_4219_311#_c_2842_n 0.0405252f $X=25.16 $Y=1.16 $X2=0
+ $Y2=0
cc_1328 N_D[3]_M1035_g N_A_4219_311#_c_2846_n 5.79575e-19 $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_1329 N_D[3]_M1070_g N_A_4219_311#_c_2846_n 0.00215964f $X=25.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1330 N_D[3]_c_1685_n N_A_4219_311#_c_2846_n 0.022724f $X=25.16 $Y=1.16 $X2=0
+ $Y2=0
cc_1331 N_D[3]_c_1686_n N_A_4219_311#_c_2846_n 8.03631e-19 $X=25.265 $Y=1.16
+ $X2=0 $Y2=0
cc_1332 N_D[3]_M1027_g N_A_4219_311#_c_2850_n 5.91934e-19 $X=24.325 $Y=1.985
+ $X2=0 $Y2=0
cc_1333 N_D[3]_M1035_g N_A_4219_311#_c_2850_n 0.0100233f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_1334 N_D[3]_M1070_g N_A_4219_311#_c_2850_n 0.00897418f $X=25.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1335 N_D[3]_M1010_g N_A_4219_311#_c_2853_n 8.61029e-19 $X=23.855 $Y=1.985
+ $X2=0 $Y2=0
cc_1336 N_D[3]_M1027_g N_A_4219_311#_c_2853_n 5.79575e-19 $X=24.325 $Y=1.985
+ $X2=0 $Y2=0
cc_1337 N_D[3]_c_1684_n N_A_4219_311#_c_2853_n 8.03631e-19 $X=24.415 $Y=1.16
+ $X2=0 $Y2=0
cc_1338 N_D[3]_c_1685_n N_A_4219_311#_c_2853_n 0.0199757f $X=25.16 $Y=1.16 $X2=0
+ $Y2=0
cc_1339 N_D[3]_M1013_g N_VGND_c_2927_n 0.00321269f $X=23.88 $Y=0.56 $X2=0 $Y2=0
cc_1340 N_D[3]_M1032_g N_VGND_c_2927_n 2.6376e-19 $X=24.3 $Y=0.56 $X2=0 $Y2=0
cc_1341 N_D[3]_M1032_g N_VGND_c_2928_n 0.0019152f $X=24.3 $Y=0.56 $X2=0 $Y2=0
cc_1342 N_D[3]_M1040_g N_VGND_c_2928_n 0.00166854f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_1343 N_D[3]_M1054_g N_VGND_c_2928_n 2.64031e-19 $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_1344 N_D[3]_M1054_g N_VGND_c_2930_n 0.00345859f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_1345 N_D[3]_M1013_g VGND 0.00702263f $X=23.88 $Y=0.56 $X2=0 $Y2=0
cc_1346 N_D[3]_M1032_g VGND 0.00624811f $X=24.3 $Y=0.56 $X2=0 $Y2=0
cc_1347 N_D[3]_M1040_g VGND 0.00593887f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_1348 N_D[3]_M1054_g VGND 0.0107845f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_1349 N_D[3]_M1013_g N_VGND_c_2956_n 0.00422241f $X=23.88 $Y=0.56 $X2=0 $Y2=0
cc_1350 N_D[3]_M1032_g N_VGND_c_2956_n 0.00430643f $X=24.3 $Y=0.56 $X2=0 $Y2=0
cc_1351 N_D[3]_M1040_g N_VGND_c_2957_n 0.00422241f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_1352 N_D[3]_M1054_g N_VGND_c_2957_n 0.00551064f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_1353 N_D[3]_M1013_g N_A_4269_66#_c_3500_n 0.00261078f $X=23.88 $Y=0.56 $X2=0
+ $Y2=0
cc_1354 N_D[3]_M1013_g N_A_4269_66#_c_3501_n 0.0121912f $X=23.88 $Y=0.56 $X2=0
+ $Y2=0
cc_1355 N_D[3]_M1013_g N_A_4269_66#_c_3521_n 0.00699463f $X=23.88 $Y=0.56 $X2=0
+ $Y2=0
cc_1356 N_D[3]_M1032_g N_A_4269_66#_c_3521_n 0.00661764f $X=24.3 $Y=0.56 $X2=0
+ $Y2=0
cc_1357 N_D[3]_M1040_g N_A_4269_66#_c_3521_n 5.22365e-19 $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_1358 N_D[3]_M1032_g N_A_4269_66#_c_3503_n 0.00900364f $X=24.3 $Y=0.56 $X2=0
+ $Y2=0
cc_1359 N_D[3]_M1040_g N_A_4269_66#_c_3503_n 0.00986515f $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_1360 N_D[3]_M1054_g N_A_4269_66#_c_3503_n 0.00228093f $X=25.24 $Y=0.56 $X2=0
+ $Y2=0
cc_1361 N_D[3]_c_1683_n N_A_4269_66#_c_3503_n 0.00463549f $X=24.705 $Y=1.16
+ $X2=0 $Y2=0
cc_1362 N_D[3]_c_1685_n N_A_4269_66#_c_3503_n 0.0608884f $X=25.16 $Y=1.16 $X2=0
+ $Y2=0
cc_1363 N_D[3]_c_1686_n N_A_4269_66#_c_3503_n 0.00208088f $X=25.265 $Y=1.16
+ $X2=0 $Y2=0
cc_1364 N_D[3]_M1032_g N_A_4269_66#_c_3530_n 5.22365e-19 $X=24.3 $Y=0.56 $X2=0
+ $Y2=0
cc_1365 N_D[3]_M1040_g N_A_4269_66#_c_3530_n 0.00661134f $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_1366 N_D[3]_M1054_g N_A_4269_66#_c_3530_n 0.00529286f $X=25.24 $Y=0.56 $X2=0
+ $Y2=0
cc_1367 N_D[3]_M1013_g N_A_4269_66#_c_3504_n 0.00128201f $X=23.88 $Y=0.56 $X2=0
+ $Y2=0
cc_1368 N_D[3]_M1032_g N_A_4269_66#_c_3504_n 8.68782e-19 $X=24.3 $Y=0.56 $X2=0
+ $Y2=0
cc_1369 N_D[3]_c_1684_n N_A_4269_66#_c_3504_n 0.00208088f $X=24.415 $Y=1.16
+ $X2=0 $Y2=0
cc_1370 N_D[3]_c_1685_n N_A_4269_66#_c_3504_n 0.018367f $X=25.16 $Y=1.16 $X2=0
+ $Y2=0
cc_1371 VPWR N_A_117_297#_M1003_s 0.00231261f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_1372 VPWR N_A_117_297#_M1055_s 0.00231261f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1373 VPWR N_A_117_297#_c_2114_n 0.0123132f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1374 N_VPWR_c_1801_n N_A_117_297#_c_2114_n 0.0189467f $X=1.065 $Y=2.72 $X2=0
+ $Y2=0
cc_1375 N_VPWR_M1041_d N_A_117_297#_c_2117_n 0.00350459f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_1376 N_VPWR_c_1759_n N_A_117_297#_c_2117_n 0.0143191f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_1377 N_VPWR_c_1760_n N_A_117_297#_c_2121_n 0.0189467f $X=2.005 $Y=2.72 $X2=0
+ $Y2=0
cc_1378 VPWR N_A_117_297#_c_2121_n 0.0123132f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1379 N_VPWR_M1071_d N_A_117_297#_c_2102_n 0.00737891f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_1380 N_VPWR_c_1761_n N_A_117_297#_c_2102_n 0.0180895f $X=2.14 $Y=2 $X2=0
+ $Y2=0
cc_1381 N_VPWR_c_1761_n N_A_117_297#_c_2103_n 0.03124f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_1382 N_VPWR_c_1784_n N_A_117_297#_c_2104_n 0.0420587f $X=4.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1383 VPWR N_A_117_297#_c_2104_n 0.0138198f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1384 N_VPWR_c_1761_n N_A_117_297#_c_2105_n 0.0123662f $X=2.14 $Y=2 $X2=0
+ $Y2=0
cc_1385 N_VPWR_c_1784_n N_A_117_297#_c_2105_n 0.0215086f $X=4.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1386 VPWR N_A_117_297#_c_2105_n 0.0115535f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1387 N_VPWR_c_1762_n N_A_117_297#_c_2107_n 0.0114906f $X=5.115 $Y=1.77 $X2=0
+ $Y2=0
cc_1388 N_VPWR_c_1784_n N_A_117_297#_c_2107_n 0.0635672f $X=4.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1389 VPWR N_A_117_297#_c_2107_n 0.0159283f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1390 N_VPWR_c_1762_n N_A_117_297#_c_2108_n 0.0417486f $X=5.115 $Y=1.77 $X2=0
+ $Y2=0
cc_1391 N_VPWR_c_1784_n N_A_117_297#_c_2109_n 0.0193577f $X=4.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1392 VPWR N_A_117_297#_c_2109_n 0.00495316f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1393 N_VPWR_M1004_d N_Z_c_2219_n 8.15553e-19 $X=4.99 $Y=1.625 $X2=0 $Y2=0
cc_1394 N_VPWR_M1018_d N_Z_c_2219_n 2.0504e-19 $X=5.91 $Y=1.625 $X2=0 $Y2=0
cc_1395 N_VPWR_M1036_d N_Z_c_2219_n 2.0504e-19 $X=6.7 $Y=1.625 $X2=0 $Y2=0
cc_1396 N_VPWR_M1050_d N_Z_c_2219_n 8.15553e-19 $X=7.62 $Y=1.625 $X2=0 $Y2=0
cc_1397 N_VPWR_c_1762_n N_Z_c_2219_n 0.0196216f $X=5.115 $Y=1.77 $X2=0 $Y2=0
cc_1398 N_VPWR_c_1763_n N_Z_c_2219_n 0.0222682f $X=6.055 $Y=1.77 $X2=0 $Y2=0
cc_1399 N_VPWR_c_1765_n N_Z_c_2219_n 0.0222682f $X=6.825 $Y=1.77 $X2=0 $Y2=0
cc_1400 N_VPWR_c_1766_n N_Z_c_2219_n 0.0196216f $X=7.765 $Y=1.77 $X2=0 $Y2=0
cc_1401 VPWR N_Z_c_2219_n 0.209432f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1402 VPWR N_Z_c_2421_n 0.0146963f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1403 N_VPWR_M1001_s N_Z_c_2220_n 0.00217353f $X=10.615 $Y=1.485 $X2=0 $Y2=0
cc_1404 N_VPWR_M1006_s N_Z_c_2220_n 0.00243967f $X=11.535 $Y=1.485 $X2=0 $Y2=0
cc_1405 N_VPWR_M1065_s N_Z_c_2220_n 2.0504e-19 $X=12.475 $Y=1.485 $X2=0 $Y2=0
cc_1406 N_VPWR_M1005_s N_Z_c_2220_n 2.0504e-19 $X=13.015 $Y=1.485 $X2=0 $Y2=0
cc_1407 N_VPWR_M1019_s N_Z_c_2220_n 0.00243967f $X=13.935 $Y=1.485 $X2=0 $Y2=0
cc_1408 N_VPWR_M1074_s N_Z_c_2220_n 0.00217353f $X=14.875 $Y=1.485 $X2=0 $Y2=0
cc_1409 N_VPWR_c_1767_n N_Z_c_2220_n 0.0138089f $X=10.74 $Y=2 $X2=0 $Y2=0
cc_1410 N_VPWR_c_1768_n N_Z_c_2220_n 0.0135506f $X=11.68 $Y=2 $X2=0 $Y2=0
cc_1411 N_VPWR_c_1769_n N_Z_c_2220_n 0.0276847f $X=12.62 $Y=1.66 $X2=0 $Y2=0
cc_1412 N_VPWR_c_1771_n N_Z_c_2220_n 0.0276847f $X=13.14 $Y=1.66 $X2=0 $Y2=0
cc_1413 N_VPWR_c_1772_n N_Z_c_2220_n 0.0135506f $X=14.08 $Y=2 $X2=0 $Y2=0
cc_1414 N_VPWR_c_1774_n N_Z_c_2220_n 0.0138089f $X=15.02 $Y=2 $X2=0 $Y2=0
cc_1415 VPWR N_Z_c_2220_n 0.275096f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1416 VPWR N_Z_c_2435_n 0.0146963f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1417 N_VPWR_M1020_s N_Z_c_2221_n 8.15553e-19 $X=17.87 $Y=1.625 $X2=0 $Y2=0
cc_1418 N_VPWR_M1076_s N_Z_c_2221_n 2.0504e-19 $X=18.79 $Y=1.625 $X2=0 $Y2=0
cc_1419 N_VPWR_M1045_s N_Z_c_2221_n 2.0504e-19 $X=19.58 $Y=1.625 $X2=0 $Y2=0
cc_1420 N_VPWR_M1067_s N_Z_c_2221_n 8.15553e-19 $X=20.5 $Y=1.625 $X2=0 $Y2=0
cc_1421 N_VPWR_c_1775_n N_Z_c_2221_n 0.0196216f $X=17.995 $Y=1.77 $X2=0 $Y2=0
cc_1422 N_VPWR_c_1776_n N_Z_c_2221_n 0.0222682f $X=18.935 $Y=1.77 $X2=0 $Y2=0
cc_1423 N_VPWR_c_1778_n N_Z_c_2221_n 0.0222682f $X=19.705 $Y=1.77 $X2=0 $Y2=0
cc_1424 N_VPWR_c_1779_n N_Z_c_2221_n 0.0196216f $X=20.645 $Y=1.77 $X2=0 $Y2=0
cc_1425 VPWR N_Z_c_2221_n 0.209432f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1426 VPWR N_Z_c_2445_n 0.0146963f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1427 VPWR N_Z_c_2298_n 0.0307257f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1428 VPWR N_Z_c_2447_n 0.0146963f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1429 VPWR N_Z_c_2398_n 0.0307257f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1430 VPWR N_Z_c_2449_n 0.0146963f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1431 VPWR Z 0.0307257f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1432 VPWR Z 0.0146963f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1433 VPWR Z 0.0307257f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1434 VPWR Z 0.0146963f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1435 VPWR N_Z_c_2454_n 0.0146963f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1436 VPWR N_A_1643_311#_M1001_d 0.00190235f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1437 VPWR N_A_1643_311#_M1038_d 0.00190235f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1438 N_VPWR_c_1766_n N_A_1643_311#_c_2607_n 0.0417486f $X=7.765 $Y=1.77 $X2=0
+ $Y2=0
cc_1439 N_VPWR_c_1790_n N_A_1643_311#_c_2608_n 0.0420587f $X=10.605 $Y=2.72
+ $X2=0 $Y2=0
cc_1440 VPWR N_A_1643_311#_c_2608_n 0.0104248f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1441 N_VPWR_c_1766_n N_A_1643_311#_c_2609_n 0.0114906f $X=7.765 $Y=1.77 $X2=0
+ $Y2=0
cc_1442 N_VPWR_c_1790_n N_A_1643_311#_c_2609_n 0.0215086f $X=10.605 $Y=2.72
+ $X2=0 $Y2=0
cc_1443 VPWR N_A_1643_311#_c_2609_n 0.00550351f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1444 N_VPWR_c_1767_n N_A_1643_311#_c_2611_n 0.0123662f $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_1445 N_VPWR_c_1790_n N_A_1643_311#_c_2611_n 0.0635672f $X=10.605 $Y=2.72
+ $X2=0 $Y2=0
cc_1446 VPWR N_A_1643_311#_c_2611_n 0.0159283f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1447 N_VPWR_c_1767_n N_A_1643_311#_c_2612_n 0.0299454f $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_1448 N_VPWR_M1001_s N_A_1643_311#_c_2613_n 0.00715085f $X=10.615 $Y=1.485
+ $X2=0 $Y2=0
cc_1449 N_VPWR_c_1767_n N_A_1643_311#_c_2613_n 0.0152464f $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_1450 N_VPWR_c_1767_n N_A_1643_311#_c_2633_n 0.0250039f $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_1451 N_VPWR_c_1768_n N_A_1643_311#_c_2633_n 0.0250039f $X=11.68 $Y=2 $X2=0
+ $Y2=0
cc_1452 VPWR N_A_1643_311#_c_2633_n 0.00586606f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1453 N_VPWR_c_1802_n N_A_1643_311#_c_2633_n 0.0189467f $X=11.545 $Y=2.72
+ $X2=0 $Y2=0
cc_1454 N_VPWR_M1006_s N_A_1643_311#_c_2636_n 0.00331615f $X=11.535 $Y=1.485
+ $X2=0 $Y2=0
cc_1455 N_VPWR_c_1768_n N_A_1643_311#_c_2636_n 0.0130979f $X=11.68 $Y=2 $X2=0
+ $Y2=0
cc_1456 N_VPWR_c_1768_n N_A_1643_311#_c_2644_n 0.0250039f $X=11.68 $Y=2 $X2=0
+ $Y2=0
cc_1457 N_VPWR_c_1769_n N_A_1643_311#_c_2644_n 0.0318001f $X=12.62 $Y=1.66 $X2=0
+ $Y2=0
cc_1458 VPWR N_A_1643_311#_c_2644_n 0.00586606f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1459 N_VPWR_c_1803_n N_A_1643_311#_c_2644_n 0.0189467f $X=12.485 $Y=2.72
+ $X2=0 $Y2=0
cc_1460 N_VPWR_c_1790_n N_A_1643_311#_c_2615_n 0.0193577f $X=10.605 $Y=2.72
+ $X2=0 $Y2=0
cc_1461 VPWR N_A_1643_311#_c_2615_n 0.00495316f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1462 VPWR N_A_2693_297#_M1005_d 0.00190235f $X=25.445 $Y=2.635 $X2=-0.19
+ $Y2=-0.24
cc_1463 VPWR N_A_2693_297#_M1047_d 0.00190235f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1464 N_VPWR_c_1771_n N_A_2693_297#_c_2724_n 0.0318001f $X=13.14 $Y=1.66 $X2=0
+ $Y2=0
cc_1465 N_VPWR_c_1772_n N_A_2693_297#_c_2724_n 0.0250039f $X=14.08 $Y=2 $X2=0
+ $Y2=0
cc_1466 VPWR N_A_2693_297#_c_2724_n 0.00586606f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1467 N_VPWR_c_1804_n N_A_2693_297#_c_2724_n 0.0189467f $X=13.945 $Y=2.72
+ $X2=0 $Y2=0
cc_1468 N_VPWR_M1019_s N_A_2693_297#_c_2727_n 0.00331615f $X=13.935 $Y=1.485
+ $X2=0 $Y2=0
cc_1469 N_VPWR_c_1772_n N_A_2693_297#_c_2727_n 0.0130979f $X=14.08 $Y=2 $X2=0
+ $Y2=0
cc_1470 N_VPWR_c_1772_n N_A_2693_297#_c_2731_n 0.0250039f $X=14.08 $Y=2 $X2=0
+ $Y2=0
cc_1471 N_VPWR_c_1773_n N_A_2693_297#_c_2731_n 0.0189467f $X=14.885 $Y=2.72
+ $X2=0 $Y2=0
cc_1472 N_VPWR_c_1774_n N_A_2693_297#_c_2731_n 0.0250039f $X=15.02 $Y=2 $X2=0
+ $Y2=0
cc_1473 VPWR N_A_2693_297#_c_2731_n 0.00586606f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1474 N_VPWR_M1074_s N_A_2693_297#_c_2712_n 0.00715085f $X=14.875 $Y=1.485
+ $X2=0 $Y2=0
cc_1475 N_VPWR_c_1774_n N_A_2693_297#_c_2712_n 0.0152464f $X=15.02 $Y=2 $X2=0
+ $Y2=0
cc_1476 N_VPWR_c_1774_n N_A_2693_297#_c_2713_n 0.0299454f $X=15.02 $Y=2 $X2=0
+ $Y2=0
cc_1477 N_VPWR_c_1792_n N_A_2693_297#_c_2714_n 0.0420587f $X=17.83 $Y=2.72 $X2=0
+ $Y2=0
cc_1478 VPWR N_A_2693_297#_c_2714_n 0.0104248f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1479 N_VPWR_c_1774_n N_A_2693_297#_c_2715_n 0.0123662f $X=15.02 $Y=2 $X2=0
+ $Y2=0
cc_1480 N_VPWR_c_1792_n N_A_2693_297#_c_2715_n 0.0215086f $X=17.83 $Y=2.72 $X2=0
+ $Y2=0
cc_1481 VPWR N_A_2693_297#_c_2715_n 0.00550351f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1482 N_VPWR_c_1775_n N_A_2693_297#_c_2717_n 0.0114906f $X=17.995 $Y=1.77
+ $X2=0 $Y2=0
cc_1483 N_VPWR_c_1792_n N_A_2693_297#_c_2717_n 0.0635672f $X=17.83 $Y=2.72 $X2=0
+ $Y2=0
cc_1484 VPWR N_A_2693_297#_c_2717_n 0.0159283f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1485 N_VPWR_c_1775_n N_A_2693_297#_c_2718_n 0.0417486f $X=17.995 $Y=1.77
+ $X2=0 $Y2=0
cc_1486 N_VPWR_c_1792_n N_A_2693_297#_c_2719_n 0.0193577f $X=17.83 $Y=2.72 $X2=0
+ $Y2=0
cc_1487 VPWR N_A_2693_297#_c_2719_n 0.00495316f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1488 VPWR N_A_4219_311#_M1010_s 0.00231261f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1489 VPWR N_A_4219_311#_M1035_s 0.00231261f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1490 N_VPWR_c_1779_n N_A_4219_311#_c_2814_n 0.0417486f $X=20.645 $Y=1.77
+ $X2=0 $Y2=0
cc_1491 N_VPWR_c_1798_n N_A_4219_311#_c_2815_n 0.0420587f $X=23.485 $Y=2.72
+ $X2=0 $Y2=0
cc_1492 VPWR N_A_4219_311#_c_2815_n 0.0104248f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1493 N_VPWR_c_1779_n N_A_4219_311#_c_2816_n 0.0114906f $X=20.645 $Y=1.77
+ $X2=0 $Y2=0
cc_1494 N_VPWR_c_1798_n N_A_4219_311#_c_2816_n 0.0215086f $X=23.485 $Y=2.72
+ $X2=0 $Y2=0
cc_1495 VPWR N_A_4219_311#_c_2816_n 0.00550351f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1496 N_VPWR_c_1780_n N_A_4219_311#_c_2818_n 0.0123662f $X=23.62 $Y=2 $X2=0
+ $Y2=0
cc_1497 N_VPWR_c_1798_n N_A_4219_311#_c_2818_n 0.0635672f $X=23.485 $Y=2.72
+ $X2=0 $Y2=0
cc_1498 VPWR N_A_4219_311#_c_2818_n 0.0253734f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1499 N_VPWR_c_1780_n N_A_4219_311#_c_2819_n 0.03124f $X=23.62 $Y=2 $X2=0
+ $Y2=0
cc_1500 N_VPWR_M1010_d N_A_4219_311#_c_2820_n 0.00737891f $X=23.495 $Y=1.485
+ $X2=0 $Y2=0
cc_1501 N_VPWR_c_1780_n N_A_4219_311#_c_2820_n 0.0180895f $X=23.62 $Y=2 $X2=0
+ $Y2=0
cc_1502 VPWR N_A_4219_311#_c_2839_n 0.0123132f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1503 N_VPWR_c_1805_n N_A_4219_311#_c_2839_n 0.0189467f $X=24.425 $Y=2.72
+ $X2=0 $Y2=0
cc_1504 N_VPWR_M1027_d N_A_4219_311#_c_2842_n 0.00350459f $X=24.415 $Y=1.485
+ $X2=0 $Y2=0
cc_1505 N_VPWR_c_1781_n N_A_4219_311#_c_2842_n 0.0143191f $X=24.56 $Y=2 $X2=0
+ $Y2=0
cc_1506 VPWR N_A_4219_311#_c_2850_n 0.0123132f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1507 N_VPWR_c_1806_n N_A_4219_311#_c_2850_n 0.0189467f $X=25.365 $Y=2.72
+ $X2=0 $Y2=0
cc_1508 N_VPWR_c_1798_n N_A_4219_311#_c_2822_n 0.0193577f $X=23.485 $Y=2.72
+ $X2=0 $Y2=0
cc_1509 VPWR N_A_4219_311#_c_2822_n 0.00495316f $X=25.445 $Y=2.635 $X2=0 $Y2=0
cc_1510 N_VPWR_c_1758_n N_VGND_c_2907_n 0.00764703f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_1511 N_VPWR_c_1769_n N_VGND_c_2917_n 0.00764703f $X=12.62 $Y=1.66 $X2=0 $Y2=0
cc_1512 N_VPWR_c_1771_n N_VGND_c_2919_n 0.00764703f $X=13.14 $Y=1.66 $X2=0 $Y2=0
cc_1513 N_VPWR_c_1783_n N_VGND_c_2930_n 0.00764703f $X=25.5 $Y=1.66 $X2=0 $Y2=0
cc_1514 N_A_117_297#_c_2104_n N_Z_M1042_s 0.00176676f $X=3.465 $Y=2.38 $X2=0
+ $Y2=0
cc_1515 N_A_117_297#_c_2107_n N_Z_M1063_s 0.00176676f $X=4.405 $Y=2.38 $X2=0
+ $Y2=0
cc_1516 N_A_117_297#_c_2106_n N_Z_c_2192_n 0.0192125f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_1517 N_A_117_297#_c_2106_n N_Z_c_2205_n 0.0024794f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_1518 N_A_117_297#_M1072_d N_Z_c_2219_n 2.07056e-19 $X=4.395 $Y=1.555 $X2=0
+ $Y2=0
cc_1519 N_A_117_297#_c_2107_n N_Z_c_2219_n 0.00349489f $X=4.405 $Y=2.38 $X2=0
+ $Y2=0
cc_1520 N_A_117_297#_c_2108_n N_Z_c_2219_n 0.0209902f $X=4.54 $Y=1.73 $X2=0
+ $Y2=0
cc_1521 N_A_117_297#_c_2106_n N_Z_c_2421_n 6.68271e-19 $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_1522 N_A_117_297#_c_2107_n N_Z_c_2421_n 9.16304e-19 $X=4.405 $Y=2.38 $X2=0
+ $Y2=0
cc_1523 N_A_117_297#_c_2108_n N_Z_c_2421_n 6.74054e-19 $X=4.54 $Y=1.73 $X2=0
+ $Y2=0
cc_1524 N_A_117_297#_M1056_d Z 3.24931e-19 $X=3.455 $Y=1.555 $X2=0 $Y2=0
cc_1525 N_A_117_297#_c_2104_n Z 0.00349489f $X=3.465 $Y=2.38 $X2=0 $Y2=0
cc_1526 N_A_117_297#_c_2106_n Z 0.0189041f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_1527 N_A_117_297#_c_2107_n Z 0.00349489f $X=4.405 $Y=2.38 $X2=0 $Y2=0
cc_1528 N_A_117_297#_c_2102_n N_Z_c_2239_n 0.00915958f $X=2.495 $Y=1.58 $X2=0
+ $Y2=0
cc_1529 N_A_117_297#_c_2104_n N_Z_c_2239_n 0.0151266f $X=3.465 $Y=2.38 $X2=0
+ $Y2=0
cc_1530 N_A_117_297#_c_2106_n N_Z_c_2239_n 0.0247248f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_1531 N_A_117_297#_c_2106_n N_Z_c_2245_n 0.0247248f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_1532 N_A_117_297#_c_2107_n N_Z_c_2245_n 0.0150524f $X=4.405 $Y=2.38 $X2=0
+ $Y2=0
cc_1533 N_A_117_297#_c_2108_n N_Z_c_2245_n 0.0228406f $X=4.54 $Y=1.73 $X2=0
+ $Y2=0
cc_1534 N_A_117_297#_c_2103_n N_Z_c_2454_n 0.00168706f $X=2.66 $Y=1.7 $X2=0
+ $Y2=0
cc_1535 N_A_117_297#_c_2104_n N_Z_c_2454_n 9.16304e-19 $X=3.465 $Y=2.38 $X2=0
+ $Y2=0
cc_1536 N_A_117_297#_c_2106_n N_Z_c_2454_n 6.68271e-19 $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_1537 N_A_117_297#_c_2102_n N_A_119_47#_c_3247_n 0.0247972f $X=2.495 $Y=1.58
+ $X2=0 $Y2=0
cc_1538 N_A_117_297#_c_2126_n N_A_119_47#_c_3253_n 6.95815e-19 $X=1.67 $Y=1.66
+ $X2=0 $Y2=0
cc_1539 N_Z_c_2219_n N_A_1643_311#_M1000_s 2.07056e-19 $X=8.665 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_1540 N_Z_c_2298_n N_A_1643_311#_M1014_s 3.24931e-19 $X=9.605 $Y=1.87 $X2=0
+ $Y2=0
cc_1541 N_Z_c_2220_n N_A_1643_311#_M1066_s 2.07056e-19 $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1542 N_Z_c_2219_n N_A_1643_311#_c_2607_n 0.0209902f $X=8.665 $Y=1.87 $X2=0
+ $Y2=0
cc_1543 Z N_A_1643_311#_c_2607_n 6.74054e-19 $X=8.785 $Y=1.785 $X2=0 $Y2=0
cc_1544 N_Z_c_2300_n N_A_1643_311#_c_2607_n 0.0228406f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_1545 N_Z_M1000_d N_A_1643_311#_c_2608_n 0.00176676f $X=8.665 $Y=1.555 $X2=0
+ $Y2=0
cc_1546 N_Z_c_2219_n N_A_1643_311#_c_2608_n 0.00349489f $X=8.665 $Y=1.87 $X2=0
+ $Y2=0
cc_1547 N_Z_c_2298_n N_A_1643_311#_c_2608_n 0.00349489f $X=9.605 $Y=1.87 $X2=0
+ $Y2=0
cc_1548 Z N_A_1643_311#_c_2608_n 9.16304e-19 $X=8.785 $Y=1.785 $X2=0 $Y2=0
cc_1549 N_Z_c_2300_n N_A_1643_311#_c_2608_n 0.0150524f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_1550 N_Z_c_2195_n N_A_1643_311#_c_2610_n 0.0192125f $X=9.585 $Y=1.215 $X2=0
+ $Y2=0
cc_1551 N_Z_c_2206_n N_A_1643_311#_c_2610_n 0.0024794f $X=8.91 $Y=1.215 $X2=0
+ $Y2=0
cc_1552 N_Z_c_2435_n N_A_1643_311#_c_2610_n 6.68271e-19 $X=9.895 $Y=1.87 $X2=0
+ $Y2=0
cc_1553 N_Z_c_2298_n N_A_1643_311#_c_2610_n 0.0189041f $X=9.605 $Y=1.87 $X2=0
+ $Y2=0
cc_1554 Z N_A_1643_311#_c_2610_n 6.68271e-19 $X=8.785 $Y=1.785 $X2=0 $Y2=0
cc_1555 N_Z_c_2300_n N_A_1643_311#_c_2610_n 0.0247248f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_1556 N_Z_c_2307_n N_A_1643_311#_c_2610_n 0.0247248f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_1557 N_Z_M1043_d N_A_1643_311#_c_2611_n 0.00176676f $X=9.605 $Y=1.555 $X2=0
+ $Y2=0
cc_1558 N_Z_c_2220_n N_A_1643_311#_c_2611_n 0.00349489f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1559 N_Z_c_2435_n N_A_1643_311#_c_2611_n 9.16304e-19 $X=9.895 $Y=1.87 $X2=0
+ $Y2=0
cc_1560 N_Z_c_2298_n N_A_1643_311#_c_2611_n 0.00349489f $X=9.605 $Y=1.87 $X2=0
+ $Y2=0
cc_1561 N_Z_c_2307_n N_A_1643_311#_c_2611_n 0.0150524f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_1562 N_Z_c_2220_n N_A_1643_311#_c_2612_n 0.0307463f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1563 N_Z_c_2435_n N_A_1643_311#_c_2612_n 6.74054e-19 $X=9.895 $Y=1.87 $X2=0
+ $Y2=0
cc_1564 N_Z_c_2307_n N_A_1643_311#_c_2612_n 0.0190884f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_1565 N_Z_c_2220_n N_A_1643_311#_c_2613_n 0.0242319f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1566 N_Z_c_2307_n N_A_1643_311#_c_2614_n 0.00915958f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_1567 N_Z_c_2220_n N_A_1643_311#_c_2633_n 0.0250077f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1568 N_Z_c_2220_n N_A_1643_311#_c_2636_n 0.020688f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1569 N_Z_c_2220_n N_A_1643_311#_c_2644_n 0.0230384f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1570 N_Z_c_2220_n N_A_2693_297#_M1025_d 2.07056e-19 $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1571 Z N_A_2693_297#_M1044_d 3.24931e-19 $X=16.805 $Y=1.785 $X2=0 $Y2=0
cc_1572 N_Z_c_2221_n N_A_2693_297#_M1064_d 2.07056e-19 $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_1573 N_Z_c_2220_n N_A_2693_297#_c_2724_n 0.0230384f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1574 N_Z_c_2220_n N_A_2693_297#_c_2727_n 0.020688f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1575 N_Z_c_2220_n N_A_2693_297#_c_2731_n 0.0250077f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1576 N_Z_c_2220_n N_A_2693_297#_c_2712_n 0.0242319f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1577 N_Z_c_2340_n N_A_2693_297#_c_2712_n 0.00915958f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_1578 N_Z_c_2220_n N_A_2693_297#_c_2713_n 0.0307463f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1579 N_Z_c_2447_n N_A_2693_297#_c_2713_n 6.74054e-19 $X=16.155 $Y=1.87 $X2=0
+ $Y2=0
cc_1580 N_Z_c_2340_n N_A_2693_297#_c_2713_n 0.0190884f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_1581 N_Z_M1025_s N_A_2693_297#_c_2714_n 0.00176676f $X=15.865 $Y=1.555 $X2=0
+ $Y2=0
cc_1582 N_Z_c_2220_n N_A_2693_297#_c_2714_n 0.00349489f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_1583 N_Z_c_2447_n N_A_2693_297#_c_2714_n 9.16304e-19 $X=16.155 $Y=1.87 $X2=0
+ $Y2=0
cc_1584 Z N_A_2693_297#_c_2714_n 0.00349489f $X=16.805 $Y=1.785 $X2=0 $Y2=0
cc_1585 N_Z_c_2340_n N_A_2693_297#_c_2714_n 0.0150524f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_1586 N_Z_c_2198_n N_A_2693_297#_c_2716_n 0.0192125f $X=16.585 $Y=1.215 $X2=0
+ $Y2=0
cc_1587 N_Z_c_2211_n N_A_2693_297#_c_2716_n 0.0024794f $X=16.85 $Y=1.215 $X2=0
+ $Y2=0
cc_1588 N_Z_c_2445_n N_A_2693_297#_c_2716_n 6.68271e-19 $X=17.095 $Y=1.87 $X2=0
+ $Y2=0
cc_1589 N_Z_c_2447_n N_A_2693_297#_c_2716_n 6.68271e-19 $X=16.155 $Y=1.87 $X2=0
+ $Y2=0
cc_1590 Z N_A_2693_297#_c_2716_n 0.0189041f $X=16.805 $Y=1.785 $X2=0 $Y2=0
cc_1591 N_Z_c_2340_n N_A_2693_297#_c_2716_n 0.0247248f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_1592 N_Z_c_2346_n N_A_2693_297#_c_2716_n 0.0247248f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_1593 N_Z_M1051_s N_A_2693_297#_c_2717_n 0.00176676f $X=16.805 $Y=1.555 $X2=0
+ $Y2=0
cc_1594 N_Z_c_2221_n N_A_2693_297#_c_2717_n 0.00349489f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_1595 N_Z_c_2445_n N_A_2693_297#_c_2717_n 9.16304e-19 $X=17.095 $Y=1.87 $X2=0
+ $Y2=0
cc_1596 Z N_A_2693_297#_c_2717_n 0.00349489f $X=16.805 $Y=1.785 $X2=0 $Y2=0
cc_1597 N_Z_c_2346_n N_A_2693_297#_c_2717_n 0.0150524f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_1598 N_Z_c_2221_n N_A_2693_297#_c_2718_n 0.0209902f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_1599 N_Z_c_2445_n N_A_2693_297#_c_2718_n 6.74054e-19 $X=17.095 $Y=1.87 $X2=0
+ $Y2=0
cc_1600 N_Z_c_2346_n N_A_2693_297#_c_2718_n 0.0228406f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_1601 N_Z_c_2221_n N_A_4219_311#_M1039_d 2.07056e-19 $X=21.545 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_1602 N_Z_c_2398_n N_A_4219_311#_M1048_d 3.24931e-19 $X=22.485 $Y=1.87 $X2=0
+ $Y2=0
cc_1603 N_Z_c_2221_n N_A_4219_311#_c_2814_n 0.0209902f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_1604 Z N_A_4219_311#_c_2814_n 6.74054e-19 $X=21.665 $Y=1.785 $X2=0 $Y2=0
cc_1605 N_Z_c_2400_n N_A_4219_311#_c_2814_n 0.0228406f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_1606 N_Z_M1039_s N_A_4219_311#_c_2815_n 0.00176676f $X=21.545 $Y=1.555 $X2=0
+ $Y2=0
cc_1607 N_Z_c_2221_n N_A_4219_311#_c_2815_n 0.00349489f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_1608 N_Z_c_2398_n N_A_4219_311#_c_2815_n 0.00349489f $X=22.485 $Y=1.87 $X2=0
+ $Y2=0
cc_1609 Z N_A_4219_311#_c_2815_n 9.16304e-19 $X=21.665 $Y=1.785 $X2=0 $Y2=0
cc_1610 N_Z_c_2400_n N_A_4219_311#_c_2815_n 0.0150524f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_1611 N_Z_c_2201_n N_A_4219_311#_c_2817_n 0.0192125f $X=22.465 $Y=1.215 $X2=0
+ $Y2=0
cc_1612 N_Z_c_2212_n N_A_4219_311#_c_2817_n 0.0024794f $X=21.79 $Y=1.215 $X2=0
+ $Y2=0
cc_1613 N_Z_c_2398_n N_A_4219_311#_c_2817_n 0.0189041f $X=22.485 $Y=1.87 $X2=0
+ $Y2=0
cc_1614 N_Z_c_2449_n N_A_4219_311#_c_2817_n 6.68271e-19 $X=22.63 $Y=1.87 $X2=0
+ $Y2=0
cc_1615 Z N_A_4219_311#_c_2817_n 6.68271e-19 $X=21.665 $Y=1.785 $X2=0 $Y2=0
cc_1616 N_Z_c_2400_n N_A_4219_311#_c_2817_n 0.0247248f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_1617 N_Z_c_2407_n N_A_4219_311#_c_2817_n 0.0247248f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_1618 N_Z_M1060_s N_A_4219_311#_c_2818_n 0.00176676f $X=22.485 $Y=1.555 $X2=0
+ $Y2=0
cc_1619 N_Z_c_2398_n N_A_4219_311#_c_2818_n 0.00349489f $X=22.485 $Y=1.87 $X2=0
+ $Y2=0
cc_1620 N_Z_c_2449_n N_A_4219_311#_c_2818_n 9.16304e-19 $X=22.63 $Y=1.87 $X2=0
+ $Y2=0
cc_1621 N_Z_c_2407_n N_A_4219_311#_c_2818_n 0.0151266f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_1622 N_Z_c_2449_n N_A_4219_311#_c_2819_n 0.00168706f $X=22.63 $Y=1.87 $X2=0
+ $Y2=0
cc_1623 N_Z_c_2407_n N_A_4219_311#_c_2821_n 0.00915958f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_1624 N_Z_c_2203_n N_A_119_47#_c_3247_n 0.00799417f $X=3.03 $Y=0.68 $X2=0
+ $Y2=0
cc_1625 N_Z_M1015_s N_A_119_47#_c_3249_n 0.00165831f $X=2.895 $Y=0.33 $X2=0
+ $Y2=0
cc_1626 N_Z_c_2192_n N_A_119_47#_c_3249_n 0.00133192f $X=3.705 $Y=1.215 $X2=0
+ $Y2=0
cc_1627 N_Z_c_2203_n N_A_119_47#_c_3249_n 0.0157607f $X=3.03 $Y=0.68 $X2=0 $Y2=0
cc_1628 N_Z_c_2204_n N_A_119_47#_c_3249_n 0.00293855f $X=3.13 $Y=1.215 $X2=0
+ $Y2=0
cc_1629 N_Z_c_2192_n N_A_119_47#_c_3274_n 0.00918654f $X=3.705 $Y=1.215 $X2=0
+ $Y2=0
cc_1630 N_Z_M1028_s N_A_119_47#_c_3251_n 0.00165831f $X=3.735 $Y=0.33 $X2=0
+ $Y2=0
cc_1631 N_Z_c_2192_n N_A_119_47#_c_3251_n 0.00405549f $X=3.705 $Y=1.215 $X2=0
+ $Y2=0
cc_1632 N_Z_c_2193_n N_A_119_47#_c_3251_n 0.015949f $X=3.87 $Y=0.68 $X2=0 $Y2=0
cc_1633 N_Z_c_2205_n N_A_119_47#_c_3251_n 0.00443806f $X=3.97 $Y=1.215 $X2=0
+ $Y2=0
cc_1634 N_Z_c_2205_n N_A_119_47#_c_3252_n 0.00158445f $X=3.97 $Y=1.215 $X2=0
+ $Y2=0
cc_1635 N_Z_c_2206_n N_A_1693_66#_c_3329_n 0.00158445f $X=8.91 $Y=1.215 $X2=0
+ $Y2=0
cc_1636 N_Z_M1007_d N_A_1693_66#_c_3330_n 0.00165831f $X=8.875 $Y=0.33 $X2=0
+ $Y2=0
cc_1637 N_Z_c_2194_n N_A_1693_66#_c_3330_n 0.015949f $X=9.01 $Y=0.68 $X2=0 $Y2=0
cc_1638 N_Z_c_2195_n N_A_1693_66#_c_3330_n 0.00405549f $X=9.585 $Y=1.215 $X2=0
+ $Y2=0
cc_1639 N_Z_c_2206_n N_A_1693_66#_c_3330_n 0.00443806f $X=8.91 $Y=1.215 $X2=0
+ $Y2=0
cc_1640 N_Z_c_2195_n N_A_1693_66#_c_3351_n 0.00918654f $X=9.585 $Y=1.215 $X2=0
+ $Y2=0
cc_1641 N_Z_M1026_d N_A_1693_66#_c_3332_n 0.00165831f $X=9.715 $Y=0.33 $X2=0
+ $Y2=0
cc_1642 N_Z_c_2195_n N_A_1693_66#_c_3332_n 0.00133192f $X=9.585 $Y=1.215 $X2=0
+ $Y2=0
cc_1643 N_Z_c_2207_n N_A_1693_66#_c_3332_n 0.00293855f $X=9.75 $Y=1.215 $X2=0
+ $Y2=0
cc_1644 N_Z_c_2208_n N_A_1693_66#_c_3332_n 0.0157607f $X=9.85 $Y=0.68 $X2=0
+ $Y2=0
cc_1645 N_Z_c_2208_n N_A_1693_66#_c_3335_n 0.00799417f $X=9.85 $Y=0.68 $X2=0
+ $Y2=0
cc_1646 N_Z_c_2209_n N_A_2695_47#_c_3414_n 0.00799417f $X=15.91 $Y=0.68 $X2=0
+ $Y2=0
cc_1647 N_Z_M1008_d N_A_2695_47#_c_3416_n 0.00165831f $X=15.775 $Y=0.33 $X2=0
+ $Y2=0
cc_1648 N_Z_c_2198_n N_A_2695_47#_c_3416_n 0.00133192f $X=16.585 $Y=1.215 $X2=0
+ $Y2=0
cc_1649 N_Z_c_2209_n N_A_2695_47#_c_3416_n 0.0157607f $X=15.91 $Y=0.68 $X2=0
+ $Y2=0
cc_1650 N_Z_c_2210_n N_A_2695_47#_c_3416_n 0.00293855f $X=16.01 $Y=1.215 $X2=0
+ $Y2=0
cc_1651 N_Z_c_2198_n N_A_2695_47#_c_3441_n 0.00918654f $X=16.585 $Y=1.215 $X2=0
+ $Y2=0
cc_1652 N_Z_M1030_d N_A_2695_47#_c_3418_n 0.00165831f $X=16.615 $Y=0.33 $X2=0
+ $Y2=0
cc_1653 N_Z_c_2198_n N_A_2695_47#_c_3418_n 0.00405549f $X=16.585 $Y=1.215 $X2=0
+ $Y2=0
cc_1654 N_Z_c_2199_n N_A_2695_47#_c_3418_n 0.015949f $X=16.75 $Y=0.68 $X2=0
+ $Y2=0
cc_1655 N_Z_c_2211_n N_A_2695_47#_c_3418_n 0.00443806f $X=16.85 $Y=1.215 $X2=0
+ $Y2=0
cc_1656 N_Z_c_2211_n N_A_2695_47#_c_3419_n 0.00158445f $X=16.85 $Y=1.215 $X2=0
+ $Y2=0
cc_1657 N_Z_c_2212_n N_A_4269_66#_c_3496_n 0.00158445f $X=21.79 $Y=1.215 $X2=0
+ $Y2=0
cc_1658 N_Z_M1011_d N_A_4269_66#_c_3497_n 0.00165831f $X=21.755 $Y=0.33 $X2=0
+ $Y2=0
cc_1659 N_Z_c_2200_n N_A_4269_66#_c_3497_n 0.015949f $X=21.89 $Y=0.68 $X2=0
+ $Y2=0
cc_1660 N_Z_c_2201_n N_A_4269_66#_c_3497_n 0.00405549f $X=22.465 $Y=1.215 $X2=0
+ $Y2=0
cc_1661 N_Z_c_2212_n N_A_4269_66#_c_3497_n 0.00443806f $X=21.79 $Y=1.215 $X2=0
+ $Y2=0
cc_1662 N_Z_c_2201_n N_A_4269_66#_c_3518_n 0.00918654f $X=22.465 $Y=1.215 $X2=0
+ $Y2=0
cc_1663 N_Z_M1022_d N_A_4269_66#_c_3499_n 0.00165831f $X=22.595 $Y=0.33 $X2=0
+ $Y2=0
cc_1664 N_Z_c_2201_n N_A_4269_66#_c_3499_n 0.00133192f $X=22.465 $Y=1.215 $X2=0
+ $Y2=0
cc_1665 N_Z_c_2213_n N_A_4269_66#_c_3499_n 0.00293855f $X=22.63 $Y=1.215 $X2=0
+ $Y2=0
cc_1666 N_Z_c_2214_n N_A_4269_66#_c_3499_n 0.0157607f $X=22.73 $Y=0.68 $X2=0
+ $Y2=0
cc_1667 N_Z_c_2214_n N_A_4269_66#_c_3502_n 0.00799417f $X=22.73 $Y=0.68 $X2=0
+ $Y2=0
cc_1668 N_A_1643_311#_c_2613_n N_A_1693_66#_c_3334_n 0.0147893f $X=11.045
+ $Y=1.58 $X2=0 $Y2=0
cc_1669 N_A_1643_311#_c_2613_n N_A_1693_66#_c_3335_n 0.00239279f $X=11.045
+ $Y=1.58 $X2=0 $Y2=0
cc_1670 N_A_1643_311#_c_2614_n N_A_1693_66#_c_3335_n 0.00761509f $X=10.385
+ $Y=1.58 $X2=0 $Y2=0
cc_1671 N_A_1643_311#_c_2647_n N_A_1693_66#_c_3337_n 6.95815e-19 $X=11.21
+ $Y=1.66 $X2=0 $Y2=0
cc_1672 N_A_2693_297#_c_2712_n N_A_2695_47#_c_3414_n 0.0247972f $X=15.375
+ $Y=1.58 $X2=0 $Y2=0
cc_1673 N_A_2693_297#_c_2736_n N_A_2695_47#_c_3420_n 6.95815e-19 $X=14.55
+ $Y=1.66 $X2=0 $Y2=0
cc_1674 N_A_4219_311#_c_2820_n N_A_4269_66#_c_3501_n 0.0147893f $X=23.925
+ $Y=1.58 $X2=0 $Y2=0
cc_1675 N_A_4219_311#_c_2820_n N_A_4269_66#_c_3502_n 0.00239279f $X=23.925
+ $Y=1.58 $X2=0 $Y2=0
cc_1676 N_A_4219_311#_c_2821_n N_A_4269_66#_c_3502_n 0.00761509f $X=23.265
+ $Y=1.58 $X2=0 $Y2=0
cc_1677 N_A_4219_311#_c_2853_n N_A_4269_66#_c_3504_n 6.95815e-19 $X=24.09
+ $Y=1.66 $X2=0 $Y2=0
cc_1678 VGND N_A_119_47#_M1024_s 0.00215201f $X=25.445 $Y=-0.085 $X2=-0.19
+ $Y2=-0.24
cc_1679 VGND N_A_119_47#_M1073_s 0.00215201f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1680 VGND N_A_119_47#_c_3254_n 0.0121968f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1681 N_VGND_c_2952_n N_A_119_47#_c_3254_n 0.0188215f $X=1.065 $Y=0 $X2=0
+ $Y2=0
cc_1682 N_VGND_M1057_d N_A_119_47#_c_3257_n 0.00501873f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_1683 N_VGND_c_2908_n N_A_119_47#_c_3257_n 0.0199861f $X=1.2 $Y=0.38 $X2=0
+ $Y2=0
cc_1684 N_VGND_c_2909_n N_A_119_47#_c_3257_n 0.0020257f $X=2.005 $Y=0 $X2=0
+ $Y2=0
cc_1685 VGND N_A_119_47#_c_3257_n 0.00880092f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1686 N_VGND_c_2952_n N_A_119_47#_c_3257_n 0.0020257f $X=1.065 $Y=0 $X2=0
+ $Y2=0
cc_1687 N_VGND_c_2909_n N_A_119_47#_c_3265_n 0.0188215f $X=2.005 $Y=0 $X2=0
+ $Y2=0
cc_1688 VGND N_A_119_47#_c_3265_n 0.0121968f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1689 N_VGND_M1078_d N_A_119_47#_c_3247_n 0.00692362f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_1690 N_VGND_c_2909_n N_A_119_47#_c_3247_n 0.0020257f $X=2.005 $Y=0 $X2=0
+ $Y2=0
cc_1691 N_VGND_c_2910_n N_A_119_47#_c_3247_n 0.0190091f $X=2.09 $Y=0.38 $X2=0
+ $Y2=0
cc_1692 N_VGND_c_2931_n N_A_119_47#_c_3247_n 0.00262594f $X=4.96 $Y=0 $X2=0
+ $Y2=0
cc_1693 VGND N_A_119_47#_c_3247_n 0.00940109f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1694 N_VGND_c_2910_n N_A_119_47#_c_3248_n 0.00959666f $X=2.09 $Y=0.38 $X2=0
+ $Y2=0
cc_1695 N_VGND_c_2931_n N_A_119_47#_c_3249_n 0.0422314f $X=4.96 $Y=0 $X2=0 $Y2=0
cc_1696 VGND N_A_119_47#_c_3249_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1697 N_VGND_c_2910_n N_A_119_47#_c_3250_n 0.0147456f $X=2.09 $Y=0.38 $X2=0
+ $Y2=0
cc_1698 N_VGND_c_2931_n N_A_119_47#_c_3250_n 0.0192461f $X=4.96 $Y=0 $X2=0 $Y2=0
cc_1699 VGND N_A_119_47#_c_3250_n 0.0103774f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1700 N_VGND_c_2911_n N_A_119_47#_c_3251_n 0.00694621f $X=5.165 $Y=0.445 $X2=0
+ $Y2=0
cc_1701 N_VGND_c_2931_n N_A_119_47#_c_3251_n 0.0589406f $X=4.96 $Y=0 $X2=0 $Y2=0
cc_1702 VGND N_A_119_47#_c_3251_n 0.030408f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1703 N_VGND_c_2911_n N_A_119_47#_c_3252_n 0.00696245f $X=5.165 $Y=0.445 $X2=0
+ $Y2=0
cc_1704 N_VGND_c_2931_n N_A_119_47#_c_3287_n 0.0113631f $X=4.96 $Y=0 $X2=0 $Y2=0
cc_1705 VGND N_A_119_47#_c_3287_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1706 VGND N_A_1693_66#_M1017_s 0.00215201f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1707 VGND N_A_1693_66#_M1049_s 0.00215201f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1708 N_VGND_c_2914_n N_A_1693_66#_c_3329_n 0.00696245f $X=7.715 $Y=0.445
+ $X2=0 $Y2=0
cc_1709 N_VGND_c_2939_n N_A_1693_66#_c_3330_n 0.0422314f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_1710 VGND N_A_1693_66#_c_3330_n 0.0219908f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1711 N_VGND_c_2914_n N_A_1693_66#_c_3331_n 0.00694621f $X=7.715 $Y=0.445
+ $X2=0 $Y2=0
cc_1712 N_VGND_c_2939_n N_A_1693_66#_c_3331_n 0.0167092f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_1713 VGND N_A_1693_66#_c_3331_n 0.00841721f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1714 N_VGND_c_2915_n N_A_1693_66#_c_3332_n 0.0147456f $X=10.79 $Y=0.38 $X2=0
+ $Y2=0
cc_1715 N_VGND_c_2939_n N_A_1693_66#_c_3332_n 0.0614775f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_1716 VGND N_A_1693_66#_c_3332_n 0.0325967f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1717 N_VGND_c_2915_n N_A_1693_66#_c_3333_n 0.00959666f $X=10.79 $Y=0.38 $X2=0
+ $Y2=0
cc_1718 N_VGND_M1017_d N_A_1693_66#_c_3334_n 0.00692362f $X=10.665 $Y=0.235
+ $X2=0 $Y2=0
cc_1719 N_VGND_c_2915_n N_A_1693_66#_c_3334_n 0.0190091f $X=10.79 $Y=0.38 $X2=0
+ $Y2=0
cc_1720 N_VGND_c_2939_n N_A_1693_66#_c_3334_n 0.00262594f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_1721 VGND N_A_1693_66#_c_3334_n 0.00940109f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1722 N_VGND_c_2953_n N_A_1693_66#_c_3334_n 0.0020257f $X=11.545 $Y=0 $X2=0
+ $Y2=0
cc_1723 VGND N_A_1693_66#_c_3354_n 0.0121968f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1724 N_VGND_c_2953_n N_A_1693_66#_c_3354_n 0.0188215f $X=11.545 $Y=0 $X2=0
+ $Y2=0
cc_1725 N_VGND_M1029_d N_A_1693_66#_c_3336_n 0.00501873f $X=11.495 $Y=0.235
+ $X2=0 $Y2=0
cc_1726 N_VGND_c_2916_n N_A_1693_66#_c_3336_n 0.0199861f $X=11.68 $Y=0.38 $X2=0
+ $Y2=0
cc_1727 VGND N_A_1693_66#_c_3336_n 0.00880092f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1728 N_VGND_c_2953_n N_A_1693_66#_c_3336_n 0.0020257f $X=11.545 $Y=0 $X2=0
+ $Y2=0
cc_1729 N_VGND_c_2954_n N_A_1693_66#_c_3336_n 0.0020257f $X=12.485 $Y=0 $X2=0
+ $Y2=0
cc_1730 VGND N_A_1693_66#_c_3363_n 0.0121968f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1731 N_VGND_c_2954_n N_A_1693_66#_c_3363_n 0.0188215f $X=12.485 $Y=0 $X2=0
+ $Y2=0
cc_1732 N_VGND_c_2939_n N_A_1693_66#_c_3348_n 0.0113631f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_1733 VGND N_A_1693_66#_c_3348_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1734 VGND N_A_2695_47#_M1002_d 0.00215201f $X=25.445 $Y=-0.085 $X2=-0.19
+ $Y2=-0.24
cc_1735 VGND N_A_2695_47#_M1034_d 0.00215201f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1736 VGND N_A_2695_47#_c_3421_n 0.0121968f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1737 N_VGND_c_2955_n N_A_2695_47#_c_3421_n 0.0188215f $X=13.945 $Y=0 $X2=0
+ $Y2=0
cc_1738 N_VGND_M1021_s N_A_2695_47#_c_3424_n 0.00501873f $X=13.895 $Y=0.235
+ $X2=0 $Y2=0
cc_1739 N_VGND_c_2920_n N_A_2695_47#_c_3424_n 0.0199861f $X=14.08 $Y=0.38 $X2=0
+ $Y2=0
cc_1740 N_VGND_c_2921_n N_A_2695_47#_c_3424_n 0.0020257f $X=14.885 $Y=0 $X2=0
+ $Y2=0
cc_1741 VGND N_A_2695_47#_c_3424_n 0.00880092f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1742 N_VGND_c_2955_n N_A_2695_47#_c_3424_n 0.0020257f $X=13.945 $Y=0 $X2=0
+ $Y2=0
cc_1743 N_VGND_c_2921_n N_A_2695_47#_c_3432_n 0.0188215f $X=14.885 $Y=0 $X2=0
+ $Y2=0
cc_1744 VGND N_A_2695_47#_c_3432_n 0.0121968f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1745 N_VGND_M1052_s N_A_2695_47#_c_3414_n 0.00692362f $X=14.835 $Y=0.235
+ $X2=0 $Y2=0
cc_1746 N_VGND_c_2921_n N_A_2695_47#_c_3414_n 0.0020257f $X=14.885 $Y=0 $X2=0
+ $Y2=0
cc_1747 N_VGND_c_2922_n N_A_2695_47#_c_3414_n 0.0190091f $X=14.97 $Y=0.38 $X2=0
+ $Y2=0
cc_1748 N_VGND_c_2941_n N_A_2695_47#_c_3414_n 0.00262594f $X=17.84 $Y=0 $X2=0
+ $Y2=0
cc_1749 VGND N_A_2695_47#_c_3414_n 0.00940109f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1750 N_VGND_c_2922_n N_A_2695_47#_c_3415_n 0.00959666f $X=14.97 $Y=0.38 $X2=0
+ $Y2=0
cc_1751 N_VGND_c_2941_n N_A_2695_47#_c_3416_n 0.0422314f $X=17.84 $Y=0 $X2=0
+ $Y2=0
cc_1752 VGND N_A_2695_47#_c_3416_n 0.0222193f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1753 N_VGND_c_2922_n N_A_2695_47#_c_3417_n 0.0147456f $X=14.97 $Y=0.38 $X2=0
+ $Y2=0
cc_1754 N_VGND_c_2941_n N_A_2695_47#_c_3417_n 0.0192461f $X=17.84 $Y=0 $X2=0
+ $Y2=0
cc_1755 VGND N_A_2695_47#_c_3417_n 0.0103774f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1756 N_VGND_c_2923_n N_A_2695_47#_c_3418_n 0.00694621f $X=18.045 $Y=0.445
+ $X2=0 $Y2=0
cc_1757 N_VGND_c_2941_n N_A_2695_47#_c_3418_n 0.0589406f $X=17.84 $Y=0 $X2=0
+ $Y2=0
cc_1758 VGND N_A_2695_47#_c_3418_n 0.030408f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1759 N_VGND_c_2923_n N_A_2695_47#_c_3419_n 0.00696245f $X=18.045 $Y=0.445
+ $X2=0 $Y2=0
cc_1760 N_VGND_c_2941_n N_A_2695_47#_c_3454_n 0.0113631f $X=17.84 $Y=0 $X2=0
+ $Y2=0
cc_1761 VGND N_A_2695_47#_c_3454_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1762 VGND N_A_4269_66#_M1013_s 0.00215201f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1763 VGND N_A_4269_66#_M1040_s 0.00215201f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1764 N_VGND_c_2926_n N_A_4269_66#_c_3496_n 0.00696245f $X=20.595 $Y=0.445
+ $X2=0 $Y2=0
cc_1765 N_VGND_c_2949_n N_A_4269_66#_c_3497_n 0.0422314f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_1766 VGND N_A_4269_66#_c_3497_n 0.0219908f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1767 N_VGND_c_2926_n N_A_4269_66#_c_3498_n 0.00694621f $X=20.595 $Y=0.445
+ $X2=0 $Y2=0
cc_1768 N_VGND_c_2949_n N_A_4269_66#_c_3498_n 0.0167092f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_1769 VGND N_A_4269_66#_c_3498_n 0.00841721f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1770 N_VGND_c_2927_n N_A_4269_66#_c_3499_n 0.0147456f $X=23.67 $Y=0.38 $X2=0
+ $Y2=0
cc_1771 N_VGND_c_2949_n N_A_4269_66#_c_3499_n 0.0614775f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_1772 VGND N_A_4269_66#_c_3499_n 0.0325967f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1773 N_VGND_c_2927_n N_A_4269_66#_c_3500_n 0.00959666f $X=23.67 $Y=0.38 $X2=0
+ $Y2=0
cc_1774 N_VGND_M1013_d N_A_4269_66#_c_3501_n 0.00692362f $X=23.545 $Y=0.235
+ $X2=0 $Y2=0
cc_1775 N_VGND_c_2927_n N_A_4269_66#_c_3501_n 0.0190091f $X=23.67 $Y=0.38 $X2=0
+ $Y2=0
cc_1776 N_VGND_c_2949_n N_A_4269_66#_c_3501_n 0.00262594f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_1777 VGND N_A_4269_66#_c_3501_n 0.00940109f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1778 N_VGND_c_2956_n N_A_4269_66#_c_3501_n 0.0020257f $X=24.425 $Y=0 $X2=0
+ $Y2=0
cc_1779 VGND N_A_4269_66#_c_3521_n 0.0121968f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1780 N_VGND_c_2956_n N_A_4269_66#_c_3521_n 0.0188215f $X=24.425 $Y=0 $X2=0
+ $Y2=0
cc_1781 N_VGND_M1032_d N_A_4269_66#_c_3503_n 0.00501873f $X=24.375 $Y=0.235
+ $X2=0 $Y2=0
cc_1782 N_VGND_c_2928_n N_A_4269_66#_c_3503_n 0.0199861f $X=24.56 $Y=0.38 $X2=0
+ $Y2=0
cc_1783 VGND N_A_4269_66#_c_3503_n 0.00880092f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1784 N_VGND_c_2956_n N_A_4269_66#_c_3503_n 0.0020257f $X=24.425 $Y=0 $X2=0
+ $Y2=0
cc_1785 N_VGND_c_2957_n N_A_4269_66#_c_3503_n 0.0020257f $X=25.365 $Y=0 $X2=0
+ $Y2=0
cc_1786 VGND N_A_4269_66#_c_3530_n 0.0121968f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
cc_1787 N_VGND_c_2957_n N_A_4269_66#_c_3530_n 0.0188215f $X=25.365 $Y=0 $X2=0
+ $Y2=0
cc_1788 N_VGND_c_2949_n N_A_4269_66#_c_3515_n 0.0113631f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_1789 VGND N_A_4269_66#_c_3515_n 0.00572388f $X=25.445 $Y=-0.085 $X2=0 $Y2=0
