# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o2bb2a_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.820000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.615000 1.075000 3.995000 1.445000 ;
        RECT 3.615000 1.445000 5.465000 1.615000 ;
        RECT 5.055000 1.075000 5.465000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 1.075000 4.885000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.625000 1.445000 ;
        RECT 0.085000 1.445000 2.095000 1.615000 ;
        RECT 1.715000 1.075000 2.095000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 1.075000 1.445000 1.275000 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.735000 0.275000 6.115000 0.725000 ;
        RECT 5.735000 0.725000 7.710000 0.905000 ;
        RECT 5.825000 1.785000 7.015000 1.955000 ;
        RECT 5.825000 1.955000 6.075000 2.465000 ;
        RECT 6.675000 0.275000 7.055000 0.725000 ;
        RECT 6.765000 1.415000 7.710000 1.655000 ;
        RECT 6.765000 1.655000 7.015000 1.785000 ;
        RECT 6.765000 1.955000 7.015000 2.465000 ;
        RECT 7.405000 0.905000 7.710000 1.415000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.725000 ;
      RECT 0.095000  0.725000 1.365000 0.735000 ;
      RECT 0.095000  0.735000 2.225000 0.905000 ;
      RECT 0.140000  1.795000 0.345000 2.635000 ;
      RECT 0.605000  1.785000 0.855000 2.295000 ;
      RECT 0.605000  2.295000 1.795000 2.465000 ;
      RECT 0.645000  0.085000 0.815000 0.555000 ;
      RECT 0.985000  0.255000 1.365000 0.725000 ;
      RECT 1.075000  1.785000 2.865000 1.955000 ;
      RECT 1.075000  1.955000 1.325000 2.125000 ;
      RECT 1.545000  2.125000 1.795000 2.295000 ;
      RECT 1.585000  0.085000 1.755000 0.555000 ;
      RECT 1.925000  0.255000 3.245000 0.475000 ;
      RECT 1.925000  0.475000 2.225000 0.735000 ;
      RECT 2.015000  2.125000 2.265000 2.635000 ;
      RECT 2.265000  1.075000 2.695000 1.415000 ;
      RECT 2.265000  1.415000 2.865000 1.785000 ;
      RECT 2.395000  0.645000 2.775000 0.815000 ;
      RECT 2.395000  0.815000 2.695000 1.075000 ;
      RECT 2.485000  1.955000 2.865000 1.965000 ;
      RECT 2.485000  1.965000 2.775000 2.465000 ;
      RECT 2.865000  1.075000 3.445000 1.245000 ;
      RECT 2.995000  2.135000 3.725000 2.635000 ;
      RECT 3.255000  0.725000 4.705000 0.905000 ;
      RECT 3.255000  0.905000 3.445000 1.075000 ;
      RECT 3.255000  1.245000 3.445000 1.785000 ;
      RECT 3.255000  1.785000 5.135000 1.965000 ;
      RECT 3.515000  0.085000 3.685000 0.555000 ;
      RECT 3.855000  0.305000 5.175000 0.475000 ;
      RECT 3.945000  1.965000 4.195000 2.125000 ;
      RECT 4.325000  0.645000 4.705000 0.725000 ;
      RECT 4.415000  2.135000 4.665000 2.635000 ;
      RECT 4.885000  1.965000 5.135000 2.465000 ;
      RECT 4.925000  0.475000 5.175000 0.895000 ;
      RECT 5.355000  1.795000 5.605000 2.635000 ;
      RECT 5.395000  0.085000 5.565000 0.895000 ;
      RECT 5.665000  1.075000 7.085000 1.245000 ;
      RECT 5.665000  1.245000 6.005000 1.615000 ;
      RECT 6.295000  2.165000 6.545000 2.635000 ;
      RECT 6.335000  0.085000 6.505000 0.555000 ;
      RECT 7.235000  1.825000 7.485000 2.635000 ;
      RECT 7.275000  0.085000 7.445000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.695000  1.435000 2.865000 1.605000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.725000  1.445000 5.895000 1.615000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 2.635000 1.385000 2.975000 1.460000 ;
      RECT 2.635000 1.460000 5.960000 1.600000 ;
      RECT 2.635000 1.600000 2.975000 1.635000 ;
      RECT 5.665000 1.395000 5.960000 1.460000 ;
      RECT 5.665000 1.600000 5.960000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2a_4
END LIBRARY
