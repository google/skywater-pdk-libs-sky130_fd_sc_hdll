* NGSPICE file created from sky130_fd_sc_hdll__diode_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__diode_4 DIODE VGND VNB VPB VPWR
D0 VNB DIODE ndiode p=9.88e+06u a=1.0557e+12p
.ends

