* NGSPICE file created from sky130_fd_sc_hdll__inv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__inv_2 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=5.4e+11p ps=5.08e+06u
M1001 VGND A Y VNB nshort w=650000u l=150000u
+  ad=3.705e+11p pd=3.74e+06u as=2.08e+11p ps=1.94e+06u
M1002 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

