* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor4_6 A B C D VGND VNB VPB VPWR Y
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=2.01e+12p ps=1.802e+07u
M1001 a_1263_297# C a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.02e+12p pd=1.804e+07u as=1.74e+12p ps=1.548e+07u
M1002 Y D a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=0p ps=0u
M1003 VGND B Y VNB nshort w=650000u l=150000u
+  ad=3.419e+12p pd=2.742e+07u as=2.106e+12p ps=2.208e+07u
M1004 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_685_297# C a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_685_297# C a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1263_297# C a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_685_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1263_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_297# B a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1263_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y D a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y D a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_27_297# B a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_685_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1263_297# D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_685_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_685_297# C a_1263_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_1263_297# C a_685_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND D Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
