* File: sky130_fd_sc_hdll__inputiso1n_1.pex.spice
* Created: Wed Sep  2 08:32:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%SLEEP_B 1 3 6 8 13 16
r28 13 14 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r29 11 13 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r30 8 16 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.2 $X2=0.23
+ $Y2=1.2
r31 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r32 4 14 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r33 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.475
r34 1 13 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r35 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%A_27_53# 1 2 7 9 12 16 18 19 22 26 29
+ 34
c49 26 0 7.50303e-20 $X=1.27 $Y=1.16
r50 34 35 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=1.505 $Y=1.202
+ $X2=1.53 $Y2=1.202
r51 27 34 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=1.27 $Y=1.202
+ $X2=1.505 $Y2=1.202
r52 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r53 24 32 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.16
+ $X2=0.77 $Y2=1.325
r54 24 29 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.77 $Y=1.16
+ $X2=0.77 $Y2=0.82
r55 24 26 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.895 $Y=1.16
+ $X2=1.27 $Y2=1.16
r56 22 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=1.62
+ $X2=0.73 $Y2=1.325
r57 18 29 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.77 $Y2=0.82
r58 18 19 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.42 $Y2=0.82
r59 14 19 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.42 $Y2=0.82
r60 14 16 10.7809 $w=3.08e-07 $l=2.9e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.265 $Y2=0.445
r61 10 35 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=1.202
r62 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=0.475
r63 7 34 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.505 $Y=1.41
+ $X2=1.505 $Y2=1.202
r64 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.505 $Y=1.41
+ $X2=1.505 $Y2=1.695
r65 2 22 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.62
r66 1 16 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%A 1 3 4 5 8 11 14 16 22 26
c46 11 0 7.50303e-20 $X=2 $Y=0.475
c47 4 0 8.49032e-20 $X=1.975 $Y=1.31
r48 20 26 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.06 $Y=2.25
+ $X2=1.155 $Y2=2.25
r49 19 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=2.28
+ $X2=1.225 $Y2=2.28
r50 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=2.28 $X2=1.06 $Y2=2.28
r51 16 26 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.205 $Y=2.25
+ $X2=1.155 $Y2=2.25
r52 11 13 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2 $Y=0.475 $X2=2
+ $Y2=1.015
r53 6 14 101.939 $w=2e-07 $l=3.05e-07 $layer=POLY_cond $X=1.975 $Y=2.035
+ $X2=1.975 $Y2=2.34
r54 6 8 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.975 $Y=2.035
+ $X2=1.975 $Y2=1.695
r55 5 8 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.975 $Y=1.41
+ $X2=1.975 $Y2=1.695
r56 4 5 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.975 $Y=1.31 $X2=1.975
+ $Y2=1.41
r57 3 13 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.975 $Y=1.115 $X2=1.975
+ $Y2=1.015
r58 3 4 64.6575 $w=2e-07 $l=1.95e-07 $layer=POLY_cond $X=1.975 $Y=1.115
+ $X2=1.975 $Y2=1.31
r59 1 14 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.875 $Y=2.34 $X2=1.975
+ $Y2=2.34
r60 1 22 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.875 $Y=2.34
+ $X2=1.225 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%A_229_297# 1 2 7 9 10 12 13 17 19 20
+ 24 26
c58 24 0 1.12758e-19 $X=2.42 $Y=1.16
r59 26 29 2.88111 $w=4.18e-07 $l=1.05e-07 $layer=LI1_cond $X=1.25 $Y=1.58
+ $X2=1.25 $Y2=1.685
r60 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.16 $X2=2.42 $Y2=1.16
r61 22 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.42 $Y=1.495
+ $X2=2.42 $Y2=1.16
r62 21 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.42 $Y=0.825
+ $X2=2.42 $Y2=1.16
r63 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.335 $Y=0.74
+ $X2=2.42 $Y2=0.825
r64 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.335 $Y=0.74
+ $X2=1.825 $Y2=0.74
r65 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.74 $Y=0.655
+ $X2=1.825 $Y2=0.74
r66 15 17 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.74 $Y=0.655
+ $X2=1.74 $Y2=0.47
r67 14 26 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.46 $Y=1.58 $X2=1.25
+ $Y2=1.58
r68 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.335 $Y=1.58
+ $X2=2.42 $Y2=1.495
r69 13 14 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.335 $Y=1.58
+ $X2=1.46 $Y2=1.58
r70 10 25 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.54 $Y=0.995
+ $X2=2.45 $Y2=1.16
r71 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.54 $Y=0.995
+ $X2=2.54 $Y2=0.56
r72 7 25 47.6478 $w=3.03e-07 $l=2.80624e-07 $layer=POLY_cond $X=2.515 $Y=1.41
+ $X2=2.45 $Y2=1.16
r73 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.515 $Y=1.41
+ $X2=2.515 $Y2=1.985
r74 2 29 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.485 $X2=1.27 $Y2=1.685
r75 1 17 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.265 $X2=1.74 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%VPWR 1 2 7 9 13 16 17 18 28 29
c32 2 0 1.12758e-19 $X=2.065 $Y=1.485
r33 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r34 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r35 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r36 23 26 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 22 25 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r38 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r39 20 32 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r40 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 18 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 18 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r43 16 25 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 16 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.265 $Y2=2.72
r45 15 28 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.405 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 15 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.405 $Y=2.72
+ $X2=2.265 $Y2=2.72
r47 11 17 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.265 $Y=2.635
+ $X2=2.265 $Y2=2.72
r48 11 13 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.265 $Y=2.635
+ $X2=2.265 $Y2=2
r49 7 32 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r50 7 9 44.064 $w=2.53e-07 $l=9.75e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=1.66
r51 2 13 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=2.065
+ $Y=1.485 $X2=2.275 $Y2=2
r52 1 9 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%X 1 2 12 14 15 16
r18 14 16 4.2114 $w=4.03e-07 $l=1.48e-07 $layer=LI1_cond $X=2.877 $Y=1.697
+ $X2=2.877 $Y2=1.845
r19 14 15 9.72165 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=2.877 $Y=1.697
+ $X2=2.877 $Y2=1.495
r20 10 12 7.84997 $w=3.43e-07 $l=2.35e-07 $layer=LI1_cond $X=2.76 $Y=0.587
+ $X2=2.995 $Y2=0.587
r21 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.995 $Y=0.76
+ $X2=2.995 $Y2=0.587
r22 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.995 $Y=0.76
+ $X2=2.995 $Y2=1.495
r23 2 16 300 $w=1.7e-07 $l=4.30581e-07 $layer=licon1_PDIFF $count=2 $X=2.605
+ $Y=1.485 $X2=2.76 $Y2=1.845
r24 1 10 182 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.235 $X2=2.76 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%VGND 1 2 9 11 15 16 19 27 30
r40 30 33 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.21
+ $Y2=0.4
r41 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r42 26 27 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=0.24
+ $X2=1.375 $Y2=0.24
r43 24 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r44 23 26 1.10407 $w=6.48e-07 $l=6e-08 $layer=LI1_cond $X=1.15 $Y=0.24 $X2=1.21
+ $Y2=0.24
r45 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r46 20 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r47 19 23 8.46455 $w=6.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.24
+ $X2=1.15 $Y2=0.24
r48 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r49 16 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r50 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r51 13 30 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.21
+ $Y2=0
r52 13 15 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.99
+ $Y2=0
r53 11 20 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r54 9 30 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=2.21
+ $Y2=0
r55 9 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=1.375
+ $Y2=0
r56 2 33 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.265 $X2=2.26 $Y2=0.4
r57 1 26 91 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.265 $X2=1.21 $Y2=0.4
.ends

