* File: sky130_fd_sc_hdll__clkinv_1.pex.spice
* Created: Wed Sep  2 08:26:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKINV_1%A 1 3 4 6 9 11 12 13 21
r30 21 22 2.75744 $w=4.37e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.282
+ $X2=0.99 $Y2=1.282
r31 20 21 51.8398 $w=4.37e-07 $l=4.7e-07 $layer=POLY_cond $X=0.495 $Y=1.282
+ $X2=0.965 $Y2=1.282
r32 18 20 28.1259 $w=4.37e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=1.282
+ $X2=0.495 $Y2=1.282
r33 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r34 12 13 14.8857 $w=2.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.205 $Y=0.85
+ $X2=0.205 $Y2=1.16
r35 11 12 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.205 $Y=0.51
+ $X2=0.205 $Y2=0.85
r36 7 22 28.039 $w=1.5e-07 $l=2.87e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.282
r37 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.445
r38 4 21 23.583 $w=1.8e-07 $l=2.88e-07 $layer=POLY_cond $X=0.965 $Y=1.57
+ $X2=0.965 $Y2=1.282
r39 4 6 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=0.965 $Y=1.57
+ $X2=0.965 $Y2=2.065
r40 1 20 23.583 $w=1.8e-07 $l=2.88e-07 $layer=POLY_cond $X=0.495 $Y=1.57
+ $X2=0.495 $Y2=1.282
r41 1 3 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=1.57
+ $X2=0.495 $Y2=2.065
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_1%VPWR 1 2 7 9 11 15 17 21 22 28
r22 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r23 22 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r24 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r25 19 28 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.255 $Y2=2.72
r26 19 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.61 $Y2=2.72
r27 17 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r28 17 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r29 13 28 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=2.635
+ $X2=1.255 $Y2=2.72
r30 13 15 33.1327 $w=2.78e-07 $l=8.05e-07 $layer=LI1_cond $X=1.255 $Y=2.635
+ $X2=1.255 $Y2=1.83
r31 12 25 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r32 11 28 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.255 $Y2=2.72
r33 11 12 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r34 7 25 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r35 7 9 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=1.83
r36 2 15 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.645 $X2=1.2 $Y2=1.83
r37 1 9 300 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.645 $X2=0.26 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_1%Y 1 2 9 11 13 14 28 35
r24 31 32 0.0677026 $w=5.28e-07 $l=3e-09 $layer=LI1_cond $X=0.702 $Y=1.025
+ $X2=0.705 $Y2=1.025
r25 28 31 0.27081 $w=5.28e-07 $l=1.2e-08 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.702 $Y2=1.025
r26 21 32 2.68659 $w=3.8e-07 $l=2.65e-07 $layer=LI1_cond $X=0.705 $Y=1.29
+ $X2=0.705 $Y2=1.025
r27 14 35 2.25675 $w=5.28e-07 $l=1e-07 $layer=LI1_cond $X=1.25 $Y=1.025 $X2=1.15
+ $Y2=1.025
r28 13 25 9.09823 $w=3.78e-07 $l=3e-07 $layer=LI1_cond $X=0.705 $Y=1.53
+ $X2=0.705 $Y2=1.83
r29 13 21 7.27859 $w=3.78e-07 $l=2.4e-07 $layer=LI1_cond $X=0.705 $Y=1.53
+ $X2=0.705 $Y2=1.29
r30 11 35 9.25268 $w=5.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.74 $Y=1.025
+ $X2=1.15 $Y2=1.025
r31 11 32 0.789863 $w=5.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.74 $Y=1.025
+ $X2=0.705 $Y2=1.025
r32 7 31 2.77529 $w=3.75e-07 $l=2.65e-07 $layer=LI1_cond $X=0.702 $Y=0.76
+ $X2=0.702 $Y2=1.025
r33 7 9 9.98784 $w=3.73e-07 $l=3.25e-07 $layer=LI1_cond $X=0.702 $Y=0.76
+ $X2=0.702 $Y2=0.435
r34 2 25 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.645 $X2=0.73 $Y2=1.83
r35 1 9 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.725 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_1%VGND 1 6 8 10 17 18 21
r16 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r17 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r18 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r19 15 21 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.255
+ $Y2=0
r20 15 17 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.61
+ $Y2=0
r21 10 21 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.255
+ $Y2=0
r22 10 12 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.23
+ $Y2=0
r23 8 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r24 8 12 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r25 4 21 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=0.085
+ $X2=1.255 $Y2=0
r26 4 6 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.255 $Y=0.085
+ $X2=1.255 $Y2=0.425
r27 1 6 182 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.425
.ends

