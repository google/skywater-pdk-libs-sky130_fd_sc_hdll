* File: sky130_fd_sc_hdll__ebufn_1.pex.spice
* Created: Thu Aug 27 19:06:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EBUFN_1%A 2 3 5 8 10 11 19
r28 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r29 15 18 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.16
+ $X2=0.495 $Y2=1.16
r30 10 11 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.16
+ $X2=0.22 $Y2=1.53
r31 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r32 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r33 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r34 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r35 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.67 $X2=0.495
+ $Y2=1.77
r36 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r37 1 2 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_1%TE_B 2 3 5 6 8 9 11 13 14 15 16
c51 3 0 1.98005e-19 $X=0.965 $Y=1.77
r52 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.125 $Y=1.16
+ $X2=1.125 $Y2=1.53
r53 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.125
+ $Y=1.16 $X2=1.125 $Y2=1.16
r54 14 20 129.397 $w=3.3e-07 $l=7.4e-07 $layer=POLY_cond $X=1.865 $Y=1.16
+ $X2=1.125 $Y2=1.16
r55 12 20 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.1 $Y=1.16
+ $X2=1.125 $Y2=1.16
r56 12 13 3.18546 $w=3.3e-07 $l=1.18e-07 $layer=POLY_cond $X=1.1 $Y=1.16
+ $X2=0.982 $Y2=1.16
r57 9 14 30.0773 $w=3.3e-07 $l=2.95804e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.865 $Y2=1.16
r58 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.985
r59 6 13 33.332 $w=1.75e-07 $l=1.85257e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=0.982 $Y2=1.16
r60 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=0.675
r61 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.77
+ $X2=0.965 $Y2=2.165
r62 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.67 $X2=0.965
+ $Y2=1.77
r63 1 13 33.332 $w=1.75e-07 $l=1.73292e-07 $layer=POLY_cond $X=0.965 $Y=1.325
+ $X2=0.982 $Y2=1.16
r64 1 2 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.965 $Y=1.325
+ $X2=0.965 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_1%A_211_369# 1 2 9 12 16 19 22 23 29 31
c55 19 0 5.53896e-20 $X=1.682 $Y=1.8
r56 23 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.16
+ $X2=2.58 $Y2=0.995
r57 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.16 $X2=2.58 $Y2=1.16
r58 20 29 2.95888 $w=2.5e-07 $l=2.23e-07 $layer=LI1_cond $X=1.905 $Y=1.2
+ $X2=1.682 $Y2=1.2
r59 20 22 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.905 $Y=1.2
+ $X2=2.58 $Y2=1.2
r60 18 29 3.53812 $w=3.87e-07 $l=1.25e-07 $layer=LI1_cond $X=1.682 $Y=1.325
+ $X2=1.682 $Y2=1.2
r61 18 19 12.3014 $w=4.43e-07 $l=4.75e-07 $layer=LI1_cond $X=1.682 $Y=1.325
+ $X2=1.682 $Y2=1.8
r62 14 29 3.53812 $w=3.87e-07 $l=1.50831e-07 $layer=LI1_cond $X=1.625 $Y=1.075
+ $X2=1.682 $Y2=1.2
r63 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.625 $Y=1.075
+ $X2=1.625 $Y2=0.76
r64 10 19 23.8049 $w=2.03e-07 $l=4.4e-07 $layer=LI1_cond $X=1.242 $Y=1.902
+ $X2=1.682 $Y2=1.902
r65 10 12 11.7504 $w=2.53e-07 $l=2.6e-07 $layer=LI1_cond $X=1.242 $Y=2.005
+ $X2=1.242 $Y2=2.265
r66 9 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.64 $Y=0.56 $X2=2.64
+ $Y2=0.995
r67 2 12 600 $w=1.7e-07 $l=4.87134e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.845 $X2=1.2 $Y2=2.265
r68 1 16 182 $w=1.7e-07 $l=6.56125e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.465 $X2=1.625 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_1%A_27_47# 1 2 7 9 10 12 15 19 22 23 24 26
+ 27 28 30 31 32 40
c104 22 0 1.98005e-19 $X=0.657 $Y=1.785
r105 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=1.16 $X2=3.06 $Y2=1.16
r106 40 42 20.4335 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=3.03 $Y=0.82
+ $X2=3.03 $Y2=1.16
r107 31 40 1.77774 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.915 $Y=0.82
+ $X2=3.03 $Y2=0.82
r108 31 32 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.915 $Y=0.82
+ $X2=2.175 $Y2=0.82
r109 30 32 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=2.067 $Y=0.735
+ $X2=2.175 $Y2=0.82
r110 29 30 14.4725 $w=2.13e-07 $l=2.7e-07 $layer=LI1_cond $X=2.067 $Y=0.465
+ $X2=2.067 $Y2=0.735
r111 27 29 6.81772 $w=2.1e-07 $l=1.50612e-07 $layer=LI1_cond $X=1.96 $Y=0.36
+ $X2=2.067 $Y2=0.465
r112 27 28 38.29 $w=2.08e-07 $l=7.25e-07 $layer=LI1_cond $X=1.96 $Y=0.36
+ $X2=1.235 $Y2=0.36
r113 25 28 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.15 $Y=0.465
+ $X2=1.235 $Y2=0.36
r114 25 26 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.15 $Y=0.465
+ $X2=1.15 $Y2=0.615
r115 23 26 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.065 $Y=0.72
+ $X2=1.15 $Y2=0.615
r116 23 24 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.065 $Y=0.72
+ $X2=0.79 $Y2=0.72
r117 21 24 7.02424 $w=2.08e-07 $l=1.33e-07 $layer=LI1_cond $X=0.657 $Y=0.72
+ $X2=0.79 $Y2=0.72
r118 21 22 41.7489 $w=2.63e-07 $l=9.6e-07 $layer=LI1_cond $X=0.657 $Y=0.825
+ $X2=0.657 $Y2=1.785
r119 17 22 23.1536 $w=2.18e-07 $l=4.42e-07 $layer=LI1_cond $X=0.215 $Y=1.895
+ $X2=0.657 $Y2=1.895
r120 17 19 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.215 $Y=2.005
+ $X2=0.215 $Y2=2.22
r121 13 21 23.3437 $w=2.08e-07 $l=4.42e-07 $layer=LI1_cond $X=0.215 $Y=0.72
+ $X2=0.657 $Y2=0.72
r122 13 15 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.215 $Y=0.615
+ $X2=0.215 $Y2=0.445
r123 10 43 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.025 $Y=1.41
+ $X2=3.06 $Y2=1.16
r124 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.025 $Y=1.41
+ $X2=3.025 $Y2=1.985
r125 7 43 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3 $Y=0.995
+ $X2=3.06 $Y2=1.16
r126 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3 $Y=0.995 $X2=3
+ $Y2=0.56
r127 2 19 600 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.22
r128 1 15 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_1%VPWR 1 2 9 11 15 17 19 29 30 33 36
c45 29 0 5.53896e-20 $X=3.45 $Y=2.72
r46 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r47 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r49 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r50 27 30 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r51 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 26 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 24 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.9 $Y=2.72 $X2=1.72
+ $Y2=2.72
r55 24 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.9 $Y=2.72 $X2=2.07
+ $Y2=2.72
r56 19 33 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.702 $Y2=2.72
r57 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 17 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r60 13 36 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.72
r61 13 15 12.0046 $w=3.58e-07 $l=3.75e-07 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.26
r62 12 33 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.89 $Y=2.72
+ $X2=0.702 $Y2=2.72
r63 11 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.54 $Y=2.72 $X2=1.72
+ $Y2=2.72
r64 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.54 $Y=2.72
+ $X2=0.89 $Y2=2.72
r65 7 33 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.702 $Y=2.635
+ $X2=0.702 $Y2=2.72
r66 7 9 8.45125 $w=3.73e-07 $l=2.75e-07 $layer=LI1_cond $X=0.702 $Y=2.635
+ $X2=0.702 $Y2=2.36
r67 2 15 600 $w=1.7e-07 $l=8.35165e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.485 $X2=1.72 $Y2=2.26
r68 1 9 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.845 $X2=0.73 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_1%Z 1 2 7 9 11 13 14 15 16 33 37 44 48 53 55
r27 55 61 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.45 $Y=0.85
+ $X2=3.45 $Y2=0.825
r28 33 44 2.26392 $w=9.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.315 $Y=1.98
+ $X2=3.135 $Y2=1.98
r29 16 53 7.9237 $w=2.7e-07 $l=4.85e-07 $layer=LI1_cond $X=3.45 $Y=1.98 $X2=3.45
+ $Y2=1.495
r30 16 33 2.20557 $w=9.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.45 $Y=1.98
+ $X2=3.315 $Y2=1.98
r31 16 53 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.45 $Y=1.47
+ $X2=3.45 $Y2=1.495
r32 15 16 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.45 $Y=1.19
+ $X2=3.45 $Y2=1.47
r33 14 61 1.46269 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=3.42 $Y=0.795 $X2=3.42
+ $Y2=0.825
r34 14 46 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.42 $Y=0.795
+ $X2=3.42 $Y2=0.66
r35 14 15 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.45 $Y=0.88
+ $X2=3.45 $Y2=1.19
r36 14 55 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=3.45 $Y=0.88 $X2=3.45
+ $Y2=0.85
r37 13 46 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.42 $Y=0.51
+ $X2=3.42 $Y2=0.66
r38 13 48 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.42 $Y=0.51
+ $X2=3.42 $Y2=0.4
r39 11 44 0.125773 $w=9.68e-07 $l=1e-08 $layer=LI1_cond $X=3.125 $Y=1.98
+ $X2=3.135 $Y2=1.98
r40 9 11 5.53402 $w=9.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.685 $Y=1.98
+ $X2=3.125 $Y2=1.98
r41 9 37 5.53402 $w=9.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.685 $Y=1.98
+ $X2=2.245 $Y2=1.98
r42 7 37 0.251546 $w=9.68e-07 $l=2e-08 $layer=LI1_cond $X=2.225 $Y=1.98
+ $X2=2.245 $Y2=1.98
r43 2 16 300 $w=1.7e-07 $l=4.44972e-07 $layer=licon1_PDIFF $count=2 $X=3.115
+ $Y=1.485 $X2=3.385 $Y2=1.815
r44 1 48 91 $w=1.7e-07 $l=4.19464e-07 $layer=licon1_NDIFF $count=2 $X=3.075
+ $Y=0.235 $X2=3.42 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_1%VGND 1 2 7 9 24 25 29 36 43
r43 41 43 9.19385 $w=6.48e-07 $l=9.5e-08 $layer=LI1_cond $X=2.99 $Y=0.24
+ $X2=3.085 $Y2=0.24
r44 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r45 39 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r46 38 41 8.46455 $w=6.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=0.24
+ $X2=2.99 $Y2=0.24
r47 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r48 35 38 1.84012 $w=6.48e-07 $l=1e-07 $layer=LI1_cond $X=2.43 $Y=0.24 $X2=2.53
+ $Y2=0.24
r49 35 36 9.00983 $w=6.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=0.24
+ $X2=2.345 $Y2=0.24
r50 29 32 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.705
+ $Y2=0.36
r51 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r52 25 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r53 24 43 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.085
+ $Y2=0
r54 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r55 21 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r56 20 36 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.345
+ $Y2=0
r57 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r58 18 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r59 18 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r60 17 20 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r61 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r62 15 29 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r63 15 17 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r64 9 29 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r65 9 11 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r66 7 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r67 7 11 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r68 2 35 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.235 $X2=2.43 $Y2=0.38
r69 1 32 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.36
.ends

