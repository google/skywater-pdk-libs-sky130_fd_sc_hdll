* File: sky130_fd_sc_hdll__nand2b_4.pex.spice
* Created: Wed Sep  2 08:37:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2B_4%A_N 1 3 6 8 13
c31 8 0 1.24063e-19 $X=0.235 $Y=1.19
r32 13 14 3.61862 $w=3.33e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.212
+ $X2=0.52 $Y2=1.212
r33 11 13 31.8438 $w=3.33e-07 $l=2.2e-07 $layer=POLY_cond $X=0.275 $Y=1.212
+ $X2=0.495 $Y2=1.212
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r35 4 14 21.4384 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=1.212
r36 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=0.56
r37 1 13 17.1428 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.212
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_4%A_27_47# 1 2 7 9 12 14 16 19 21 23 26 28
+ 30 33 37 39 41 43 44 45 48 50 56 61 62 72
c128 62 0 1.24063e-19 $X=1.385 $Y=1.16
r129 72 73 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.895 $Y=1.217
+ $X2=2.92 $Y2=1.217
r130 71 72 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=2.45 $Y=1.217
+ $X2=2.895 $Y2=1.217
r131 70 71 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.425 $Y=1.217
+ $X2=2.45 $Y2=1.217
r132 67 68 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.955 $Y=1.217
+ $X2=1.98 $Y2=1.217
r133 66 67 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=1.51 $Y=1.217
+ $X2=1.955 $Y2=1.217
r134 65 66 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.217
+ $X2=1.51 $Y2=1.217
r135 62 65 16.3472 $w=3.27e-07 $l=1.253e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.485 $Y2=1.217
r136 57 70 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=2.19 $Y=1.217
+ $X2=2.425 $Y2=1.217
r137 57 68 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=2.19 $Y=1.217
+ $X2=1.98 $Y2=1.217
r138 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.16 $X2=2.19 $Y2=1.16
r139 54 62 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.16
+ $X2=1.385 $Y2=1.16
r140 53 56 53.7909 $w=1.98e-07 $l=9.7e-07 $layer=LI1_cond $X=1.22 $Y=1.175
+ $X2=2.19 $Y2=1.175
r141 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.16 $X2=1.22 $Y2=1.16
r142 51 61 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=1.175
+ $X2=0.745 $Y2=1.175
r143 51 53 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=0.83 $Y=1.175
+ $X2=1.22 $Y2=1.175
r144 49 61 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.745 $Y=1.275
+ $X2=0.745 $Y2=1.175
r145 49 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.745 $Y=1.275
+ $X2=0.745 $Y2=1.445
r146 48 61 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.745 $Y=1.075
+ $X2=0.745 $Y2=1.175
r147 47 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.745 $Y=0.905
+ $X2=0.745 $Y2=1.075
r148 46 60 4.35361 $w=2.2e-07 $l=1.68e-07 $layer=LI1_cond $X=0.425 $Y=1.555
+ $X2=0.257 $Y2=1.555
r149 45 50 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.66 $Y=1.555
+ $X2=0.745 $Y2=1.445
r150 45 46 12.3102 $w=2.18e-07 $l=2.35e-07 $layer=LI1_cond $X=0.66 $Y=1.555
+ $X2=0.425 $Y2=1.555
r151 43 47 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.66 $Y=0.81
+ $X2=0.745 $Y2=0.905
r152 43 44 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=0.66 $Y=0.81
+ $X2=0.425 $Y2=0.81
r153 39 60 2.85058 $w=3.35e-07 $l=1.1e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=1.555
r154 39 41 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=2.34
r155 35 44 7.51555 $w=1.9e-07 $l=2.102e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.425 $Y2=0.81
r156 35 37 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.257 $Y2=0.38
r157 31 73 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.92 $Y=1.025
+ $X2=2.92 $Y2=1.217
r158 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.92 $Y=1.025
+ $X2=2.92 $Y2=0.56
r159 28 72 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.217
r160 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
r161 24 71 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=1.217
r162 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=0.56
r163 21 70 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.217
r164 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
r165 17 68 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.98 $Y=1.025
+ $X2=1.98 $Y2=1.217
r166 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.98 $Y=1.025
+ $X2=1.98 $Y2=0.56
r167 14 67 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.217
r168 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r169 10 66 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.51 $Y=1.025
+ $X2=1.51 $Y2=1.217
r170 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.51 $Y=1.025
+ $X2=1.51 $Y2=0.56
r171 7 65 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.217
r172 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r173 2 60 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r174 2 41 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r175 1 37 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_4%B 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 32 37 39 54 61 63 65 69
c86 5 0 1.59283e-19 $X=3.38 $Y=1.41
r87 63 65 0.0554545 $w=1.98e-07 $l=1e-09 $layer=LI1_cond $X=4.744 $Y=1.175
+ $X2=4.745 $Y2=1.175
r88 61 63 20.1855 $w=1.98e-07 $l=3.64e-07 $layer=LI1_cond $X=4.38 $Y=1.175
+ $X2=4.744 $Y2=1.175
r89 51 52 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.79 $Y=1.217
+ $X2=4.815 $Y2=1.217
r90 50 51 69.2783 $w=3.27e-07 $l=4.7e-07 $layer=POLY_cond $X=4.32 $Y=1.217
+ $X2=4.79 $Y2=1.217
r91 49 50 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.295 $Y=1.217
+ $X2=4.32 $Y2=1.217
r92 48 49 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=3.85 $Y=1.217
+ $X2=4.295 $Y2=1.217
r93 47 48 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.825 $Y=1.217
+ $X2=3.85 $Y2=1.217
r94 46 54 8.04091 $w=1.98e-07 $l=1.45e-07 $layer=LI1_cond $X=3.62 $Y=1.175
+ $X2=3.475 $Y2=1.175
r95 45 47 30.2171 $w=3.27e-07 $l=2.05e-07 $layer=POLY_cond $X=3.62 $Y=1.217
+ $X2=3.825 $Y2=1.217
r96 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.62
+ $Y=1.16 $X2=3.62 $Y2=1.16
r97 43 45 35.3761 $w=3.27e-07 $l=2.4e-07 $layer=POLY_cond $X=3.38 $Y=1.217
+ $X2=3.62 $Y2=1.217
r98 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.355 $Y=1.217
+ $X2=3.38 $Y2=1.217
r99 40 69 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=5.055 $Y=1.175
+ $X2=5.19 $Y2=1.175
r100 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.055
+ $Y=1.16 $X2=5.055 $Y2=1.16
r101 37 52 12.6622 $w=3.27e-07 $l=9.94987e-08 $layer=POLY_cond $X=4.89 $Y=1.16
+ $X2=4.815 $Y2=1.217
r102 37 39 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.16
+ $X2=5.055 $Y2=1.16
r103 32 69 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=5.305 $Y=1.175
+ $X2=5.19 $Y2=1.175
r104 31 40 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=4.83 $Y=1.175
+ $X2=5.055 $Y2=1.175
r105 31 65 4.71364 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=4.83 $Y=1.175
+ $X2=4.745 $Y2=1.175
r106 30 61 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=4.375 $Y=1.175
+ $X2=4.38 $Y2=1.175
r107 29 30 25.7864 $w=1.98e-07 $l=4.65e-07 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=4.375 $Y2=1.175
r108 29 46 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=3.62 $Y2=1.175
r109 25 52 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.815 $Y=1.025
+ $X2=4.815 $Y2=1.217
r110 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.815 $Y=1.025
+ $X2=4.815 $Y2=0.56
r111 22 51 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.79 $Y=1.41
+ $X2=4.79 $Y2=1.217
r112 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.79 $Y=1.41
+ $X2=4.79 $Y2=1.985
r113 19 50 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.32 $Y=1.41
+ $X2=4.32 $Y2=1.217
r114 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.32 $Y=1.41
+ $X2=4.32 $Y2=1.985
r115 15 49 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.295 $Y=1.025
+ $X2=4.295 $Y2=1.217
r116 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.295 $Y=1.025
+ $X2=4.295 $Y2=0.56
r117 12 48 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.85 $Y=1.41
+ $X2=3.85 $Y2=1.217
r118 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.85 $Y=1.41
+ $X2=3.85 $Y2=1.985
r119 8 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.825 $Y=1.025
+ $X2=3.825 $Y2=1.217
r120 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.825 $Y=1.025
+ $X2=3.825 $Y2=0.56
r121 5 43 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.217
r122 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.985
r123 1 42 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.355 $Y=1.025
+ $X2=3.355 $Y2=1.217
r124 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.355 $Y=1.025
+ $X2=3.355 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_4%VPWR 1 2 3 4 5 6 24 27 31 35 39 41 43 48
+ 51 52 54 55 57 58 59 71 76 82
r87 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r88 77 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 76 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r91 74 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r92 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r93 71 81 4.54404 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=4.97 $Y=2.72
+ $X2=5.245 $Y2=2.72
r94 71 73 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.97 $Y=2.72
+ $X2=4.83 $Y2=2.72
r95 70 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r96 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r97 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r98 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r99 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r100 64 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r101 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r102 61 76 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=0.99 $Y2=2.72
r103 61 63 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r104 59 79 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r105 57 69 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4 $Y=2.72 $X2=3.91
+ $Y2=2.72
r106 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4 $Y=2.72 $X2=4.085
+ $Y2=2.72
r107 56 73 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.17 $Y=2.72
+ $X2=4.83 $Y2=2.72
r108 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=2.72
+ $X2=4.085 $Y2=2.72
r109 54 66 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.06 $Y=2.72 $X2=2.99
+ $Y2=2.72
r110 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=2.72
+ $X2=3.145 $Y2=2.72
r111 53 69 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.23 $Y=2.72
+ $X2=3.91 $Y2=2.72
r112 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=2.72
+ $X2=3.145 $Y2=2.72
r113 51 63 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r114 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.19 $Y2=2.72
r115 50 66 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.99 $Y2=2.72
r116 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.19 $Y2=2.72
r117 48 49 6.43014 $w=6.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=2 $X2=0.99
+ $Y2=1.835
r118 43 46 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.135 $Y=1.66
+ $X2=5.135 $Y2=2.34
r119 41 81 3.22214 $w=3.3e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.135 $Y=2.635
+ $X2=5.245 $Y2=2.72
r120 41 46 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.135 $Y=2.635
+ $X2=5.135 $Y2=2.34
r121 37 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=2.635
+ $X2=4.085 $Y2=2.72
r122 37 39 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.085 $Y=2.635
+ $X2=4.085 $Y2=2
r123 33 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=2.635
+ $X2=3.145 $Y2=2.72
r124 33 35 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.145 $Y=2.635
+ $X2=3.145 $Y2=2
r125 29 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r126 29 31 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2
r127 27 49 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=1.177 $Y=1.66
+ $X2=1.177 $Y2=1.835
r128 22 76 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=2.635
+ $X2=0.99 $Y2=2.72
r129 22 24 5.11367 $w=6.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.99 $Y=2.635
+ $X2=0.99 $Y2=2.34
r130 21 48 3.1202 $w=6.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.99 $Y=2.18
+ $X2=0.99 $Y2=2
r131 21 24 2.77352 $w=6.88e-07 $l=1.6e-07 $layer=LI1_cond $X=0.99 $Y=2.18
+ $X2=0.99 $Y2=2.34
r132 6 46 400 $w=1.7e-07 $l=9.74192e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.485 $X2=5.135 $Y2=2.34
r133 6 43 400 $w=1.7e-07 $l=3.31134e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.485 $X2=5.135 $Y2=1.66
r134 5 39 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.94
+ $Y=1.485 $X2=4.085 $Y2=2
r135 4 35 300 $w=1.7e-07 $l=5.89597e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.485 $X2=3.145 $Y2=2
r136 3 31 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2
r137 2 27 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=1.66
r138 2 24 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=2.34
r139 1 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_4%Y 1 2 3 4 5 6 19 23 25 27 29 30 31 35 37
+ 39 41 48 51 52 53
c104 48 0 1.4834e-19 $X=3.615 $Y=1.66
c105 30 0 1.59283e-19 $X=2.707 $Y=1.445
c106 29 0 1.21227e-19 $X=2.707 $Y=0.905
r107 53 65 3.35521 $w=3.93e-07 $l=1.15e-07 $layer=LI1_cond $X=2.642 $Y=2.225
+ $X2=2.642 $Y2=2.34
r108 52 53 9.91976 $w=3.93e-07 $l=3.4e-07 $layer=LI1_cond $X=2.642 $Y=1.885
+ $X2=2.642 $Y2=2.225
r109 52 57 6.41867 $w=3.93e-07 $l=2.2e-07 $layer=LI1_cond $X=2.642 $Y=1.885
+ $X2=2.642 $Y2=1.665
r110 51 57 1.91251 $w=3.95e-07 $l=1.1e-07 $layer=LI1_cond $X=2.642 $Y=1.555
+ $X2=2.642 $Y2=1.665
r111 39 50 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=4.53 $Y=1.665
+ $X2=4.53 $Y2=1.555
r112 39 41 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.53 $Y=1.665
+ $X2=4.53 $Y2=2.34
r113 38 48 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.78 $Y=1.555
+ $X2=3.59 $Y2=1.555
r114 37 50 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.34 $Y=1.555
+ $X2=4.53 $Y2=1.555
r115 37 38 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=4.34 $Y=1.555
+ $X2=3.78 $Y2=1.555
r116 33 48 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=3.59 $Y=1.665
+ $X2=3.59 $Y2=1.555
r117 33 35 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.59 $Y=1.665
+ $X2=3.59 $Y2=2.34
r118 32 51 4.36787 $w=2.2e-07 $l=1.98e-07 $layer=LI1_cond $X=2.84 $Y=1.555
+ $X2=2.642 $Y2=1.555
r119 31 48 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.4 $Y=1.555
+ $X2=3.59 $Y2=1.555
r120 31 32 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=3.4 $Y=1.555
+ $X2=2.84 $Y2=1.555
r121 30 51 1.91251 $w=2.65e-07 $l=1.38744e-07 $layer=LI1_cond $X=2.707 $Y=1.445
+ $X2=2.642 $Y2=1.555
r122 29 46 3.44693 $w=2.65e-07 $l=1.35e-07 $layer=LI1_cond $X=2.707 $Y=0.905
+ $X2=2.707 $Y2=0.77
r123 29 30 23.4837 $w=2.63e-07 $l=5.4e-07 $layer=LI1_cond $X=2.707 $Y=0.905
+ $X2=2.707 $Y2=1.445
r124 28 44 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.885 $Y=1.555
+ $X2=1.695 $Y2=1.555
r125 27 51 4.36787 $w=2.2e-07 $l=1.97e-07 $layer=LI1_cond $X=2.445 $Y=1.555
+ $X2=2.642 $Y2=1.555
r126 27 28 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=2.445 $Y=1.555
+ $X2=1.885 $Y2=1.555
r127 23 44 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.555
r128 23 25 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=2.34
r129 19 46 3.37033 $w=2.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.575 $Y=0.77
+ $X2=2.707 $Y2=0.77
r130 19 21 36.494 $w=2.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.575 $Y=0.77
+ $X2=1.72 $Y2=0.77
r131 6 50 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.485 $X2=4.555 $Y2=1.66
r132 6 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.485 $X2=4.555 $Y2=2.34
r133 5 48 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.485 $X2=3.615 $Y2=1.66
r134 5 35 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.485 $X2=3.615 $Y2=2.34
r135 4 51 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=1.66
r136 4 65 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=2.34
r137 3 44 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=1.66
r138 3 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=2.34
r139 2 46 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.235 $X2=2.66 $Y2=0.72
r140 1 21 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.72 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_4%VGND 1 2 3 14 18 22 25 26 28 29 30 43 44
+ 47 50
r74 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r75 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r76 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r77 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r78 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r79 37 38 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r80 35 38 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r81 35 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r82 34 37 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r83 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r84 32 47 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=0.84 $Y=0 $X2=0.742
+ $Y2=0
r85 32 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.84 $Y=0 $X2=1.15
+ $Y2=0
r86 30 48 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r87 30 50 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r88 28 40 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.37
+ $Y2=0
r89 28 29 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.59
+ $Y2=0
r90 27 43 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.71 $Y=0 $X2=5.29
+ $Y2=0
r91 27 29 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.71 $Y=0 $X2=4.59
+ $Y2=0
r92 25 37 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.53 $Y=0 $X2=3.45
+ $Y2=0
r93 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=0 $X2=3.615
+ $Y2=0
r94 24 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=4.37
+ $Y2=0
r95 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.615
+ $Y2=0
r96 20 29 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0
r97 20 22 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0.38
r98 16 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=0.085
+ $X2=3.615 $Y2=0
r99 16 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.615 $Y=0.085
+ $X2=3.615 $Y2=0.38
r100 12 47 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.742 $Y=0.085
+ $X2=0.742 $Y2=0
r101 12 14 16.7786 $w=1.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.742 $Y=0.085
+ $X2=0.742 $Y2=0.38
r102 3 22 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=4.37
+ $Y=0.235 $X2=4.555 $Y2=0.38
r103 2 18 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.235 $X2=3.615 $Y2=0.38
r104 1 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2B_4%A_225_47# 1 2 3 4 5 16 18 20 24 25 26 30
+ 32 36 44
c80 26 0 1.4834e-19 $X=3.87 $Y=0.81
r81 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.135 $Y=0.715
+ $X2=5.135 $Y2=0.38
r82 33 44 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.25 $Y=0.81 $X2=4.06
+ $Y2=0.81
r83 32 34 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=4.97 $Y=0.81
+ $X2=5.135 $Y2=0.715
r84 32 33 42.0287 $w=1.88e-07 $l=7.2e-07 $layer=LI1_cond $X=4.97 $Y=0.81
+ $X2=4.25 $Y2=0.81
r85 28 44 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.06 $Y=0.715
+ $X2=4.06 $Y2=0.81
r86 28 30 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.06 $Y=0.715
+ $X2=4.06 $Y2=0.38
r87 27 43 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.31 $Y=0.81
+ $X2=3.185 $Y2=0.81
r88 26 44 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.87 $Y=0.81 $X2=4.06
+ $Y2=0.81
r89 26 27 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=3.87 $Y=0.81 $X2=3.31
+ $Y2=0.81
r90 25 43 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=3.185 $Y=0.715
+ $X2=3.185 $Y2=0.81
r91 24 41 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.185 $Y=0.465
+ $X2=3.185 $Y2=0.36
r92 24 25 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=3.185 $Y=0.465
+ $X2=3.185 $Y2=0.715
r93 21 39 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.335 $Y=0.36
+ $X2=1.21 $Y2=0.36
r94 21 23 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=1.335 $Y=0.36
+ $X2=2.19 $Y2=0.36
r95 20 41 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.06 $Y=0.36
+ $X2=3.185 $Y2=0.36
r96 20 23 45.9481 $w=2.08e-07 $l=8.7e-07 $layer=LI1_cond $X=3.06 $Y=0.36
+ $X2=2.19 $Y2=0.36
r97 16 39 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.21 $Y=0.465
+ $X2=1.21 $Y2=0.36
r98 16 18 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.21 $Y=0.465
+ $X2=1.21 $Y2=0.72
r99 5 36 91 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=2 $X=4.89
+ $Y=0.235 $X2=5.135 $Y2=0.38
r100 4 30 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.9
+ $Y=0.235 $X2=4.085 $Y2=0.38
r101 3 43 182 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.235 $X2=3.145 $Y2=0.72
r102 3 41 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.235 $X2=3.145 $Y2=0.38
r103 2 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.38
r104 1 39 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.38
r105 1 18 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.72
.ends

