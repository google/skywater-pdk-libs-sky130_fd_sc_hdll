* File: sky130_fd_sc_hdll__nor2_1.pex.spice
* Created: Wed Sep  2 08:39:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR2_1%B 1 3 4 6 7
r25 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r26 4 10 40.1292 $w=4.26e-07 $l=2.36525e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.352 $Y2=1.16
r27 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r28 1 10 44.7281 $w=4.26e-07 $l=3.13449e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.352 $Y2=1.16
r29 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_1%A 1 3 4 6 7 10
r26 10 12 32.5317 $w=3.63e-07 $l=2.45e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.21 $Y2=1.202
r27 9 10 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r28 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.16 $X2=1.21 $Y2=1.16
r29 4 10 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r30 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r31 1 9 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_1%Y 1 2 7 11 14 15 18 19
c32 14 0 1.00411e-19 $X=0.69 $Y=1.495
r33 19 24 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=2.21
+ $X2=0.26 $Y2=2.34
r34 15 19 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.21
r35 15 17 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.665 $X2=0.26
+ $Y2=1.58
r36 14 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.69 $Y=1.495 $X2=0.69
+ $Y2=0.895
r37 9 18 7.683 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=0.705 $Y=0.705
+ $X2=0.705 $Y2=0.895
r38 9 11 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=0.705
+ $X2=0.705 $Y2=0.39
r39 8 17 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=1.58
+ $X2=0.26 $Y2=1.58
r40 7 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=1.58
+ $X2=0.69 $Y2=1.495
r41 7 8 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.605 $Y=1.58
+ $X2=0.425 $Y2=1.58
r42 2 24 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r43 2 17 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r44 1 11 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_1%VPWR 1 4 6 10 12 19
r18 19 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r19 18 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r20 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r21 12 18 6.08638 $w=1.7e-07 $l=3.62e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.477 $Y2=2.72
r22 12 14 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.23 $Y2=2.72
r23 10 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r24 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r25 6 9 15.9477 $w=5.08e-07 $l=6.8e-07 $layer=LI1_cond $X=1.37 $Y=1.66 $X2=1.37
+ $Y2=2.34
r26 4 18 3.22813 $w=5.1e-07 $l=1.43332e-07 $layer=LI1_cond $X=1.37 $Y=2.635
+ $X2=1.477 $Y2=2.72
r27 4 9 6.91849 $w=5.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.37 $Y=2.635
+ $X2=1.37 $Y2=2.34
r28 1 9 200 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=3 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r29 1 6 200 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=3 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_1%VGND 1 2 7 9 11 13 15 17 27
r22 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r23 21 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r24 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r25 18 23 3.93736 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r26 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r27 17 26 5.96807 $w=1.7e-07 $l=3.87e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.452
+ $Y2=0
r28 17 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.69
+ $Y2=0
r29 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r30 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r31 11 26 3.34644 $w=5.1e-07 $l=1.69245e-07 $layer=LI1_cond $X=1.32 $Y=0.085
+ $X2=1.452 $Y2=0
r32 11 13 7.15302 $w=5.08e-07 $l=3.05e-07 $layer=LI1_cond $X=1.32 $Y=0.085
+ $X2=1.32 $Y2=0.39
r33 7 23 3.14078 $w=2.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.172 $Y2=0
r34 7 9 14.6456 $w=2.38e-07 $l=3.05e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.39
r35 2 13 45.5 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_NDIFF $count=4 $X=1.015
+ $Y=0.235 $X2=1.49 $Y2=0.39
r36 1 9 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

