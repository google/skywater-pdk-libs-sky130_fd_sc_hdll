* File: sky130_fd_sc_hdll__a21boi_4.pxi.spice
* Created: Thu Aug 27 18:52:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21BOI_4%B1_N N_B1_N_c_91_n N_B1_N_M1010_g N_B1_N_c_92_n
+ N_B1_N_M1015_g B1_N PM_SKY130_FD_SC_HDLL__A21BOI_4%B1_N
x_PM_SKY130_FD_SC_HDLL__A21BOI_4%A_27_47# N_A_27_47#_M1015_s N_A_27_47#_M1010_s
+ N_A_27_47#_c_123_n N_A_27_47#_M1002_g N_A_27_47#_c_132_n N_A_27_47#_M1005_g
+ N_A_27_47#_c_124_n N_A_27_47#_M1018_g N_A_27_47#_c_133_n N_A_27_47#_M1008_g
+ N_A_27_47#_c_125_n N_A_27_47#_M1019_g N_A_27_47#_c_134_n N_A_27_47#_M1016_g
+ N_A_27_47#_c_126_n N_A_27_47#_M1025_g N_A_27_47#_c_135_n N_A_27_47#_M1022_g
+ N_A_27_47#_c_127_n N_A_27_47#_c_128_n N_A_27_47#_c_136_n N_A_27_47#_c_149_n
+ N_A_27_47#_c_129_n N_A_27_47#_c_137_n N_A_27_47#_c_138_n N_A_27_47#_c_139_n
+ N_A_27_47#_c_130_n N_A_27_47#_c_131_n PM_SKY130_FD_SC_HDLL__A21BOI_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__A21BOI_4%A2 N_A2_c_241_n N_A2_M1003_g N_A2_c_242_n
+ N_A2_M1000_g N_A2_c_243_n N_A2_M1001_g N_A2_c_251_n N_A2_M1006_g N_A2_c_252_n
+ N_A2_M1011_g N_A2_c_244_n N_A2_M1004_g N_A2_c_253_n N_A2_M1023_g N_A2_c_245_n
+ N_A2_M1012_g N_A2_c_246_n N_A2_c_263_n N_A2_c_247_n N_A2_c_256_n A2
+ N_A2_c_248_n N_A2_c_249_n A2 PM_SKY130_FD_SC_HDLL__A21BOI_4%A2
x_PM_SKY130_FD_SC_HDLL__A21BOI_4%A1 N_A1_c_366_n N_A1_M1007_g N_A1_c_372_n
+ N_A1_M1014_g N_A1_c_373_n N_A1_M1017_g N_A1_c_367_n N_A1_M1009_g N_A1_c_374_n
+ N_A1_M1021_g N_A1_c_368_n N_A1_M1013_g N_A1_c_375_n N_A1_M1024_g N_A1_c_369_n
+ N_A1_M1020_g A1 N_A1_c_370_n N_A1_c_371_n A1 PM_SKY130_FD_SC_HDLL__A21BOI_4%A1
x_PM_SKY130_FD_SC_HDLL__A21BOI_4%VPWR N_VPWR_M1010_d N_VPWR_M1003_d
+ N_VPWR_M1017_d N_VPWR_M1024_d N_VPWR_M1011_d N_VPWR_c_440_n N_VPWR_c_441_n
+ N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n VPWR N_VPWR_c_445_n
+ N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_439_n N_VPWR_c_449_n N_VPWR_c_450_n
+ N_VPWR_c_451_n PM_SKY130_FD_SC_HDLL__A21BOI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A21BOI_4%A_227_297# N_A_227_297#_M1005_d
+ N_A_227_297#_M1008_d N_A_227_297#_M1022_d N_A_227_297#_M1014_s
+ N_A_227_297#_M1021_s N_A_227_297#_M1006_s N_A_227_297#_M1023_s
+ N_A_227_297#_c_597_n N_A_227_297#_c_556_n N_A_227_297#_c_560_n
+ N_A_227_297#_c_570_n N_A_227_297#_c_562_n N_A_227_297#_c_613_n
+ N_A_227_297#_c_575_n N_A_227_297#_c_620_n N_A_227_297#_c_577_n
+ N_A_227_297#_c_554_n N_A_227_297#_c_555_n N_A_227_297#_c_583_n
+ N_A_227_297#_c_584_n PM_SKY130_FD_SC_HDLL__A21BOI_4%A_227_297#
x_PM_SKY130_FD_SC_HDLL__A21BOI_4%Y N_Y_M1002_s N_Y_M1019_s N_Y_M1007_d
+ N_Y_M1013_d N_Y_M1005_s N_Y_M1016_s N_Y_c_641_n N_Y_c_699_p N_Y_c_645_n
+ N_Y_c_636_n N_Y_c_637_n N_Y_c_638_n N_Y_c_653_n N_Y_c_658_n N_Y_c_660_n
+ N_Y_c_661_n N_Y_c_639_n Y Y PM_SKY130_FD_SC_HDLL__A21BOI_4%Y
x_PM_SKY130_FD_SC_HDLL__A21BOI_4%VGND N_VGND_M1015_d N_VGND_M1018_d
+ N_VGND_M1025_d N_VGND_M1001_s N_VGND_M1012_s N_VGND_c_724_n N_VGND_c_725_n
+ N_VGND_c_726_n N_VGND_c_727_n N_VGND_c_728_n N_VGND_c_729_n VGND
+ N_VGND_c_730_n N_VGND_c_731_n N_VGND_c_732_n N_VGND_c_733_n N_VGND_c_734_n
+ N_VGND_c_735_n PM_SKY130_FD_SC_HDLL__A21BOI_4%VGND
x_PM_SKY130_FD_SC_HDLL__A21BOI_4%A_724_47# N_A_724_47#_M1000_d
+ N_A_724_47#_M1009_s N_A_724_47#_M1020_s N_A_724_47#_M1004_d
+ N_A_724_47#_c_829_n N_A_724_47#_c_830_n N_A_724_47#_c_831_n
+ N_A_724_47#_c_827_n N_A_724_47#_c_828_n N_A_724_47#_c_842_n
+ PM_SKY130_FD_SC_HDLL__A21BOI_4%A_724_47#
cc_1 VNB N_B1_N_c_91_n 0.0348363f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_2 VNB N_B1_N_c_92_n 0.0231164f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=0.995
cc_3 VNB B1_N 0.0147405f $X=-0.19 $Y=-0.24 $X2=0.175 $Y2=1.445
cc_4 VNB N_A_27_47#_c_123_n 0.016884f $X=-0.19 $Y=-0.24 $X2=0.175 $Y2=1.445
cc_5 VNB N_A_27_47#_c_124_n 0.0171475f $X=-0.19 $Y=-0.24 $X2=0.392 $Y2=1.53
cc_6 VNB N_A_27_47#_c_125_n 0.0166697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_126_n 0.0197746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_127_n 0.0088069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_128_n 0.0144029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_129_n 0.00160741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_130_n 0.00260583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_131_n 0.0940855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_241_n 0.0267652f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_14 VNB N_A2_c_242_n 0.0197241f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=0.995
cc_15 VNB N_A2_c_243_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0.175 $Y2=1.445
cc_16 VNB N_A2_c_244_n 0.0172939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A2_c_245_n 0.0224545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_246_n 0.00160282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_247_n 0.00239395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_248_n 0.0706013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A2_c_249_n 0.00961897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A1_c_366_n 0.0166783f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_23 VNB N_A1_c_367_n 0.0170186f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.16
cc_24 VNB N_A1_c_368_n 0.0169333f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A1_c_369_n 0.016668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A1_c_370_n 0.00170867f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A1_c_371_n 0.100169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_439_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_636_n 0.00434246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_637_n 2.63992e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_638_n 0.0110398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_639_n 0.00691285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_724_n 0.00479809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_725_n 0.0106437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_726_n 0.0344016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_727_n 0.0311056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_728_n 0.0619488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_729_n 0.00362451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_730_n 0.0165531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_731_n 0.0185827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_732_n 0.00796566f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_733_n 0.0139287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_734_n 0.019048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_735_n 0.353209f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_724_47#_c_827_n 0.00534476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_724_47#_c_828_n 0.00280167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VPB N_B1_N_c_91_n 0.0365574f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_48 VPB B1_N 0.014796f $X=-0.19 $Y=1.305 $X2=0.175 $Y2=1.445
cc_49 VPB N_A_27_47#_c_132_n 0.0196741f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.16
cc_50 VPB N_A_27_47#_c_133_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_134_n 0.0164114f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_135_n 0.0159808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_136_n 0.00467003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_137_n 0.00818434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_138_n 0.0121935f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_139_n 0.0282991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_130_n 0.00629939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_131_n 0.059011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A2_c_241_n 0.0268118f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_60 VPB N_A2_c_251_n 0.015356f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.16
cc_61 VPB N_A2_c_252_n 0.0152328f $X=-0.19 $Y=1.305 $X2=0.392 $Y2=1.53
cc_62 VPB N_A2_c_253_n 0.0189747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A2_c_246_n 0.00280652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A2_c_247_n 0.00198511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A2_c_256_n 0.013033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A2_c_248_n 0.0382325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A2_c_249_n 0.00733094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A1_c_372_n 0.0162831f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=0.995
cc_69 VPB N_A1_c_373_n 0.0158207f $X=-0.19 $Y=1.305 $X2=0.175 $Y2=1.445
cc_70 VPB N_A1_c_374_n 0.0161f $X=-0.19 $Y=1.305 $X2=0.392 $Y2=1.53
cc_71 VPB N_A1_c_375_n 0.015854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A1_c_370_n 0.00799673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A1_c_371_n 0.0253835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_440_n 0.00884045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_441_n 0.00547506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_442_n 0.060246f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_443_n 0.00538475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_444_n 0.01367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_445_n 0.0127542f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_446_n 0.0127781f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_447_n 0.0158513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_439_n 0.0523356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_449_n 0.0235893f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_450_n 0.00538475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_451_n 0.00547506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_227_297#_c_554_n 0.0107834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_227_297#_c_555_n 0.0135274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_Y_c_636_n 0.00274377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 B1_N N_A_27_47#_M1010_s 0.003021f $X=0.175 $Y=1.445 $X2=0 $Y2=0
cc_90 N_B1_N_c_92_n N_A_27_47#_c_123_n 0.0149279f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B1_N_c_91_n N_A_27_47#_c_127_n 0.00121693f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_92 B1_N N_A_27_47#_c_127_n 0.0202789f $X=0.175 $Y=1.445 $X2=0 $Y2=0
cc_93 N_B1_N_c_92_n N_A_27_47#_c_128_n 0.0106217f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B1_N_c_91_n N_A_27_47#_c_136_n 0.0171888f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_95 B1_N N_A_27_47#_c_136_n 0.0145323f $X=0.175 $Y=1.445 $X2=0 $Y2=0
cc_96 N_B1_N_c_91_n N_A_27_47#_c_149_n 0.00100586f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_97 N_B1_N_c_92_n N_A_27_47#_c_149_n 0.0169343f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_98 B1_N N_A_27_47#_c_149_n 0.0133962f $X=0.175 $Y=1.445 $X2=0 $Y2=0
cc_99 N_B1_N_c_92_n N_A_27_47#_c_129_n 0.0057172f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_100 B1_N N_A_27_47#_c_129_n 0.0030372f $X=0.175 $Y=1.445 $X2=0 $Y2=0
cc_101 N_B1_N_c_91_n N_A_27_47#_c_137_n 0.006996f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_102 B1_N N_A_27_47#_c_137_n 0.0219923f $X=0.175 $Y=1.445 $X2=0 $Y2=0
cc_103 N_B1_N_c_91_n N_A_27_47#_c_139_n 0.0117399f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_104 B1_N N_A_27_47#_c_139_n 0.0224148f $X=0.175 $Y=1.445 $X2=0 $Y2=0
cc_105 N_B1_N_c_91_n N_A_27_47#_c_130_n 0.00296664f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_106 B1_N N_A_27_47#_c_130_n 0.0271084f $X=0.175 $Y=1.445 $X2=0 $Y2=0
cc_107 N_B1_N_c_91_n N_A_27_47#_c_131_n 0.0149279f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_108 B1_N N_A_27_47#_c_131_n 2.47758e-19 $X=0.175 $Y=1.445 $X2=0 $Y2=0
cc_109 B1_N N_VPWR_M1010_d 0.00168767f $X=0.175 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_110 N_B1_N_c_91_n N_VPWR_c_440_n 0.00451579f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_111 N_B1_N_c_91_n N_VPWR_c_439_n 0.00898818f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B1_N_c_91_n N_VPWR_c_449_n 0.0051742f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B1_N_c_91_n N_A_227_297#_c_556_n 0.00439456f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B1_N_c_92_n N_VGND_c_727_n 0.00872204f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B1_N_c_92_n N_VGND_c_735_n 0.00705857f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_135_n N_A2_c_241_n 0.0303905f $X=2.99 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_117 N_A_27_47#_c_131_n N_A2_c_241_n 0.0242965f $X=2.645 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_118 N_A_27_47#_c_135_n N_A2_c_246_n 2.305e-19 $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_131_n N_A2_c_246_n 5.82523e-19 $X=2.645 $Y=1.202 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_135_n N_A2_c_263_n 8.31559e-19 $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_136_n N_VPWR_M1010_d 0.00834721f $X=0.84 $Y=1.895 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_27_47#_c_137_n N_VPWR_M1010_d 0.00358753f $X=0.925 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_123 N_A_27_47#_c_132_n N_VPWR_c_440_n 0.00208699f $X=1.55 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_136_n N_VPWR_c_440_n 0.0208991f $X=0.84 $Y=1.895 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_135_n N_VPWR_c_441_n 0.00101785f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_132_n N_VPWR_c_442_n 0.00429453f $X=1.55 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_133_n N_VPWR_c_442_n 0.00429362f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_134_n N_VPWR_c_442_n 0.00429201f $X=2.51 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_135_n N_VPWR_c_442_n 0.00429201f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_27_47#_c_136_n N_VPWR_c_442_n 0.0018132f $X=0.84 $Y=1.895 $X2=0 $Y2=0
cc_131 N_A_27_47#_M1010_s N_VPWR_c_439_n 0.00221616f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_132 N_A_27_47#_c_132_n N_VPWR_c_439_n 0.0073737f $X=1.55 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_133_n N_VPWR_c_439_n 0.00611667f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_27_47#_c_134_n N_VPWR_c_439_n 0.00611655f $X=2.51 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_135_n N_VPWR_c_439_n 0.00620861f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_136_n N_VPWR_c_439_n 0.00911427f $X=0.84 $Y=1.895 $X2=0
+ $Y2=0
cc_137 N_A_27_47#_c_139_n N_VPWR_c_439_n 0.0124954f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_136_n N_VPWR_c_449_n 0.00271905f $X=0.84 $Y=1.895 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_c_139_n N_VPWR_c_449_n 0.0210703f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_136_n N_A_227_297#_c_556_n 0.0178879f $X=0.84 $Y=1.895 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_c_138_n N_A_227_297#_c_556_n 0.00995594f $X=2.325 $Y=1.16
+ $X2=0 $Y2=0
cc_142 N_A_27_47#_c_131_n N_A_227_297#_c_556_n 0.00150138f $X=2.645 $Y=1.202
+ $X2=0 $Y2=0
cc_143 N_A_27_47#_c_132_n N_A_227_297#_c_560_n 0.0171395f $X=1.55 $Y=1.41 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_c_133_n N_A_227_297#_c_560_n 0.00841764f $X=2.03 $Y=1.41 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_c_133_n N_A_227_297#_c_562_n 0.00317151f $X=2.03 $Y=1.41 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_c_134_n N_A_227_297#_c_562_n 0.0116963f $X=2.51 $Y=1.41 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_c_135_n N_A_227_297#_c_562_n 0.0188757f $X=2.99 $Y=1.41 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_124_n N_Y_c_641_n 0.013028f $X=1.685 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_125_n N_Y_c_641_n 0.0115201f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_138_n N_Y_c_641_n 0.049103f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_131_n N_Y_c_641_n 0.00393251f $X=2.645 $Y=1.202 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_126_n N_Y_c_645_n 0.0148814f $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_138_n N_Y_c_645_n 0.00519128f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_131_n N_Y_c_645_n 0.00287285f $X=2.645 $Y=1.202 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_134_n N_Y_c_636_n 0.00386811f $X=2.51 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_126_n N_Y_c_636_n 0.00393201f $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_135_n N_Y_c_636_n 0.00491499f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_138_n N_Y_c_636_n 0.0216407f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_131_n N_Y_c_636_n 0.0270154f $X=2.645 $Y=1.202 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_123_n N_Y_c_653_n 0.00496059f $X=1.205 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_149_n N_Y_c_653_n 0.0116742f $X=0.84 $Y=0.705 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_129_n N_Y_c_653_n 0.00422784f $X=0.997 $Y=1.035 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_138_n N_Y_c_653_n 0.0145985f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_131_n N_Y_c_653_n 0.00374018f $X=2.645 $Y=1.202 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_138_n N_Y_c_658_n 0.0149565f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_131_n N_Y_c_658_n 0.00378594f $X=2.645 $Y=1.202 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_126_n N_Y_c_660_n 0.00133073f $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_133_n N_Y_c_661_n 0.0196012f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_134_n N_Y_c_661_n 0.0201998f $X=2.51 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_135_n N_Y_c_661_n 0.0142997f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_138_n N_Y_c_661_n 0.0516637f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_131_n N_Y_c_661_n 0.0103522f $X=2.645 $Y=1.202 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_149_n N_VGND_M1015_d 0.00422601f $X=0.84 $Y=0.705 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_27_47#_c_129_n N_VGND_M1015_d 0.00116387f $X=0.997 $Y=1.035 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A_27_47#_c_123_n N_VGND_c_727_n 0.00781765f $X=1.205 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_124_n N_VGND_c_727_n 8.10743e-19 $X=1.685 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_128_n N_VGND_c_727_n 0.0244675f $X=0.28 $Y=0.36 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_149_n N_VGND_c_727_n 0.0289997f $X=0.84 $Y=0.705 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_123_n N_VGND_c_730_n 0.00487821f $X=1.205 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_124_n N_VGND_c_730_n 0.00422112f $X=1.685 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_124_n N_VGND_c_732_n 0.00171872f $X=1.685 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_125_n N_VGND_c_732_n 0.00913379f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_126_n N_VGND_c_732_n 5.51597e-19 $X=2.645 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_125_n N_VGND_c_733_n 0.00211056f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_126_n N_VGND_c_733_n 0.00433717f $X=2.645 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_126_n N_VGND_c_734_n 0.00339683f $X=2.645 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_131_n N_VGND_c_734_n 0.00117746f $X=2.645 $Y=1.202 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_M1015_s N_VGND_c_735_n 0.00429487f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_123_n N_VGND_c_735_n 0.00843158f $X=1.205 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_124_n N_VGND_c_735_n 0.00590855f $X=1.685 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_125_n N_VGND_c_735_n 0.00284765f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_126_n N_VGND_c_735_n 0.00722501f $X=2.645 $Y=0.995 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_128_n N_VGND_c_735_n 0.0135138f $X=0.28 $Y=0.36 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_149_n N_VGND_c_735_n 0.0105612f $X=0.84 $Y=0.705 $X2=0 $Y2=0
cc_195 N_A2_c_242_n N_A1_c_366_n 0.0255706f $X=3.545 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_196 N_A2_c_241_n N_A1_c_372_n 0.0363522f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A2_c_246_n N_A1_c_372_n 0.00164446f $X=3.465 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A2_c_256_n N_A1_c_372_n 0.0143516f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_199 N_A2_c_256_n N_A1_c_373_n 0.0143377f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_200 N_A2_c_256_n N_A1_c_374_n 0.0143377f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_201 N_A2_c_251_n N_A1_c_375_n 0.0391028f $X=5.9 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A2_c_247_n N_A1_c_375_n 0.0018629f $X=6.04 $Y=1.39 $X2=0 $Y2=0
cc_203 N_A2_c_256_n N_A1_c_375_n 0.0167504f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_204 N_A2_c_243_n N_A1_c_369_n 0.0235788f $X=5.875 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A2_c_241_n N_A1_c_370_n 8.87839e-19 $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A2_c_246_n N_A1_c_370_n 0.021768f $X=3.465 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A2_c_247_n N_A1_c_370_n 0.0140887f $X=6.04 $Y=1.39 $X2=0 $Y2=0
cc_208 N_A2_c_256_n N_A1_c_370_n 0.119243f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_209 N_A2_c_248_n N_A1_c_370_n 2.90736e-19 $X=6.875 $Y=1.202 $X2=0 $Y2=0
cc_210 N_A2_c_241_n N_A1_c_371_n 0.0258418f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A2_c_246_n N_A1_c_371_n 0.00318127f $X=3.465 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A2_c_247_n N_A1_c_371_n 0.00480287f $X=6.04 $Y=1.39 $X2=0 $Y2=0
cc_213 N_A2_c_256_n N_A1_c_371_n 0.00833524f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_214 N_A2_c_248_n N_A1_c_371_n 0.0235788f $X=6.875 $Y=1.202 $X2=0 $Y2=0
cc_215 N_A2_c_263_n N_VPWR_M1003_d 5.2043e-19 $X=3.695 $Y=1.592 $X2=0 $Y2=0
cc_216 N_A2_c_256_n N_VPWR_M1003_d 0.00158005f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_217 N_A2_c_256_n N_VPWR_M1017_d 0.00199924f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_218 N_A2_c_247_n N_VPWR_M1024_d 3.10624e-19 $X=6.04 $Y=1.39 $X2=0 $Y2=0
cc_219 N_A2_c_256_n N_VPWR_M1024_d 0.00158005f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_220 N_A2_c_249_n N_VPWR_M1011_d 0.00195249f $X=6.905 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A2_c_241_n N_VPWR_c_441_n 0.00947287f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A2_c_241_n N_VPWR_c_442_n 0.0035176f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A2_c_251_n N_VPWR_c_446_n 0.00436183f $X=5.9 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A2_c_252_n N_VPWR_c_446_n 0.00379901f $X=6.37 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A2_c_253_n N_VPWR_c_447_n 0.00379901f $X=6.84 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A2_c_241_n N_VPWR_c_439_n 0.00421648f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A2_c_251_n N_VPWR_c_439_n 0.00494532f $X=5.9 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A2_c_252_n N_VPWR_c_439_n 0.00438112f $X=6.37 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A2_c_253_n N_VPWR_c_439_n 0.00531504f $X=6.84 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A2_c_251_n N_VPWR_c_450_n 0.00682926f $X=5.9 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A2_c_252_n N_VPWR_c_450_n 4.93764e-19 $X=6.37 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A2_c_251_n N_VPWR_c_451_n 5.09137e-19 $X=5.9 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A2_c_252_n N_VPWR_c_451_n 0.00783739f $X=6.37 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A2_c_253_n N_VPWR_c_451_n 0.00943405f $X=6.84 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A2_c_263_n N_A_227_297#_M1022_d 0.00251451f $X=3.695 $Y=1.592 $X2=0
+ $Y2=0
cc_236 N_A2_c_256_n N_A_227_297#_M1014_s 0.00199924f $X=5.725 $Y=1.39 $X2=0
+ $Y2=0
cc_237 N_A2_c_256_n N_A_227_297#_M1021_s 0.00199437f $X=5.725 $Y=1.39 $X2=0
+ $Y2=0
cc_238 N_A2_c_249_n N_A_227_297#_M1006_s 0.00191452f $X=6.905 $Y=1.16 $X2=0
+ $Y2=0
cc_239 N_A2_c_249_n N_A_227_297#_M1023_s 0.011381f $X=6.905 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A2_c_241_n N_A_227_297#_c_570_n 0.0153931f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A2_c_263_n N_A_227_297#_c_570_n 0.0179009f $X=3.695 $Y=1.592 $X2=0
+ $Y2=0
cc_242 N_A2_c_256_n N_A_227_297#_c_570_n 0.0775879f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_243 N_A2_c_241_n N_A_227_297#_c_562_n 2.09297e-19 $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A2_c_263_n N_A_227_297#_c_562_n 0.00470781f $X=3.695 $Y=1.592 $X2=0
+ $Y2=0
cc_245 N_A2_c_251_n N_A_227_297#_c_575_n 0.0156963f $X=5.9 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A2_c_256_n N_A_227_297#_c_575_n 0.0401943f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_247 N_A2_c_252_n N_A_227_297#_c_577_n 0.015582f $X=6.37 $Y=1.41 $X2=0 $Y2=0
cc_248 N_A2_c_253_n N_A_227_297#_c_577_n 0.0127186f $X=6.84 $Y=1.41 $X2=0 $Y2=0
cc_249 N_A2_c_248_n N_A_227_297#_c_577_n 7.66811e-19 $X=6.875 $Y=1.202 $X2=0
+ $Y2=0
cc_250 N_A2_c_249_n N_A_227_297#_c_577_n 0.0422494f $X=6.905 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A2_c_248_n N_A_227_297#_c_554_n 3.55007e-19 $X=6.875 $Y=1.202 $X2=0
+ $Y2=0
cc_252 N_A2_c_249_n N_A_227_297#_c_554_n 0.0114802f $X=6.905 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A2_c_256_n N_A_227_297#_c_583_n 0.0152498f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_254 N_A2_c_248_n N_A_227_297#_c_584_n 6.3906e-19 $X=6.875 $Y=1.202 $X2=0
+ $Y2=0
cc_255 N_A2_c_249_n N_A_227_297#_c_584_n 0.0152772f $X=6.905 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A2_c_241_n N_Y_c_636_n 0.00362136f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A2_c_242_n N_Y_c_636_n 0.00304074f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A2_c_246_n N_Y_c_636_n 0.0337243f $X=3.465 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A2_c_263_n N_Y_c_636_n 0.0048869f $X=3.695 $Y=1.592 $X2=0 $Y2=0
cc_260 N_A2_c_241_n N_Y_c_637_n 0.001467f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A2_c_242_n N_Y_c_637_n 0.00653244f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A2_c_256_n N_Y_c_638_n 0.00563538f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_263 N_A2_c_241_n N_Y_c_661_n 9.28308e-19 $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A2_c_241_n N_Y_c_639_n 0.00443783f $X=3.5 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A2_c_242_n N_Y_c_639_n 0.00953835f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A2_c_246_n N_Y_c_639_n 0.0311154f $X=3.465 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A2_c_243_n N_VGND_c_724_n 0.00519429f $X=5.875 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A2_c_244_n N_VGND_c_724_n 0.00289125f $X=6.395 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A2_c_245_n N_VGND_c_726_n 0.00448362f $X=6.875 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A2_c_248_n N_VGND_c_726_n 0.00223987f $X=6.875 $Y=1.202 $X2=0 $Y2=0
cc_271 N_A2_c_249_n N_VGND_c_726_n 0.0093319f $X=6.905 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A2_c_242_n N_VGND_c_728_n 0.00405721f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A2_c_243_n N_VGND_c_728_n 0.00403873f $X=5.875 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A2_c_244_n N_VGND_c_731_n 0.00427134f $X=6.395 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A2_c_245_n N_VGND_c_731_n 0.0054895f $X=6.875 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A2_c_242_n N_VGND_c_734_n 0.00640935f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A2_c_242_n N_VGND_c_735_n 0.006975f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A2_c_243_n N_VGND_c_735_n 0.00599083f $X=5.875 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A2_c_244_n N_VGND_c_735_n 0.00614542f $X=6.395 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A2_c_245_n N_VGND_c_735_n 0.0108057f $X=6.875 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A2_c_242_n N_A_724_47#_c_829_n 0.00442984f $X=3.545 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A2_c_243_n N_A_724_47#_c_830_n 0.0040881f $X=5.875 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A2_c_243_n N_A_724_47#_c_831_n 0.00593154f $X=5.875 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A2_c_244_n N_A_724_47#_c_831_n 5.01809e-19 $X=6.395 $Y=0.995 $X2=0
+ $Y2=0
cc_285 N_A2_c_243_n N_A_724_47#_c_827_n 0.00712827f $X=5.875 $Y=0.995 $X2=0
+ $Y2=0
cc_286 N_A2_c_244_n N_A_724_47#_c_827_n 0.0102615f $X=6.395 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A2_c_245_n N_A_724_47#_c_827_n 0.00317383f $X=6.875 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_A2_c_247_n N_A_724_47#_c_827_n 0.0449578f $X=6.04 $Y=1.39 $X2=0 $Y2=0
cc_289 N_A2_c_248_n N_A_724_47#_c_827_n 0.00852195f $X=6.875 $Y=1.202 $X2=0
+ $Y2=0
cc_290 N_A2_c_249_n N_A_724_47#_c_827_n 0.0331939f $X=6.905 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A2_c_243_n N_A_724_47#_c_828_n 0.00337814f $X=5.875 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_A2_c_247_n N_A_724_47#_c_828_n 0.0123571f $X=6.04 $Y=1.39 $X2=0 $Y2=0
cc_293 N_A2_c_256_n N_A_724_47#_c_828_n 0.00438828f $X=5.725 $Y=1.39 $X2=0 $Y2=0
cc_294 N_A2_c_243_n N_A_724_47#_c_842_n 5.87718e-19 $X=5.875 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_A2_c_244_n N_A_724_47#_c_842_n 0.00653659f $X=6.395 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A2_c_245_n N_A_724_47#_c_842_n 0.00536147f $X=6.875 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A1_c_372_n N_VPWR_c_441_n 0.00772308f $X=3.99 $Y=1.41 $X2=0 $Y2=0
cc_298 N_A1_c_373_n N_VPWR_c_441_n 0.00100586f $X=4.47 $Y=1.41 $X2=0 $Y2=0
cc_299 N_A1_c_372_n N_VPWR_c_443_n 0.00111962f $X=3.99 $Y=1.41 $X2=0 $Y2=0
cc_300 N_A1_c_373_n N_VPWR_c_443_n 0.0105269f $X=4.47 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A1_c_374_n N_VPWR_c_443_n 0.00636819f $X=4.95 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A1_c_375_n N_VPWR_c_443_n 4.76818e-19 $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A1_c_372_n N_VPWR_c_444_n 0.00464324f $X=3.99 $Y=1.41 $X2=0 $Y2=0
cc_304 N_A1_c_373_n N_VPWR_c_444_n 0.0032362f $X=4.47 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A1_c_374_n N_VPWR_c_445_n 0.00464324f $X=4.95 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A1_c_375_n N_VPWR_c_445_n 0.0032362f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A1_c_372_n N_VPWR_c_439_n 0.00529844f $X=3.99 $Y=1.41 $X2=0 $Y2=0
cc_308 N_A1_c_373_n N_VPWR_c_439_n 0.00388795f $X=4.47 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A1_c_374_n N_VPWR_c_439_n 0.00525281f $X=4.95 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A1_c_375_n N_VPWR_c_439_n 0.00384231f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A1_c_374_n N_VPWR_c_450_n 5.25185e-19 $X=4.95 $Y=1.41 $X2=0 $Y2=0
cc_312 N_A1_c_375_n N_VPWR_c_450_n 0.00888881f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_313 N_A1_c_372_n N_A_227_297#_c_570_n 0.0130725f $X=3.99 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A1_c_373_n N_A_227_297#_c_570_n 0.0126261f $X=4.47 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A1_c_374_n N_A_227_297#_c_570_n 0.0130581f $X=4.95 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A1_c_375_n N_A_227_297#_c_575_n 0.0124874f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A1_c_366_n N_Y_c_638_n 0.0128587f $X=3.965 $Y=0.99 $X2=0 $Y2=0
cc_318 N_A1_c_367_n N_Y_c_638_n 0.010275f $X=4.475 $Y=0.99 $X2=0 $Y2=0
cc_319 N_A1_c_368_n N_Y_c_638_n 0.0102726f $X=4.955 $Y=0.99 $X2=0 $Y2=0
cc_320 N_A1_c_369_n N_Y_c_638_n 0.00233957f $X=5.455 $Y=0.99 $X2=0 $Y2=0
cc_321 N_A1_c_370_n N_Y_c_638_n 0.112319f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A1_c_371_n N_Y_c_638_n 0.0121329f $X=5.43 $Y=1.2 $X2=0 $Y2=0
cc_323 N_A1_c_366_n N_VGND_c_728_n 0.00357877f $X=3.965 $Y=0.99 $X2=0 $Y2=0
cc_324 N_A1_c_367_n N_VGND_c_728_n 0.00357877f $X=4.475 $Y=0.99 $X2=0 $Y2=0
cc_325 N_A1_c_368_n N_VGND_c_728_n 0.00357877f $X=4.955 $Y=0.99 $X2=0 $Y2=0
cc_326 N_A1_c_369_n N_VGND_c_728_n 0.00357877f $X=5.455 $Y=0.99 $X2=0 $Y2=0
cc_327 N_A1_c_366_n N_VGND_c_735_n 0.00548096f $X=3.965 $Y=0.99 $X2=0 $Y2=0
cc_328 N_A1_c_367_n N_VGND_c_735_n 0.00560469f $X=4.475 $Y=0.99 $X2=0 $Y2=0
cc_329 N_A1_c_368_n N_VGND_c_735_n 0.00558119f $X=4.955 $Y=0.99 $X2=0 $Y2=0
cc_330 N_A1_c_369_n N_VGND_c_735_n 0.00545746f $X=5.455 $Y=0.99 $X2=0 $Y2=0
cc_331 N_A1_c_366_n N_A_724_47#_c_829_n 0.0104539f $X=3.965 $Y=0.99 $X2=0 $Y2=0
cc_332 N_A1_c_367_n N_A_724_47#_c_829_n 0.0104539f $X=4.475 $Y=0.99 $X2=0 $Y2=0
cc_333 N_A1_c_368_n N_A_724_47#_c_829_n 0.0103796f $X=4.955 $Y=0.99 $X2=0 $Y2=0
cc_334 N_A1_c_369_n N_A_724_47#_c_829_n 0.0139648f $X=5.455 $Y=0.99 $X2=0 $Y2=0
cc_335 N_A1_c_370_n N_A_724_47#_c_829_n 0.00148199f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A1_c_369_n N_A_724_47#_c_831_n 0.00452349f $X=5.455 $Y=0.99 $X2=0 $Y2=0
cc_337 N_A1_c_369_n N_A_724_47#_c_828_n 0.00170282f $X=5.455 $Y=0.99 $X2=0 $Y2=0
cc_338 N_VPWR_c_439_n N_A_227_297#_M1005_d 0.0041883f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_339 N_VPWR_c_439_n N_A_227_297#_M1008_d 0.00239291f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_439_n N_A_227_297#_M1022_d 0.00278173f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_439_n N_A_227_297#_M1014_s 0.00341753f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_439_n N_A_227_297#_M1021_s 0.00273993f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_439_n N_A_227_297#_M1006_s 0.00264282f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_439_n N_A_227_297#_M1023_s 0.00244747f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_440_n N_A_227_297#_c_597_n 0.0150677f $X=0.74 $Y=2.34 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_442_n N_A_227_297#_c_597_n 0.0164451f $X=3.535 $Y=2.72 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_439_n N_A_227_297#_c_597_n 0.00943173f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_440_n N_A_227_297#_c_556_n 0.00220009f $X=0.74 $Y=2.34 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_442_n N_A_227_297#_c_560_n 0.0359212f $X=3.535 $Y=2.72 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_439_n N_A_227_297#_c_560_n 0.0222394f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_351 N_VPWR_M1003_d N_A_227_297#_c_570_n 0.00408766f $X=3.59 $Y=1.485 $X2=0
+ $Y2=0
cc_352 N_VPWR_M1017_d N_A_227_297#_c_570_n 0.00373237f $X=4.56 $Y=1.485 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_441_n N_A_227_297#_c_570_n 0.0199956f $X=3.75 $Y=2.36 $X2=0
+ $Y2=0
cc_354 N_VPWR_c_442_n N_A_227_297#_c_570_n 0.00264869f $X=3.535 $Y=2.72 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_443_n N_A_227_297#_c_570_n 0.0199464f $X=4.71 $Y=2.36 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_444_n N_A_227_297#_c_570_n 0.00952824f $X=4.495 $Y=2.72 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_445_n N_A_227_297#_c_570_n 0.00344373f $X=5.455 $Y=2.72 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_439_n N_A_227_297#_c_570_n 0.0289096f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_442_n N_A_227_297#_c_562_n 0.0768983f $X=3.535 $Y=2.72 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_439_n N_A_227_297#_c_562_n 0.0472839f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_361 N_VPWR_c_445_n N_A_227_297#_c_613_n 0.0130156f $X=5.455 $Y=2.72 $X2=0
+ $Y2=0
cc_362 N_VPWR_c_439_n N_A_227_297#_c_613_n 0.00720328f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_363 N_VPWR_M1024_d N_A_227_297#_c_575_n 0.00370274f $X=5.52 $Y=1.485 $X2=0
+ $Y2=0
cc_364 N_VPWR_c_445_n N_A_227_297#_c_575_n 0.00256992f $X=5.455 $Y=2.72 $X2=0
+ $Y2=0
cc_365 N_VPWR_c_446_n N_A_227_297#_c_575_n 0.0033277f $X=6.415 $Y=2.72 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_439_n N_A_227_297#_c_575_n 0.0115583f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_450_n N_A_227_297#_c_575_n 0.0198971f $X=5.665 $Y=2.36 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_446_n N_A_227_297#_c_620_n 0.0123606f $X=6.415 $Y=2.72 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_439_n N_A_227_297#_c_620_n 0.0070216f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_450_n N_A_227_297#_c_620_n 0.0119105f $X=5.665 $Y=2.36 $X2=0
+ $Y2=0
cc_371 N_VPWR_M1011_d N_A_227_297#_c_577_n 0.00351756f $X=6.46 $Y=1.485 $X2=0
+ $Y2=0
cc_372 N_VPWR_c_446_n N_A_227_297#_c_577_n 0.00282346f $X=6.415 $Y=2.72 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_447_n N_A_227_297#_c_577_n 0.00297102f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_439_n N_A_227_297#_c_577_n 0.0112672f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_451_n N_A_227_297#_c_577_n 0.0198971f $X=6.605 $Y=2.36 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_447_n N_A_227_297#_c_555_n 0.0172982f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_439_n N_A_227_297#_c_555_n 0.00951562f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_451_n N_A_227_297#_c_555_n 0.0131293f $X=6.605 $Y=2.36 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_439_n N_Y_M1005_s 0.00240926f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_380 N_VPWR_c_439_n N_Y_M1016_s 0.00240897f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_381 N_A_227_297#_c_560_n N_Y_M1005_s 0.00382218f $X=2.055 $Y=2.34 $X2=0 $Y2=0
cc_382 N_A_227_297#_c_562_n N_Y_M1016_s 0.00375879f $X=3.365 $Y=1.99 $X2=0 $Y2=0
cc_383 N_A_227_297#_M1008_d N_Y_c_661_n 0.0038817f $X=2.12 $Y=1.485 $X2=0 $Y2=0
cc_384 N_A_227_297#_c_560_n N_Y_c_661_n 0.0213875f $X=2.055 $Y=2.34 $X2=0 $Y2=0
cc_385 N_A_227_297#_c_562_n N_Y_c_661_n 0.065672f $X=3.365 $Y=1.99 $X2=0 $Y2=0
cc_386 N_Y_c_641_n N_VGND_M1018_d 0.00419317f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_387 N_Y_c_645_n N_VGND_M1025_d 9.1036e-19 $X=2.82 $Y=0.78 $X2=0 $Y2=0
cc_388 N_Y_c_660_n N_VGND_M1025_d 0.00513258f $X=2.975 $Y=0.795 $X2=0 $Y2=0
cc_389 N_Y_c_639_n N_VGND_M1025_d 0.00429242f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_390 N_Y_c_653_n N_VGND_c_727_n 0.00463323f $X=1.47 $Y=0.535 $X2=0 $Y2=0
cc_391 N_Y_c_639_n N_VGND_c_728_n 0.00212611f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_392 N_Y_c_641_n N_VGND_c_730_n 0.00335005f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_393 N_Y_c_653_n N_VGND_c_730_n 0.0071941f $X=1.47 $Y=0.535 $X2=0 $Y2=0
cc_394 N_Y_c_641_n N_VGND_c_732_n 0.0221395f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_395 N_Y_c_699_p N_VGND_c_732_n 0.0143006f $X=2.43 $Y=0.42 $X2=0 $Y2=0
cc_396 N_Y_c_641_n N_VGND_c_733_n 0.00260346f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_397 N_Y_c_699_p N_VGND_c_733_n 0.0127385f $X=2.43 $Y=0.42 $X2=0 $Y2=0
cc_398 N_Y_c_645_n N_VGND_c_733_n 0.00271527f $X=2.82 $Y=0.78 $X2=0 $Y2=0
cc_399 N_Y_c_645_n N_VGND_c_734_n 0.00328838f $X=2.82 $Y=0.78 $X2=0 $Y2=0
cc_400 N_Y_c_660_n N_VGND_c_734_n 0.0264543f $X=2.975 $Y=0.795 $X2=0 $Y2=0
cc_401 N_Y_c_639_n N_VGND_c_734_n 0.0198737f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_402 N_Y_M1002_s N_VGND_c_735_n 0.00621961f $X=1.28 $Y=0.235 $X2=0 $Y2=0
cc_403 N_Y_M1019_s N_VGND_c_735_n 0.00315407f $X=2.24 $Y=0.235 $X2=0 $Y2=0
cc_404 N_Y_M1007_d N_VGND_c_735_n 0.00289111f $X=4.04 $Y=0.235 $X2=0 $Y2=0
cc_405 N_Y_M1013_d N_VGND_c_735_n 0.0028108f $X=5.03 $Y=0.235 $X2=0 $Y2=0
cc_406 N_Y_c_641_n N_VGND_c_735_n 0.0119527f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_407 N_Y_c_699_p N_VGND_c_735_n 0.00721967f $X=2.43 $Y=0.42 $X2=0 $Y2=0
cc_408 N_Y_c_645_n N_VGND_c_735_n 0.00538517f $X=2.82 $Y=0.78 $X2=0 $Y2=0
cc_409 N_Y_c_637_n N_VGND_c_735_n 0.00351546f $X=3.665 $Y=0.785 $X2=0 $Y2=0
cc_410 N_Y_c_653_n N_VGND_c_735_n 0.00672198f $X=1.47 $Y=0.535 $X2=0 $Y2=0
cc_411 N_Y_c_660_n N_VGND_c_735_n 0.00141155f $X=2.975 $Y=0.795 $X2=0 $Y2=0
cc_412 N_Y_c_639_n N_VGND_c_735_n 0.00519342f $X=3.555 $Y=0.785 $X2=0 $Y2=0
cc_413 N_Y_c_638_n N_A_724_47#_M1000_d 0.00162311f $X=5.22 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_414 N_Y_c_638_n N_A_724_47#_M1009_s 0.00224739f $X=5.22 $Y=0.76 $X2=0 $Y2=0
cc_415 N_Y_M1007_d N_A_724_47#_c_829_n 0.00476658f $X=4.04 $Y=0.235 $X2=0 $Y2=0
cc_416 N_Y_M1013_d N_A_724_47#_c_829_n 0.00457616f $X=5.03 $Y=0.235 $X2=0 $Y2=0
cc_417 N_Y_c_637_n N_A_724_47#_c_829_n 0.0967035f $X=3.665 $Y=0.785 $X2=0 $Y2=0
cc_418 N_Y_c_638_n N_A_724_47#_c_831_n 0.00388125f $X=5.22 $Y=0.76 $X2=0 $Y2=0
cc_419 N_Y_c_638_n N_A_724_47#_c_828_n 0.0113909f $X=5.22 $Y=0.76 $X2=0 $Y2=0
cc_420 N_VGND_c_735_n N_A_724_47#_M1000_d 0.00215227f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_421 N_VGND_c_735_n N_A_724_47#_M1009_s 0.00263412f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_735_n N_A_724_47#_M1020_s 0.00215208f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_735_n N_A_724_47#_M1004_d 0.0026338f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_728_n N_A_724_47#_c_829_n 0.116003f $X=6.085 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_734_n N_A_724_47#_c_829_n 0.0206335f $X=3.385 $Y=0.22 $X2=0
+ $Y2=0
cc_426 N_VGND_c_735_n N_A_724_47#_c_829_n 0.0732792f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_724_n N_A_724_47#_c_830_n 0.0162144f $X=6.18 $Y=0.4 $X2=0 $Y2=0
cc_428 N_VGND_c_728_n N_A_724_47#_c_830_n 0.0160793f $X=6.085 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_735_n N_A_724_47#_c_830_n 0.0096316f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_724_n N_A_724_47#_c_831_n 0.00356776f $X=6.18 $Y=0.4 $X2=0 $Y2=0
cc_431 N_VGND_M1001_s N_A_724_47#_c_827_n 0.00343275f $X=5.95 $Y=0.235 $X2=0
+ $Y2=0
cc_432 N_VGND_c_724_n N_A_724_47#_c_827_n 0.0138893f $X=6.18 $Y=0.4 $X2=0 $Y2=0
cc_433 N_VGND_c_728_n N_A_724_47#_c_827_n 0.00263884f $X=6.085 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_731_n N_A_724_47#_c_827_n 0.00196536f $X=7 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_735_n N_A_724_47#_c_827_n 0.00987199f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_731_n N_A_724_47#_c_842_n 0.0223809f $X=7 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_735_n N_A_724_47#_c_842_n 0.014176f $X=7.13 $Y=0 $X2=0 $Y2=0
