* File: sky130_fd_sc_hdll__or3_2.pxi.spice
* Created: Wed Sep  2 08:48:35 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR3_2%C N_C_c_62_n N_C_M1001_g N_C_M1008_g C N_C_c_61_n
+ PM_SKY130_FD_SC_HDLL__OR3_2%C
x_PM_SKY130_FD_SC_HDLL__OR3_2%B N_B_c_84_n N_B_c_87_n N_B_c_88_n N_B_M1009_g
+ N_B_M1004_g N_B_c_85_n N_B_c_86_n B B B B B PM_SKY130_FD_SC_HDLL__OR3_2%B
x_PM_SKY130_FD_SC_HDLL__OR3_2%A N_A_c_128_n N_A_M1006_g N_A_M1002_g A A A
+ N_A_c_130_n A N_A_c_131_n PM_SKY130_FD_SC_HDLL__OR3_2%A
x_PM_SKY130_FD_SC_HDLL__OR3_2%A_30_53# N_A_30_53#_M1008_s N_A_30_53#_M1004_d
+ N_A_30_53#_M1001_s N_A_30_53#_c_179_n N_A_30_53#_M1000_g N_A_30_53#_c_189_n
+ N_A_30_53#_M1003_g N_A_30_53#_c_190_n N_A_30_53#_M1005_g N_A_30_53#_c_180_n
+ N_A_30_53#_M1007_g N_A_30_53#_c_181_n N_A_30_53#_c_191_n N_A_30_53#_c_182_n
+ N_A_30_53#_c_183_n N_A_30_53#_c_192_n N_A_30_53#_c_193_n N_A_30_53#_c_279_p
+ N_A_30_53#_c_184_n N_A_30_53#_c_212_n N_A_30_53#_c_185_n N_A_30_53#_c_194_n
+ N_A_30_53#_c_186_n N_A_30_53#_c_195_n N_A_30_53#_c_187_n N_A_30_53#_c_188_n
+ PM_SKY130_FD_SC_HDLL__OR3_2%A_30_53#
x_PM_SKY130_FD_SC_HDLL__OR3_2%VPWR N_VPWR_M1006_d N_VPWR_M1005_d N_VPWR_c_296_n
+ N_VPWR_c_297_n N_VPWR_c_298_n VPWR N_VPWR_c_299_n N_VPWR_c_300_n
+ N_VPWR_c_301_n N_VPWR_c_295_n PM_SKY130_FD_SC_HDLL__OR3_2%VPWR
x_PM_SKY130_FD_SC_HDLL__OR3_2%X N_X_M1000_s N_X_M1003_s N_X_c_328_n N_X_c_331_n
+ N_X_c_326_n X PM_SKY130_FD_SC_HDLL__OR3_2%X
x_PM_SKY130_FD_SC_HDLL__OR3_2%VGND N_VGND_M1008_d N_VGND_M1002_d N_VGND_M1007_d
+ N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n VGND N_VGND_c_358_n
+ N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n
+ PM_SKY130_FD_SC_HDLL__OR3_2%VGND
cc_1 VNB N_C_M1008_g 0.0347457f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.475
cc_2 VNB C 0.0147109f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_C_c_61_n 0.0375861f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.202
cc_4 VNB N_B_c_84_n 0.0186323f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.695
cc_5 VNB N_B_c_85_n 0.0147582f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.202
cc_6 VNB N_B_c_86_n 0.0136004f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_7 VNB N_A_c_128_n 0.026579f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.41
cc_8 VNB N_A_M1002_g 0.0296069f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.475
cc_9 VNB N_A_c_130_n 0.00216296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_c_131_n 0.00196889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_30_53#_c_179_n 0.0184705f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.202
cc_12 VNB N_A_30_53#_c_180_n 0.0216421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_30_53#_c_181_n 0.0135183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_30_53#_c_182_n 0.00324292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_30_53#_c_183_n 0.00940378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_30_53#_c_184_n 0.00135955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_30_53#_c_185_n 0.00183221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_30_53#_c_186_n 0.00149272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_30_53#_c_187_n 0.00311809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_30_53#_c_188_n 0.0503474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_295_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_326_n 8.88908e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_355_n 0.00289919f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_24 VNB N_VGND_c_356_n 0.0111284f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.202
cc_25 VNB N_VGND_c_357_n 0.0369869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_358_n 0.0152668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_359_n 0.0199552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_360_n 0.00602632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_361_n 0.0137871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_362_n 0.0111386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_363_n 0.187351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_C_c_62_n 0.019972f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_33 VPB C 0.00405604f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_34 VPB N_C_c_61_n 0.0174587f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.202
cc_35 VPB N_B_c_87_n 0.00562437f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.695
cc_36 VPB N_B_c_88_n 0.0498999f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=0.995
cc_37 VPB N_B_M1009_g 0.0107136f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=0.475
cc_38 VPB B 0.0381946f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.202
cc_39 VPB N_A_c_128_n 0.0303869f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_40 VPB N_A_c_130_n 0.00322575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_30_53#_c_189_n 0.0190729f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.202
cc_42 VPB N_A_30_53#_c_190_n 0.0193182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_30_53#_c_191_n 0.011323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_30_53#_c_192_n 0.00349637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_30_53#_c_193_n 0.00979957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_30_53#_c_194_n 0.00242774f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_30_53#_c_195_n 0.00148365f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_30_53#_c_187_n 6.91143e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_30_53#_c_188_n 0.0249876f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_296_n 0.014331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_297_n 0.0110992f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_52 VPB N_VPWR_c_298_n 0.0510195f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.202
cc_53 VPB N_VPWR_c_299_n 0.0420274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_300_n 0.0207755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_301_n 0.00901444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_295_n 0.0595004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_X_c_326_n 0.00126197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 N_C_c_61_n N_B_c_84_n 0.0212841f $X=0.51 $Y=1.202 $X2=0 $Y2=0
cc_59 N_C_c_62_n N_B_M1009_g 0.035952f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_60 N_C_M1008_g N_B_c_85_n 0.0112369f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_61 N_C_M1008_g N_B_c_86_n 0.0212841f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_62 N_C_c_62_n B 0.00527095f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_63 N_C_c_62_n N_A_c_131_n 0.00799389f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_64 C N_A_c_131_n 0.0245564f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_65 N_C_c_61_n N_A_c_131_n 0.0149939f $X=0.51 $Y=1.202 $X2=0 $Y2=0
cc_66 C N_A_30_53#_c_191_n 0.0216023f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_67 N_C_c_61_n N_A_30_53#_c_191_n 0.00195431f $X=0.51 $Y=1.202 $X2=0 $Y2=0
cc_68 N_C_M1008_g N_A_30_53#_c_182_n 0.0152773f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_69 C N_A_30_53#_c_182_n 0.00177486f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_70 N_C_c_61_n N_A_30_53#_c_182_n 0.0031905f $X=0.51 $Y=1.202 $X2=0 $Y2=0
cc_71 C N_A_30_53#_c_183_n 0.0212035f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_72 N_C_c_61_n N_A_30_53#_c_183_n 0.00184772f $X=0.51 $Y=1.202 $X2=0 $Y2=0
cc_73 N_C_c_62_n N_A_30_53#_c_192_n 0.0138675f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_74 N_C_M1008_g N_VGND_c_355_n 0.0124881f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_75 N_C_M1008_g N_VGND_c_358_n 0.00187556f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_76 N_C_M1008_g N_VGND_c_363_n 0.00331269f $X=0.535 $Y=0.475 $X2=0 $Y2=0
cc_77 N_B_c_84_n N_A_c_128_n 0.0167852f $X=0.92 $Y=1.31 $X2=-0.19 $Y2=-0.24
cc_78 N_B_c_87_n N_A_c_128_n 0.00343361f $X=0.92 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_79 N_B_M1009_g N_A_c_128_n 0.0206987f $X=0.92 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_80 B N_A_c_128_n 6.44478e-19 $X=1.085 $Y=2.15 $X2=-0.19 $Y2=-0.24
cc_81 N_B_c_84_n N_A_M1002_g 0.00330916f $X=0.92 $Y=1.31 $X2=0 $Y2=0
cc_82 N_B_c_85_n N_A_M1002_g 0.015811f $X=0.95 $Y=0.76 $X2=0 $Y2=0
cc_83 N_B_c_84_n N_A_c_130_n 0.0103585f $X=0.92 $Y=1.31 $X2=0 $Y2=0
cc_84 N_B_c_87_n N_A_c_130_n 0.00369388f $X=0.92 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B_c_86_n N_A_c_130_n 0.00177283f $X=0.95 $Y=0.91 $X2=0 $Y2=0
cc_86 N_B_c_84_n N_A_c_131_n 0.00632891f $X=0.92 $Y=1.31 $X2=0 $Y2=0
cc_87 N_B_c_87_n N_A_c_131_n 0.00309614f $X=0.92 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B_M1009_g N_A_c_131_n 0.00648038f $X=0.92 $Y=1.695 $X2=0 $Y2=0
cc_89 N_B_c_85_n N_A_30_53#_c_182_n 0.00747646f $X=0.95 $Y=0.76 $X2=0 $Y2=0
cc_90 N_B_c_86_n N_A_30_53#_c_182_n 0.00793181f $X=0.95 $Y=0.91 $X2=0 $Y2=0
cc_91 N_B_c_88_n N_A_30_53#_c_192_n 0.00124804f $X=0.92 $Y=2.035 $X2=0 $Y2=0
cc_92 N_B_M1009_g N_A_30_53#_c_192_n 0.0123508f $X=0.92 $Y=1.695 $X2=0 $Y2=0
cc_93 B N_A_30_53#_c_192_n 0.059861f $X=1.085 $Y=2.15 $X2=0 $Y2=0
cc_94 B N_A_30_53#_c_193_n 0.0230159f $X=1.085 $Y=2.15 $X2=0 $Y2=0
cc_95 B N_A_30_53#_c_212_n 3.54753e-19 $X=1.085 $Y=2.15 $X2=0 $Y2=0
cc_96 N_B_M1009_g N_A_30_53#_c_195_n 0.00472277f $X=0.92 $Y=1.695 $X2=0 $Y2=0
cc_97 B N_A_30_53#_c_195_n 0.0137701f $X=1.085 $Y=2.15 $X2=0 $Y2=0
cc_98 N_B_c_88_n N_VPWR_c_296_n 0.00371783f $X=0.92 $Y=2.035 $X2=0 $Y2=0
cc_99 B N_VPWR_c_296_n 0.0218015f $X=1.085 $Y=2.15 $X2=0 $Y2=0
cc_100 N_B_c_88_n N_VPWR_c_299_n 0.00793506f $X=0.92 $Y=2.035 $X2=0 $Y2=0
cc_101 B N_VPWR_c_299_n 0.0649251f $X=1.085 $Y=2.15 $X2=0 $Y2=0
cc_102 N_B_c_88_n N_VPWR_c_295_n 0.0113914f $X=0.92 $Y=2.035 $X2=0 $Y2=0
cc_103 B N_VPWR_c_295_n 0.0471615f $X=1.085 $Y=2.15 $X2=0 $Y2=0
cc_104 N_B_c_85_n N_VGND_c_355_n 0.00166757f $X=0.95 $Y=0.76 $X2=0 $Y2=0
cc_105 N_B_c_86_n N_VGND_c_355_n 4.40092e-19 $X=0.95 $Y=0.91 $X2=0 $Y2=0
cc_106 N_B_c_85_n N_VGND_c_361_n 0.00403348f $X=0.95 $Y=0.76 $X2=0 $Y2=0
cc_107 N_B_c_85_n N_VGND_c_362_n 5.92419e-19 $X=0.95 $Y=0.76 $X2=0 $Y2=0
cc_108 N_B_c_85_n N_VGND_c_363_n 0.00564418f $X=0.95 $Y=0.76 $X2=0 $Y2=0
cc_109 N_A_M1002_g N_A_30_53#_c_179_n 0.0131287f $X=1.475 $Y=0.475 $X2=0 $Y2=0
cc_110 N_A_c_128_n N_A_30_53#_c_189_n 0.0113704f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_130_n N_A_30_53#_c_182_n 0.0184543f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_c_131_n N_A_30_53#_c_182_n 0.0261429f $X=0.717 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_c_128_n N_A_30_53#_c_192_n 2.12882e-19 $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_c_130_n N_A_30_53#_c_192_n 0.0103904f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_c_131_n N_A_30_53#_c_192_n 0.0163964f $X=0.717 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_c_128_n N_A_30_53#_c_184_n 0.0034911f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_M1002_g N_A_30_53#_c_184_n 0.0122277f $X=1.475 $Y=0.475 $X2=0 $Y2=0
cc_118 N_A_c_130_n N_A_30_53#_c_184_n 0.0204446f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_c_128_n N_A_30_53#_c_212_n 0.0153527f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_130_n N_A_30_53#_c_212_n 0.013641f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_M1002_g N_A_30_53#_c_185_n 0.00331117f $X=1.475 $Y=0.475 $X2=0 $Y2=0
cc_122 N_A_c_128_n N_A_30_53#_c_194_n 0.00334226f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_c_128_n N_A_30_53#_c_186_n 5.77159e-19 $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_130_n N_A_30_53#_c_186_n 0.0146254f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_c_128_n N_A_30_53#_c_195_n 0.0148587f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_130_n N_A_30_53#_c_195_n 0.011315f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_c_131_n N_A_30_53#_c_195_n 0.00544382f $X=0.717 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_c_128_n N_A_30_53#_c_187_n 0.00285728f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_130_n N_A_30_53#_c_187_n 0.0179327f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_c_128_n N_A_30_53#_c_188_n 0.00800977f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_c_130_n N_A_30_53#_c_188_n 3.08235e-19 $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_c_131_n A_120_297# 0.00128322f $X=0.717 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_133 N_A_c_128_n N_VPWR_c_296_n 0.00404913f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_128_n N_VPWR_c_299_n 0.00351268f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_128_n N_VPWR_c_295_n 0.00445321f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_M1002_g N_VGND_c_361_n 0.00187556f $X=1.475 $Y=0.475 $X2=0 $Y2=0
cc_137 N_A_M1002_g N_VGND_c_362_n 0.0107242f $X=1.475 $Y=0.475 $X2=0 $Y2=0
cc_138 N_A_M1002_g N_VGND_c_363_n 0.00260008f $X=1.475 $Y=0.475 $X2=0 $Y2=0
cc_139 N_A_30_53#_c_192_n A_120_297# 0.0012331f $X=1.2 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_140 N_A_30_53#_c_192_n A_202_297# 0.00258448f $X=1.2 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A_30_53#_c_195_n A_202_297# 0.00463716f $X=1.285 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_142 N_A_30_53#_c_212_n N_VPWR_M1006_d 0.0121405f $X=1.89 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_143 N_A_30_53#_c_189_n N_VPWR_c_296_n 0.0159668f $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_30_53#_c_212_n N_VPWR_c_296_n 0.0356988f $X=1.89 $Y=1.58 $X2=0 $Y2=0
cc_145 N_A_30_53#_c_195_n N_VPWR_c_296_n 0.00733636f $X=1.285 $Y=1.58 $X2=0
+ $Y2=0
cc_146 N_A_30_53#_c_190_n N_VPWR_c_298_n 0.00880278f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_30_53#_c_189_n N_VPWR_c_300_n 0.00702461f $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_30_53#_c_190_n N_VPWR_c_300_n 0.00559759f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_30_53#_c_189_n N_VPWR_c_295_n 0.0138964f $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_30_53#_c_190_n N_VPWR_c_295_n 0.0101476f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_30_53#_c_180_n N_X_c_328_n 0.00536146f $X=2.675 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_30_53#_c_184_n N_X_c_328_n 0.00703906f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_30_53#_c_188_n N_X_c_328_n 0.00549901f $X=2.65 $Y=1.202 $X2=0 $Y2=0
cc_154 N_A_30_53#_c_189_n N_X_c_331_n 0.00855852f $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_30_53#_c_190_n N_X_c_331_n 0.00408912f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_30_53#_c_212_n N_X_c_331_n 0.0114273f $X=1.89 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A_30_53#_c_188_n N_X_c_331_n 0.00617734f $X=2.65 $Y=1.202 $X2=0 $Y2=0
cc_158 N_A_30_53#_c_179_n N_X_c_326_n 0.00168199f $X=2.155 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_30_53#_c_189_n N_X_c_326_n 6.3219e-19 $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_30_53#_c_190_n N_X_c_326_n 0.00242981f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_30_53#_c_180_n N_X_c_326_n 0.00755759f $X=2.675 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_30_53#_c_184_n N_X_c_326_n 0.00287475f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_30_53#_c_185_n N_X_c_326_n 0.00700628f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_30_53#_c_194_n N_X_c_326_n 0.0070569f $X=2 $Y=1.495 $X2=0 $Y2=0
cc_165 N_A_30_53#_c_187_n N_X_c_326_n 0.024108f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_30_53#_c_188_n N_X_c_326_n 0.0308696f $X=2.65 $Y=1.202 $X2=0 $Y2=0
cc_167 N_A_30_53#_c_190_n X 0.0146614f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_30_53#_c_182_n N_VGND_M1008_d 0.00211434f $X=1.13 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_30_53#_c_184_n N_VGND_M1002_d 0.0111346f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_30_53#_c_185_n N_VGND_M1002_d 8.40753e-19 $X=2 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_30_53#_c_181_n N_VGND_c_355_n 0.0138472f $X=0.275 $Y=0.47 $X2=0 $Y2=0
cc_172 N_A_30_53#_c_182_n N_VGND_c_355_n 0.0214496f $X=1.13 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A_30_53#_c_180_n N_VGND_c_357_n 0.0103005f $X=2.675 $Y=0.995 $X2=0
+ $Y2=0
cc_174 N_A_30_53#_c_181_n N_VGND_c_358_n 0.0132481f $X=0.275 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A_30_53#_c_182_n N_VGND_c_358_n 0.0023206f $X=1.13 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_30_53#_c_179_n N_VGND_c_359_n 0.00524631f $X=2.155 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_30_53#_c_180_n N_VGND_c_359_n 0.00513402f $X=2.675 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_30_53#_c_184_n N_VGND_c_359_n 3.19125e-19 $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_30_53#_c_182_n N_VGND_c_361_n 0.0029785f $X=1.13 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A_30_53#_c_279_p N_VGND_c_361_n 0.00861358f $X=1.215 $Y=0.47 $X2=0
+ $Y2=0
cc_181 N_A_30_53#_c_184_n N_VGND_c_361_n 0.0023206f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_30_53#_c_179_n N_VGND_c_362_n 0.0143944f $X=2.155 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_30_53#_c_180_n N_VGND_c_362_n 0.00168957f $X=2.675 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_30_53#_c_279_p N_VGND_c_362_n 0.0139639f $X=1.215 $Y=0.47 $X2=0 $Y2=0
cc_185 N_A_30_53#_c_184_n N_VGND_c_362_n 0.0386993f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A_30_53#_c_179_n N_VGND_c_363_n 0.00874751f $X=2.155 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_30_53#_c_180_n N_VGND_c_363_n 0.0099569f $X=2.675 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_30_53#_c_181_n N_VGND_c_363_n 0.00942308f $X=0.275 $Y=0.47 $X2=0
+ $Y2=0
cc_189 N_A_30_53#_c_182_n N_VGND_c_363_n 0.011414f $X=1.13 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_30_53#_c_279_p N_VGND_c_363_n 0.00625722f $X=1.215 $Y=0.47 $X2=0
+ $Y2=0
cc_191 N_A_30_53#_c_184_n N_VGND_c_363_n 0.00753365f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_192 N_VPWR_c_295_n N_X_M1003_s 0.00444633f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_298_n N_X_c_326_n 0.0792653f $X=2.91 $Y=1.62 $X2=0 $Y2=0
cc_194 N_VPWR_c_300_n X 0.0205265f $X=2.825 $Y=2.72 $X2=0 $Y2=0
cc_195 N_VPWR_c_295_n X 0.0120094f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_196 N_VPWR_c_298_n N_VGND_c_357_n 0.0124587f $X=2.91 $Y=1.62 $X2=0 $Y2=0
cc_197 N_X_c_328_n N_VGND_c_357_n 0.026465f $X=2.562 $Y=0.587 $X2=0 $Y2=0
cc_198 N_X_c_326_n N_VGND_c_357_n 0.0114629f $X=2.492 $Y=1.495 $X2=0 $Y2=0
cc_199 N_X_c_328_n N_VGND_c_359_n 0.00969563f $X=2.562 $Y=0.587 $X2=0 $Y2=0
cc_200 N_X_c_328_n N_VGND_c_362_n 0.00427264f $X=2.562 $Y=0.587 $X2=0 $Y2=0
cc_201 N_X_M1000_s N_VGND_c_363_n 0.00668317f $X=2.23 $Y=0.235 $X2=0 $Y2=0
cc_202 N_X_c_328_n N_VGND_c_363_n 0.0108492f $X=2.562 $Y=0.587 $X2=0 $Y2=0
