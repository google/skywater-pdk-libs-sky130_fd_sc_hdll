* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VGND A1_N a_343_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_341_297# A2_N a_343_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X2 a_82_21# B2 a_696_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_82_21# a_343_47# a_622_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X4 VGND a_343_47# a_82_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VPWR B1 a_622_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X7 a_622_369# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X8 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_696_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_343_47# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR A1_N a_341_297# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X13 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
