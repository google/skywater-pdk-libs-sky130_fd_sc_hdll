* File: sky130_fd_sc_hdll__and2_2.pex.spice
* Created: Thu Aug 27 18:56:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND2_2%A 2 3 5 8 12 13 15 16 22 24
r37 22 24 8.36086 $w=2.53e-07 $l=1.85e-07 $layer=LI1_cond $X=0.222 $Y=1.325
+ $X2=0.222 $Y2=1.51
r38 16 24 1.80775 $w=2.53e-07 $l=4e-08 $layer=LI1_cond $X=0.222 $Y=1.55
+ $X2=0.222 $Y2=1.51
r39 15 22 3.36826 $w=2.55e-07 $l=1.25e-07 $layer=LI1_cond $X=0.222 $Y=1.2
+ $X2=0.222 $Y2=1.325
r40 13 21 37.7137 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.44 $Y=1.16
+ $X2=0.44 $Y2=1.325
r41 13 20 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.44 $Y=1.16
+ $X2=0.44 $Y2=0.995
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.45
+ $Y=1.16 $X2=0.45 $Y2=1.16
r43 10 15 3.4491 $w=2.5e-07 $l=1.28e-07 $layer=LI1_cond $X=0.35 $Y=1.2 $X2=0.222
+ $Y2=1.2
r44 10 12 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=0.35 $Y=1.2 $X2=0.45
+ $Y2=1.2
r45 8 20 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.54 $Y=0.585
+ $X2=0.54 $Y2=0.995
r46 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.515 $Y=1.78
+ $X2=0.515 $Y2=2.065
r47 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.515 $Y=1.68 $X2=0.515
+ $Y2=1.78
r48 2 21 117.71 $w=2e-07 $l=3.55e-07 $layer=POLY_cond $X=0.515 $Y=1.68 $X2=0.515
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_2%B 3 6 7 9 10 13
r41 13 16 36.565 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.16
+ $X2=1.075 $Y2=1.325
r42 13 15 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.16
+ $X2=1.075 $Y2=0.995
r43 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.16 $X2=1.05 $Y2=1.16
r44 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.985 $Y=1.78
+ $X2=0.985 $Y2=2.065
r45 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.985 $Y=1.68 $X2=0.985
+ $Y2=1.78
r46 6 16 117.71 $w=2e-07 $l=3.55e-07 $layer=POLY_cond $X=0.985 $Y=1.68 $X2=0.985
+ $Y2=1.325
r47 3 15 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.96 $Y=0.585
+ $X2=0.96 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_2%A_27_75# 1 2 7 9 10 12 13 15 17 18 20 21 24
+ 26 27 30 32 33 34 35 39
r98 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.64
+ $Y=1.16 $X2=1.64 $Y2=1.16
r99 36 38 16.6797 $w=2.56e-07 $l=3.5e-07 $layer=LI1_cond $X=1.6 $Y=0.81 $X2=1.6
+ $Y2=1.16
r100 34 38 9.24244 $w=2.56e-07 $l=2.0106e-07 $layer=LI1_cond $X=1.52 $Y=1.325
+ $X2=1.6 $Y2=1.16
r101 34 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.52 $Y=1.325
+ $X2=1.52 $Y2=1.575
r102 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=1.66
+ $X2=1.52 $Y2=1.575
r103 32 33 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.435 $Y=1.66
+ $X2=0.915 $Y2=1.66
r104 28 33 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.765 $Y=1.745
+ $X2=0.915 $Y2=1.66
r105 28 30 14.7897 $w=2.98e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=1.745
+ $X2=0.765 $Y2=2.13
r106 26 36 2.48511 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.81
+ $X2=1.6 $Y2=0.81
r107 26 27 57.7895 $w=1.88e-07 $l=9.9e-07 $layer=LI1_cond $X=1.435 $Y=0.81
+ $X2=0.445 $Y2=0.81
r108 22 27 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.28 $Y=0.715
+ $X2=0.445 $Y2=0.81
r109 22 24 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.28 $Y=0.715
+ $X2=0.28 $Y2=0.52
r110 18 21 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=2.19 $Y=0.995
+ $X2=2.165 $Y2=1.202
r111 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.19 $Y=0.995
+ $X2=2.19 $Y2=0.56
r112 15 21 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=2.165 $Y=1.41
+ $X2=2.165 $Y2=1.202
r113 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.165 $Y=1.41
+ $X2=2.165 $Y2=1.985
r114 14 39 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.675 $Y=1.16
+ $X2=1.575 $Y2=1.202
r115 13 21 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.065 $Y=1.16
+ $X2=2.165 $Y2=1.202
r116 13 14 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=2.065 $Y=1.16
+ $X2=1.675 $Y2=1.16
r117 10 39 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.575 $Y=1.41
+ $X2=1.575 $Y2=1.202
r118 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.575 $Y=1.41
+ $X2=1.575 $Y2=1.985
r119 7 39 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.55 $Y=0.995
+ $X2=1.575 $Y2=1.202
r120 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.55 $Y=0.995
+ $X2=1.55 $Y2=0.56
r121 2 30 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.855 $X2=0.75 $Y2=2.13
r122 1 24 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.375 $X2=0.28 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_2%VPWR 1 2 3 10 12 16 18 20 25 26 27 33 42
r38 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r40 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 33 41 4.40761 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.567 $Y2=2.72
r42 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 32 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r45 29 38 4.27358 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r46 29 31 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 27 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 27 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r49 25 31 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 25 26 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.335 $Y2=2.72
r51 24 35 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.505 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 24 26 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.505 $Y=2.72
+ $X2=1.335 $Y2=2.72
r53 20 23 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=2.52 $Y=1.66
+ $X2=2.52 $Y2=2.34
r54 18 41 3.03023 $w=2.9e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.52 $Y=2.635
+ $X2=2.567 $Y2=2.72
r55 18 23 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.52 $Y=2.635
+ $X2=2.52 $Y2=2.34
r56 14 26 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=2.635
+ $X2=1.335 $Y2=2.72
r57 14 16 21.5236 $w=3.38e-07 $l=6.35e-07 $layer=LI1_cond $X=1.335 $Y=2.635
+ $X2=1.335 $Y2=2
r58 10 38 3.08647 $w=2.8e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.197 $Y2=2.72
r59 10 12 20.7851 $w=2.78e-07 $l=5.05e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.255 $Y2=2.13
r60 3 23 400 $w=1.7e-07 $l=9.51998e-07 $layer=licon1_PDIFF $count=1 $X=2.255
+ $Y=1.485 $X2=2.46 $Y2=2.34
r61 3 20 400 $w=1.7e-07 $l=2.79106e-07 $layer=licon1_PDIFF $count=1 $X=2.255
+ $Y=1.485 $X2=2.46 $Y2=1.66
r62 2 16 300 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.855 $X2=1.34 $Y2=2
r63 1 12 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.855 $X2=0.28 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_2%X 1 2 7 11 12 13 14 15 16 25 36
r32 36 40 1.92074 $w=2.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.07 $Y=1.87
+ $X2=2.07 $Y2=1.915
r33 16 42 5.46036 $w=4.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.975 $Y=2.21
+ $X2=1.975 $Y2=2
r34 15 42 1.69011 $w=4.58e-07 $l=6.5e-08 $layer=LI1_cond $X=1.975 $Y=1.935
+ $X2=1.975 $Y2=2
r35 15 40 2.54368 $w=4.58e-07 $l=2e-08 $layer=LI1_cond $X=1.975 $Y=1.935
+ $X2=1.975 $Y2=1.915
r36 15 36 0.853661 $w=2.68e-07 $l=2e-08 $layer=LI1_cond $X=2.07 $Y=1.85 $X2=2.07
+ $Y2=1.87
r37 14 15 13.6586 $w=2.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.07 $Y=1.53
+ $X2=2.07 $Y2=1.85
r38 13 14 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.07 $Y=1.19
+ $X2=2.07 $Y2=1.53
r39 12 13 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.07 $Y=0.85
+ $X2=2.07 $Y2=1.19
r40 11 25 3.53583 $w=2.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.07 $Y=0.4 $X2=2.07
+ $Y2=0.545
r41 11 12 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.07 $Y=0.57
+ $X2=2.07 $Y2=0.85
r42 11 25 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.07 $Y=0.57
+ $X2=2.07 $Y2=0.545
r43 7 11 3.29198 $w=2.9e-07 $l=1.35e-07 $layer=LI1_cond $X=1.935 $Y=0.4 $X2=2.07
+ $Y2=0.4
r44 7 9 4.96743 $w=2.88e-07 $l=1.25e-07 $layer=LI1_cond $X=1.935 $Y=0.4 $X2=1.81
+ $Y2=0.4
r45 2 42 300 $w=1.7e-07 $l=6.2562e-07 $layer=licon1_PDIFF $count=2 $X=1.665
+ $Y=1.485 $X2=1.91 $Y2=2
r46 1 9 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.235 $X2=1.81 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_2%VGND 1 2 9 11 13 16 17 18 27 33
r34 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r35 30 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r36 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r37 27 32 4.40761 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.567
+ $Y2=0
r38 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.07
+ $Y2=0
r39 26 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r40 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r41 21 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r42 18 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r43 18 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r44 16 25 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.15
+ $Y2=0
r45 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.3
+ $Y2=0
r46 15 29 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=2.07
+ $Y2=0
r47 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.3
+ $Y2=0
r48 11 32 3.03023 $w=2.9e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.52 $Y=0.085
+ $X2=2.567 $Y2=0
r49 11 13 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.52 $Y=0.085
+ $X2=2.52 $Y2=0.38
r50 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=0.085
+ $X2=1.3 $Y2=0
r51 7 9 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.3 $Y=0.085 $X2=1.3
+ $Y2=0.38
r52 2 13 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=2.265
+ $Y=0.235 $X2=2.46 $Y2=0.38
r53 1 9 182 $w=1.7e-07 $l=3.0749e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.375 $X2=1.34 $Y2=0.38
.ends

