* File: sky130_fd_sc_hdll__and4_4.pex.spice
* Created: Wed Sep  2 08:23:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND4_4%A 1 3 4 6 7 8 14
r29 14 15 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r30 12 14 33.0137 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.202
+ $X2=0.495 $Y2=1.202
r31 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r32 7 8 16.7716 $w=2.03e-07 $l=3.1e-07 $layer=LI1_cond $X=0.227 $Y=0.85
+ $X2=0.227 $Y2=1.16
r33 4 15 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r35 1 14 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_4%B 1 3 4 6 7 8 9
r31 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.16 $X2=0.975 $Y2=1.16
r32 9 15 0.788623 $w=4.53e-07 $l=3e-08 $layer=LI1_cond $X=1.117 $Y=1.19
+ $X2=1.117 $Y2=1.16
r33 8 15 8.14911 $w=4.53e-07 $l=3.1e-07 $layer=LI1_cond $X=1.117 $Y=0.85
+ $X2=1.117 $Y2=1.16
r34 7 8 8.93773 $w=4.53e-07 $l=3.4e-07 $layer=LI1_cond $X=1.117 $Y=0.51
+ $X2=1.117 $Y2=0.85
r35 4 14 48.1839 $w=2.94e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=1 $Y2=1.16
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r37 1 14 38.5845 $w=2.94e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.915 $Y=0.995
+ $X2=1 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.915 $Y=0.995
+ $X2=0.915 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_4%C 1 3 4 6 7 8 9
r31 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6 $Y=1.16
+ $X2=1.6 $Y2=1.16
r32 8 9 13.4814 $w=2.63e-07 $l=3.1e-07 $layer=LI1_cond $X=1.647 $Y=0.85
+ $X2=1.647 $Y2=1.16
r33 7 8 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=1.647 $Y=0.51
+ $X2=1.647 $Y2=0.85
r34 4 14 45.3064 $w=3.7e-07 $l=2.96648e-07 $layer=POLY_cond $X=1.475 $Y=1.41
+ $X2=1.577 $Y2=1.16
r35 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.475 $Y=1.41
+ $X2=1.475 $Y2=1.985
r36 1 14 39.0558 $w=3.7e-07 $l=2.21371e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.577 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.445 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_4%D 1 3 4 6 7
r37 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.16 $X2=2.14 $Y2=1.16
r38 7 11 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=2.13 $Y=0.85 $X2=2.13
+ $Y2=1.16
r39 4 10 47.9974 $w=2.97e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.165 $Y2=1.16
r40 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.105 $Y2=1.985
r41 1 10 43.4349 $w=2.97e-07 $l=2.33666e-07 $layer=POLY_cond $X=2.08 $Y=0.965
+ $X2=2.165 $Y2=1.16
r42 1 3 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.08 $Y=0.965 $X2=2.08
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_4%A_27_47# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 35 38 40 44 46 49 50 55 61 63 64 73
c134 49 0 1.10875e-19 $X=2.53 $Y=1.495
r135 73 74 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.045 $Y=1.202
+ $X2=4.07 $Y2=1.202
r136 70 71 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.55 $Y=1.202
+ $X2=3.575 $Y2=1.202
r137 69 70 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=3.105 $Y=1.202
+ $X2=3.55 $Y2=1.202
r138 68 69 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.08 $Y=1.202
+ $X2=3.105 $Y2=1.202
r139 65 66 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.61 $Y=1.202
+ $X2=2.635 $Y2=1.202
r140 59 61 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.26 $Y=0.42
+ $X2=0.61 $Y2=0.42
r141 56 73 35.6317 $w=3.72e-07 $l=2.75e-07 $layer=POLY_cond $X=3.77 $Y=1.202
+ $X2=4.045 $Y2=1.202
r142 56 71 25.2661 $w=3.72e-07 $l=1.95e-07 $layer=POLY_cond $X=3.77 $Y=1.202
+ $X2=3.575 $Y2=1.202
r143 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.77
+ $Y=1.16 $X2=3.77 $Y2=1.16
r144 53 68 11.6613 $w=3.72e-07 $l=9e-08 $layer=POLY_cond $X=2.99 $Y=1.202
+ $X2=3.08 $Y2=1.202
r145 53 66 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=2.99 $Y=1.202
+ $X2=2.635 $Y2=1.202
r146 52 55 39.0829 $w=2.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.99 $Y=1.19
+ $X2=3.77 $Y2=1.19
r147 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.16 $X2=2.99 $Y2=1.16
r148 50 52 18.7898 $w=2.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.615 $Y=1.19
+ $X2=2.99 $Y2=1.19
r149 48 50 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.53 $Y=1.305
+ $X2=2.615 $Y2=1.19
r150 48 49 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.53 $Y=1.305
+ $X2=2.53 $Y2=1.495
r151 47 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.795 $Y=1.58
+ $X2=1.7 $Y2=1.58
r152 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=2.53 $Y2=1.495
r153 46 47 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=1.795 $Y2=1.58
r154 42 64 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=1.665
+ $X2=1.7 $Y2=1.58
r155 42 44 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.7 $Y=1.665
+ $X2=1.7 $Y2=1.96
r156 41 63 2.20034 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.815 $Y=1.58
+ $X2=0.657 $Y2=1.58
r157 40 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.605 $Y=1.58
+ $X2=1.7 $Y2=1.58
r158 40 41 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.605 $Y=1.58
+ $X2=0.815 $Y2=1.58
r159 36 63 4.23118 $w=2.15e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.71 $Y=1.665
+ $X2=0.657 $Y2=1.58
r160 36 38 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.71 $Y=1.665
+ $X2=0.71 $Y2=1.96
r161 35 63 4.23118 $w=2.15e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.61 $Y=1.495
+ $X2=0.657 $Y2=1.58
r162 34 61 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=0.585
+ $X2=0.61 $Y2=0.42
r163 34 35 47.6692 $w=2.18e-07 $l=9.1e-07 $layer=LI1_cond $X=0.61 $Y=0.585
+ $X2=0.61 $Y2=1.495
r164 31 74 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.07 $Y=0.995
+ $X2=4.07 $Y2=1.202
r165 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.07 $Y=0.995
+ $X2=4.07 $Y2=0.56
r166 28 73 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.045 $Y=1.41
+ $X2=4.045 $Y2=1.202
r167 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.045 $Y=1.41
+ $X2=4.045 $Y2=1.985
r168 25 71 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.575 $Y=1.41
+ $X2=3.575 $Y2=1.202
r169 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.575 $Y=1.41
+ $X2=3.575 $Y2=1.985
r170 22 70 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.55 $Y=0.995
+ $X2=3.55 $Y2=1.202
r171 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.55 $Y=0.995
+ $X2=3.55 $Y2=0.56
r172 19 69 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.105 $Y=1.41
+ $X2=3.105 $Y2=1.202
r173 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.105 $Y=1.41
+ $X2=3.105 $Y2=1.985
r174 16 68 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.08 $Y=0.995
+ $X2=3.08 $Y2=1.202
r175 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.08 $Y=0.995
+ $X2=3.08 $Y2=0.56
r176 13 66 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.635 $Y=1.41
+ $X2=2.635 $Y2=1.202
r177 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.635 $Y=1.41
+ $X2=2.635 $Y2=1.985
r178 10 65 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.61 $Y=0.995
+ $X2=2.61 $Y2=1.202
r179 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.61 $Y=0.995
+ $X2=2.61 $Y2=0.56
r180 3 44 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.565
+ $Y=1.485 $X2=1.71 $Y2=1.96
r181 2 38 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
r182 1 59 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_4%VPWR 1 2 3 4 5 16 18 22 26 30 32 34 37 38
+ 40 41 42 44 56 64 68
c73 3 0 1.10875e-19 $X=2.195 $Y=1.485
r74 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r75 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r76 59 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r77 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r78 56 67 5.10144 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=4.332 $Y2=2.72
r79 56 58 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=3.91 $Y2=2.72
r80 55 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r81 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r82 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 52 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r84 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r85 49 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=2.72
+ $X2=1.22 $Y2=2.72
r86 49 51 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.385 $Y=2.72
+ $X2=2.07 $Y2=2.72
r87 48 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r88 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 45 61 4.29151 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r90 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r91 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=1.22 $Y2=2.72
r92 44 47 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=0.69 $Y2=2.72
r93 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 42 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 40 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=2.72
+ $X2=2.99 $Y2=2.72
r96 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.255 $Y=2.72
+ $X2=3.38 $Y2=2.72
r97 39 58 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.505 $Y=2.72
+ $X2=3.91 $Y2=2.72
r98 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.505 $Y=2.72
+ $X2=3.38 $Y2=2.72
r99 37 51 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.07 $Y2=2.72
r100 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.39 $Y2=2.72
r101 36 54 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.555 $Y=2.72
+ $X2=2.99 $Y2=2.72
r102 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.555 $Y=2.72
+ $X2=2.39 $Y2=2.72
r103 32 67 3.09525 $w=3.8e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.255 $Y=2.635
+ $X2=4.332 $Y2=2.72
r104 32 34 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=4.255 $Y=2.635
+ $X2=4.255 $Y2=2
r105 28 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.38 $Y=2.635
+ $X2=3.38 $Y2=2.72
r106 28 30 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.38 $Y=2.635
+ $X2=3.38 $Y2=2
r107 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=2.635
+ $X2=2.39 $Y2=2.72
r108 24 26 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.39 $Y=2.635
+ $X2=2.39 $Y2=2.02
r109 20 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=2.72
r110 20 22 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=2.02
r111 16 61 3.06854 $w=2.8e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.192 $Y2=2.72
r112 16 18 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.245 $Y2=2
r113 5 34 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.135
+ $Y=1.485 $X2=4.28 $Y2=2
r114 4 30 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.195
+ $Y=1.485 $X2=3.34 $Y2=2
r115 3 26 300 $w=1.7e-07 $l=6.2494e-07 $layer=licon1_PDIFF $count=2 $X=2.195
+ $Y=1.485 $X2=2.39 $Y2=2.02
r116 2 22 300 $w=1.7e-07 $l=6.11964e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.22 $Y2=2.02
r117 1 18 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_4%X 1 2 3 4 15 19 21 22 23 24 27 31 33 35 37
+ 38 39 40 41 47 48 50
r83 47 50 1.80775 $w=2.53e-07 $l=4e-08 $layer=LI1_cond $X=4.327 $Y=0.81
+ $X2=4.327 $Y2=0.85
r84 41 48 3.44845 $w=2.55e-07 $l=1.3e-07 $layer=LI1_cond $X=4.327 $Y=1.615
+ $X2=4.327 $Y2=1.485
r85 41 48 0.903877 $w=2.53e-07 $l=2e-08 $layer=LI1_cond $X=4.327 $Y=1.465
+ $X2=4.327 $Y2=1.485
r86 40 41 12.4283 $w=2.53e-07 $l=2.75e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.327 $Y2=1.465
r87 39 47 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.327 $Y=0.725
+ $X2=4.327 $Y2=0.81
r88 39 40 14.3716 $w=2.53e-07 $l=3.18e-07 $layer=LI1_cond $X=4.327 $Y=0.872
+ $X2=4.327 $Y2=1.19
r89 39 50 0.994265 $w=2.53e-07 $l=2.2e-08 $layer=LI1_cond $X=4.327 $Y=0.872
+ $X2=4.327 $Y2=0.85
r90 36 38 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=1.615
+ $X2=3.81 $Y2=1.615
r91 35 41 3.36887 $w=2.6e-07 $l=1.27e-07 $layer=LI1_cond $X=4.2 $Y=1.615
+ $X2=4.327 $Y2=1.615
r92 35 36 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=4.2 $Y=1.615
+ $X2=3.895 $Y2=1.615
r93 34 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=0.725
+ $X2=3.81 $Y2=0.725
r94 33 39 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.2 $Y=0.725
+ $X2=4.327 $Y2=0.725
r95 33 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.2 $Y=0.725
+ $X2=3.895 $Y2=0.725
r96 29 38 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.81 $Y=1.745
+ $X2=3.81 $Y2=1.615
r97 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.81 $Y=1.745
+ $X2=3.81 $Y2=1.96
r98 25 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=0.64 $X2=3.81
+ $Y2=0.725
r99 25 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.81 $Y=0.64
+ $X2=3.81 $Y2=0.42
r100 23 38 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.725 $Y=1.57
+ $X2=3.81 $Y2=1.615
r101 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.725 $Y=1.57
+ $X2=3.035 $Y2=1.57
r102 21 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0.725
+ $X2=3.81 $Y2=0.725
r103 21 22 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.725 $Y=0.725
+ $X2=2.955 $Y2=0.725
r104 17 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.91 $Y=1.655
+ $X2=3.035 $Y2=1.57
r105 17 19 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=2.91 $Y=1.655
+ $X2=2.91 $Y2=1.96
r106 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.87 $Y=0.64
+ $X2=2.955 $Y2=0.725
r107 13 15 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.87 $Y=0.64
+ $X2=2.87 $Y2=0.42
r108 4 31 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.665
+ $Y=1.485 $X2=3.81 $Y2=1.96
r109 3 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.725
+ $Y=1.485 $X2=2.87 $Y2=1.96
r110 2 27 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=3.625
+ $Y=0.235 $X2=3.81 $Y2=0.42
r111 1 15 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=2.685
+ $Y=0.235 $X2=2.87 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4_4%VGND 1 2 3 12 16 18 20 23 24 26 27 28 40 46
r74 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r75 43 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r76 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r77 40 45 5.10144 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=4.065 $Y=0 $X2=4.332
+ $Y2=0
r78 40 42 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.065 $Y=0 $X2=3.91
+ $Y2=0
r79 39 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r80 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r81 36 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r82 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r83 31 35 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r84 28 36 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r85 28 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r86 26 38 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=2.99
+ $Y2=0
r87 26 27 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.315
+ $Y2=0
r88 25 42 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.91
+ $Y2=0
r89 25 27 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.315
+ $Y2=0
r90 23 35 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.07
+ $Y2=0
r91 23 24 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.38
+ $Y2=0
r92 22 38 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.99
+ $Y2=0
r93 22 24 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.38
+ $Y2=0
r94 18 45 3.09525 $w=3.8e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.332 $Y2=0
r95 18 20 9.09823 $w=3.78e-07 $l=3e-07 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0.385
r96 14 27 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0
r97 14 16 9.09823 $w=3.78e-07 $l=3e-07 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0.385
r98 10 24 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=0.085
+ $X2=2.38 $Y2=0
r99 10 12 11.1527 $w=3.08e-07 $l=3e-07 $layer=LI1_cond $X=2.38 $Y=0.085 $X2=2.38
+ $Y2=0.385
r100 3 20 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=4.145
+ $Y=0.235 $X2=4.28 $Y2=0.385
r101 2 16 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.235 $X2=3.34 $Y2=0.385
r102 1 12 182 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.235 $X2=2.39 $Y2=0.385
.ends

