* File: sky130_fd_sc_hdll__inv_6.spice
* Created: Thu Aug 27 19:09:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__inv_6.pex.spice"
.subckt sky130_fd_sc_hdll__inv_6  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75002.5
+ A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7 SB=75002.1
+ A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1005_d N_A_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1 SB=75001.6
+ A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_M1008_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6 SB=75001.1
+ A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1008_d N_A_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1 SB=75000.7
+ A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.65 AD=0.1755
+ AS=0.104 PD=1.84 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1002_d N_A_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1004_d N_A_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g N_Y_M1007_s VPB PHIGHVT L=0.18 W=1 AD=0.28
+ AS=0.145 PD=2.56 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX13_noxref noxref_7 A A PROBETYPE=1
pX14_noxref noxref_8 A A PROBETYPE=1
pX15_noxref noxref_9 A A PROBETYPE=1
*
.include "sky130_fd_sc_hdll__inv_6.pxi.spice"
*
.ends
*
*
