* NGSPICE file created from sky130_fd_sc_hdll__nor4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
M1000 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=4.034e+11p ps=3.96e+06u
M1001 VGND A Y VNB nshort w=650000u l=150000u
+  ad=1.1897e+12p pd=1.252e+07u as=9.295e+11p ps=8.06e+06u
M1002 VGND D_N a_754_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1003 Y a_754_21# a_514_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.3e+11p ps=7.66e+06u
M1004 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR D_N a_754_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1006 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_514_297# C a_305_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1008 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_305_297# C a_514_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# B a_305_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_754_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_305_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_754_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_514_297# a_754_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

