* File: sky130_fd_sc_hdll__buf_12.pex.spice
* Created: Thu Aug 27 18:59:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUF_12%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 49 54 56 59 62
c84 32 0 1.25463e-19 $X=1.52 $Y=1.105
r85 54 56 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.315 $Y=1.175
+ $X2=0.655 $Y2=1.175
r86 49 50 3.73065 $w=3.23e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.212
+ $X2=1.93 $Y2=1.212
r87 47 49 59.6904 $w=3.23e-07 $l=4e-07 $layer=POLY_cond $X=1.505 $Y=1.212
+ $X2=1.905 $Y2=1.212
r88 47 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.505
+ $Y=1.16 $X2=1.505 $Y2=1.16
r89 45 47 6.71517 $w=3.23e-07 $l=4.5e-08 $layer=POLY_cond $X=1.46 $Y=1.212
+ $X2=1.505 $Y2=1.212
r90 44 45 3.73065 $w=3.23e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.212
+ $X2=1.46 $Y2=1.212
r91 43 44 66.4056 $w=3.23e-07 $l=4.45e-07 $layer=POLY_cond $X=0.99 $Y=1.212
+ $X2=1.435 $Y2=1.212
r92 42 43 3.73065 $w=3.23e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.212
+ $X2=0.99 $Y2=1.212
r93 41 42 66.4056 $w=3.23e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.212
+ $X2=0.965 $Y2=1.212
r94 40 41 3.73065 $w=3.23e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.212
+ $X2=0.52 $Y2=1.212
r95 38 40 16.4149 $w=3.23e-07 $l=1.1e-07 $layer=POLY_cond $X=0.385 $Y=1.212
+ $X2=0.495 $Y2=1.212
r96 38 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.16 $X2=0.385 $Y2=1.16
r97 32 62 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=1.605 $Y=1.175
+ $X2=1.505 $Y2=1.175
r98 31 62 19.1318 $w=1.98e-07 $l=3.45e-07 $layer=LI1_cond $X=1.16 $Y=1.175
+ $X2=1.505 $Y2=1.175
r99 31 59 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=1.16 $Y=1.175
+ $X2=1.115 $Y2=1.175
r100 30 59 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=0.705 $Y=1.175
+ $X2=1.115 $Y2=1.175
r101 30 56 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=0.705 $Y=1.175
+ $X2=0.655 $Y2=1.175
r102 29 54 1.94091 $w=1.98e-07 $l=3.5e-08 $layer=LI1_cond $X=0.28 $Y=1.175
+ $X2=0.315 $Y2=1.175
r103 25 50 20.7134 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.212
r104 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r105 22 49 16.4327 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.212
r106 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r107 18 45 20.7134 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.212
r108 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r109 15 44 16.4327 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.212
r110 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r111 11 43 20.7134 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=1.212
r112 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=0.56
r113 8 42 16.4327 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.212
r114 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r115 4 41 20.7134 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=1.212
r116 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=0.56
r117 1 40 16.4327 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.212
r118 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_12%A_117_297# 1 2 3 4 15 17 19 22 24 26 29 31
+ 33 36 38 40 43 45 47 50 52 54 57 59 61 64 66 68 71 73 75 78 80 82 85 87 89 90
+ 92 95 99 105 107 108 109 110 113 119 121 123 126 128 134 137 138 139 164
c294 164 0 1.25463e-19 $X=7.545 $Y=1.217
r295 164 165 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=7.545 $Y=1.217
+ $X2=7.57 $Y2=1.217
r296 163 164 70.5732 $w=3.21e-07 $l=4.7e-07 $layer=POLY_cond $X=7.075 $Y=1.217
+ $X2=7.545 $Y2=1.217
r297 162 163 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=7.05 $Y=1.217
+ $X2=7.075 $Y2=1.217
r298 161 162 66.8193 $w=3.21e-07 $l=4.45e-07 $layer=POLY_cond $X=6.605 $Y=1.217
+ $X2=7.05 $Y2=1.217
r299 160 161 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=6.58 $Y=1.217
+ $X2=6.605 $Y2=1.217
r300 159 160 66.8193 $w=3.21e-07 $l=4.45e-07 $layer=POLY_cond $X=6.135 $Y=1.217
+ $X2=6.58 $Y2=1.217
r301 158 159 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=6.11 $Y=1.217
+ $X2=6.135 $Y2=1.217
r302 157 158 66.8193 $w=3.21e-07 $l=4.45e-07 $layer=POLY_cond $X=5.665 $Y=1.217
+ $X2=6.11 $Y2=1.217
r303 156 157 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=5.64 $Y=1.217
+ $X2=5.665 $Y2=1.217
r304 155 156 66.8193 $w=3.21e-07 $l=4.45e-07 $layer=POLY_cond $X=5.195 $Y=1.217
+ $X2=5.64 $Y2=1.217
r305 154 155 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.217
+ $X2=5.195 $Y2=1.217
r306 151 152 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.217
+ $X2=4.725 $Y2=1.217
r307 150 151 66.8193 $w=3.21e-07 $l=4.45e-07 $layer=POLY_cond $X=4.255 $Y=1.217
+ $X2=4.7 $Y2=1.217
r308 149 150 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.217
+ $X2=4.255 $Y2=1.217
r309 148 149 66.8193 $w=3.21e-07 $l=4.45e-07 $layer=POLY_cond $X=3.785 $Y=1.217
+ $X2=4.23 $Y2=1.217
r310 147 148 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.217
+ $X2=3.785 $Y2=1.217
r311 146 147 66.8193 $w=3.21e-07 $l=4.45e-07 $layer=POLY_cond $X=3.315 $Y=1.217
+ $X2=3.76 $Y2=1.217
r312 145 146 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.217
+ $X2=3.315 $Y2=1.217
r313 144 145 66.8193 $w=3.21e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=3.29 $Y2=1.217
r314 143 144 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.217
+ $X2=2.845 $Y2=1.217
r315 140 141 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r316 135 154 63.0654 $w=3.21e-07 $l=4.2e-07 $layer=POLY_cond $X=4.75 $Y=1.217
+ $X2=5.17 $Y2=1.217
r317 135 152 3.75389 $w=3.21e-07 $l=2.5e-08 $layer=POLY_cond $X=4.75 $Y=1.217
+ $X2=4.725 $Y2=1.217
r318 134 135 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=4.75
+ $Y=1.16 $X2=4.75 $Y2=1.16
r319 132 143 54.0561 $w=3.21e-07 $l=3.6e-07 $layer=POLY_cond $X=2.46 $Y=1.217
+ $X2=2.82 $Y2=1.217
r320 132 141 12.7632 $w=3.21e-07 $l=8.5e-08 $layer=POLY_cond $X=2.46 $Y=1.217
+ $X2=2.375 $Y2=1.217
r321 131 134 149.401 $w=1.68e-07 $l=2.29e-06 $layer=LI1_cond $X=2.46 $Y=1.16
+ $X2=4.75 $Y2=1.16
r322 131 132 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r323 129 139 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.215 $Y=1.16
+ $X2=2.127 $Y2=1.16
r324 129 131 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.215 $Y=1.16
+ $X2=2.46 $Y2=1.16
r325 127 139 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.127 $Y=1.245
+ $X2=2.127 $Y2=1.16
r326 127 128 12.6753 $w=1.73e-07 $l=2e-07 $layer=LI1_cond $X=2.127 $Y=1.245
+ $X2=2.127 $Y2=1.445
r327 126 139 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.127 $Y=1.075
+ $X2=2.127 $Y2=1.16
r328 125 126 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=2.127 $Y=0.905
+ $X2=2.127 $Y2=1.075
r329 124 137 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.53
+ $X2=1.645 $Y2=1.53
r330 123 128 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=2.04 $Y=1.53
+ $X2=2.127 $Y2=1.445
r331 123 124 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.04 $Y=1.53
+ $X2=1.835 $Y2=1.53
r332 122 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0.82
+ $X2=1.67 $Y2=0.82
r333 121 125 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=2.04 $Y=0.82
+ $X2=2.127 $Y2=0.905
r334 121 122 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.04 $Y=0.82
+ $X2=1.755 $Y2=0.82
r335 117 138 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.735
+ $X2=1.67 $Y2=0.82
r336 117 119 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.67 $Y=0.735
+ $X2=1.67 $Y2=0.56
r337 113 115 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.645 $Y=1.63
+ $X2=1.645 $Y2=2.31
r338 111 137 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=1.615
+ $X2=1.645 $Y2=1.53
r339 111 113 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.645 $Y=1.615
+ $X2=1.645 $Y2=1.63
r340 109 137 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.53
+ $X2=1.645 $Y2=1.53
r341 109 110 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.53
+ $X2=0.895 $Y2=1.53
r342 107 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0.82
+ $X2=1.67 $Y2=0.82
r343 107 108 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0.82
+ $X2=0.815 $Y2=0.82
r344 103 108 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.73 $Y=0.735
+ $X2=0.815 $Y2=0.82
r345 103 105 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.73 $Y=0.735
+ $X2=0.73 $Y2=0.56
r346 99 101 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.705 $Y=1.63
+ $X2=0.705 $Y2=2.31
r347 97 110 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=0.705 $Y=1.615
+ $X2=0.895 $Y2=1.53
r348 97 99 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=0.705 $Y=1.615
+ $X2=0.705 $Y2=1.63
r349 93 165 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.57 $Y=1.025
+ $X2=7.57 $Y2=1.217
r350 93 95 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.57 $Y=1.025
+ $X2=7.57 $Y2=0.56
r351 90 164 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.217
r352 90 92 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.985
r353 87 163 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.217
r354 87 89 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.985
r355 83 162 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.05 $Y=1.025
+ $X2=7.05 $Y2=1.217
r356 83 85 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.05 $Y=1.025
+ $X2=7.05 $Y2=0.56
r357 80 161 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.217
r358 80 82 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.985
r359 76 160 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.58 $Y=1.025
+ $X2=6.58 $Y2=1.217
r360 76 78 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.58 $Y=1.025
+ $X2=6.58 $Y2=0.56
r361 73 159 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.217
r362 73 75 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.985
r363 69 158 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.11 $Y=1.025
+ $X2=6.11 $Y2=1.217
r364 69 71 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.11 $Y=1.025
+ $X2=6.11 $Y2=0.56
r365 66 157 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.217
r366 66 68 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r367 62 156 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.64 $Y=1.025
+ $X2=5.64 $Y2=1.217
r368 62 64 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.64 $Y=1.025
+ $X2=5.64 $Y2=0.56
r369 59 155 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.217
r370 59 61 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r371 55 154 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=1.217
r372 55 57 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=0.56
r373 52 152 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.217
r374 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r375 48 151 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=1.217
r376 48 50 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=0.56
r377 45 150 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.217
r378 45 47 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r379 41 149 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=1.217
r380 41 43 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=0.56
r381 38 148 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.217
r382 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r383 34 147 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.76 $Y=1.025
+ $X2=3.76 $Y2=1.217
r384 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.76 $Y=1.025
+ $X2=3.76 $Y2=0.56
r385 31 146 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r386 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r387 27 145 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r388 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r389 24 144 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r390 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r391 20 143 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=1.217
r392 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=0.56
r393 17 141 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r394 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r395 13 140 20.5661 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r396 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
r397 4 115 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.31
r398 4 113 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.63
r399 3 101 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.31
r400 3 99 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.63
r401 2 119 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.56
r402 1 105 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_12%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 36 40 44 48
+ 52 54 58 60 64 66 70 74 76 78 83 88 95 96 102 104 107 110 113 116 119 122 125
+ 128 133
r149 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r150 123 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r151 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r152 120 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r153 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r154 117 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r155 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r156 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r157 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r158 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r159 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r160 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r161 102 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.2 $Y2=2.72
r162 101 133 0.12093 $w=4.8e-07 $l=4.25e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.655 $Y2=2.72
r163 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r164 98 128 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.655 $Y2=2.72
r165 98 100 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r166 96 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r167 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r168 93 125 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.945 $Y=2.72
+ $X2=7.755 $Y2=2.72
r169 93 95 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.945 $Y=2.72
+ $X2=8.05 $Y2=2.72
r170 92 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r171 92 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r172 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r173 89 113 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=3.995 $Y2=2.72
r174 89 91 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.37 $Y2=2.72
r175 88 116 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.745 $Y=2.72
+ $X2=4.935 $Y2=2.72
r176 88 91 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.745 $Y=2.72
+ $X2=4.37 $Y2=2.72
r177 87 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r178 87 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r179 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r180 84 110 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.055 $Y2=2.72
r181 84 86 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.45 $Y2=2.72
r182 83 113 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.995 $Y2=2.72
r183 83 86 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.45 $Y2=2.72
r184 82 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r185 82 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r186 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r187 79 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.14 $Y2=2.72
r188 79 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.53 $Y2=2.72
r189 78 110 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.055 $Y2=2.72
r190 78 81 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.53 $Y2=2.72
r191 76 105 0.126621 $w=4.8e-07 $l=4.45e-07 $layer=MET1_cond $X=0.705 $Y=2.72
+ $X2=1.15 $Y2=2.72
r192 76 133 0.0142271 $w=4.8e-07 $l=5e-08 $layer=MET1_cond $X=0.705 $Y=2.72
+ $X2=0.655 $Y2=2.72
r193 74 102 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.705 $Y=2.72
+ $X2=1.115 $Y2=2.72
r194 74 128 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.705 $Y=2.72
+ $X2=0.655 $Y2=2.72
r195 70 73 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=7.755 $Y=1.66
+ $X2=7.755 $Y2=2.34
r196 68 125 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.755 $Y=2.635
+ $X2=7.755 $Y2=2.72
r197 68 73 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=7.755 $Y=2.635
+ $X2=7.755 $Y2=2.34
r198 67 122 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.005 $Y=2.72
+ $X2=6.815 $Y2=2.72
r199 66 125 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.565 $Y=2.72
+ $X2=7.755 $Y2=2.72
r200 66 67 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.565 $Y=2.72
+ $X2=7.005 $Y2=2.72
r201 62 122 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=2.635
+ $X2=6.815 $Y2=2.72
r202 62 64 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=6.815 $Y=2.635
+ $X2=6.815 $Y2=2
r203 61 119 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.065 $Y=2.72
+ $X2=5.875 $Y2=2.72
r204 60 122 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.625 $Y=2.72
+ $X2=6.815 $Y2=2.72
r205 60 61 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.625 $Y=2.72
+ $X2=6.065 $Y2=2.72
r206 56 119 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=2.635
+ $X2=5.875 $Y2=2.72
r207 56 58 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=5.875 $Y=2.635
+ $X2=5.875 $Y2=2
r208 55 116 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.125 $Y=2.72
+ $X2=4.935 $Y2=2.72
r209 54 119 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.685 $Y=2.72
+ $X2=5.875 $Y2=2.72
r210 54 55 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.685 $Y=2.72
+ $X2=5.125 $Y2=2.72
r211 50 116 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.935 $Y=2.635
+ $X2=4.935 $Y2=2.72
r212 50 52 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=4.935 $Y=2.635
+ $X2=4.935 $Y2=2
r213 46 113 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=2.635
+ $X2=3.995 $Y2=2.72
r214 46 48 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.995 $Y=2.635
+ $X2=3.995 $Y2=2
r215 42 110 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=2.635
+ $X2=3.055 $Y2=2.72
r216 42 44 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.055 $Y=2.635
+ $X2=3.055 $Y2=2
r217 38 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r218 38 40 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r219 37 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.2 $Y2=2.72
r220 36 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.14 $Y2=2.72
r221 36 37 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r222 32 104 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r223 32 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r224 28 100 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.172 $Y2=2.72
r225 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2
r226 9 73 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=2.34
r227 9 70 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=1.66
r228 8 64 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=2
r229 7 58 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=2
r230 6 52 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=2
r231 5 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2
r232 4 44 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r233 3 40 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r234 2 34 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r235 1 30 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_12%X 1 2 3 4 5 6 7 8 9 10 11 12 39 43 45 46 47
+ 48 51 55 57 59 63 67 69 71 75 79 83 87 91 93 94 95 96 97 106 110 112 117
r184 116 117 13.0318 $w=8.78e-07 $l=9.4e-07 $layer=LI1_cond $X=6.37 $Y=1.175
+ $X2=7.31 $Y2=1.175
r185 115 116 13.0318 $w=8.78e-07 $l=9.4e-07 $layer=LI1_cond $X=5.43 $Y=1.175
+ $X2=6.37 $Y2=1.175
r186 110 112 0.138636 $w=8.78e-07 $l=1e-08 $layer=LI1_cond $X=5.325 $Y=1.175
+ $X2=5.335 $Y2=1.175
r187 97 115 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=5.43 $Y=1.615
+ $X2=5.43 $Y2=1.175
r188 97 115 1.17841 $w=8.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=1.175
+ $X2=5.43 $Y2=1.175
r189 97 112 0.138636 $w=8.78e-07 $l=1e-08 $layer=LI1_cond $X=5.345 $Y=1.175
+ $X2=5.335 $Y2=1.175
r190 97 106 7.61063 $w=2.53e-07 $l=1.4e-07 $layer=LI1_cond $X=5.43 $Y=1.615
+ $X2=5.43 $Y2=1.755
r191 89 117 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=7.31 $Y=1.615
+ $X2=7.31 $Y2=1.175
r192 89 91 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=7.31 $Y=1.615
+ $X2=7.31 $Y2=1.755
r193 85 117 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=7.31 $Y=0.735
+ $X2=7.31 $Y2=1.175
r194 85 87 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.31 $Y=0.735
+ $X2=7.31 $Y2=0.56
r195 81 116 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=6.37 $Y=1.615
+ $X2=6.37 $Y2=1.175
r196 81 83 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.37 $Y=1.615
+ $X2=6.37 $Y2=1.755
r197 77 116 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=6.37 $Y=0.735
+ $X2=6.37 $Y2=1.175
r198 77 79 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.37 $Y=0.735
+ $X2=6.37 $Y2=0.56
r199 73 115 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=5.43 $Y=0.735
+ $X2=5.43 $Y2=1.175
r200 73 75 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.43 $Y=0.735
+ $X2=5.43 $Y2=0.56
r201 72 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=1.53
+ $X2=4.49 $Y2=1.53
r202 71 110 4.3386 $w=4.4e-07 $l=4.08473e-07 $layer=LI1_cond $X=5.21 $Y=1.53
+ $X2=5.325 $Y2=1.175
r203 71 72 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.21 $Y=1.53
+ $X2=4.575 $Y2=1.53
r204 70 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=0.82
+ $X2=4.49 $Y2=0.82
r205 69 110 4.3386 $w=4.4e-07 $l=4.08473e-07 $layer=LI1_cond $X=5.21 $Y=0.82
+ $X2=5.325 $Y2=1.175
r206 69 70 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.21 $Y=0.82
+ $X2=4.575 $Y2=0.82
r207 65 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=1.615
+ $X2=4.49 $Y2=1.53
r208 65 67 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.49 $Y=1.615
+ $X2=4.49 $Y2=1.755
r209 61 95 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.735
+ $X2=4.49 $Y2=0.82
r210 61 63 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.49 $Y=0.735
+ $X2=4.49 $Y2=0.56
r211 60 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=1.53
+ $X2=3.55 $Y2=1.53
r212 59 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=1.53
+ $X2=4.49 $Y2=1.53
r213 59 60 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.405 $Y=1.53
+ $X2=3.635 $Y2=1.53
r214 58 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0.82
+ $X2=3.55 $Y2=0.82
r215 57 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=0.82
+ $X2=4.49 $Y2=0.82
r216 57 58 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.405 $Y=0.82
+ $X2=3.635 $Y2=0.82
r217 53 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=1.615
+ $X2=3.55 $Y2=1.53
r218 53 55 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.55 $Y=1.615
+ $X2=3.55 $Y2=1.755
r219 49 93 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.735
+ $X2=3.55 $Y2=0.82
r220 49 51 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.55 $Y=0.735
+ $X2=3.55 $Y2=0.56
r221 47 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=1.53
+ $X2=3.55 $Y2=1.53
r222 47 48 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.465 $Y=1.53
+ $X2=2.695 $Y2=1.53
r223 45 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=0.82
+ $X2=3.55 $Y2=0.82
r224 45 46 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.465 $Y=0.82
+ $X2=2.695 $Y2=0.82
r225 41 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.61 $Y=1.615
+ $X2=2.695 $Y2=1.53
r226 41 43 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.61 $Y=1.615
+ $X2=2.61 $Y2=1.755
r227 37 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.61 $Y=0.735
+ $X2=2.695 $Y2=0.82
r228 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.61 $Y=0.735
+ $X2=2.61 $Y2=0.56
r229 12 91 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=1.755
r230 11 83 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=1.755
r231 10 106 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.755
r232 9 67 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.755
r233 8 55 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.755
r234 7 43 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.755
r235 6 87 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=7.125
+ $Y=0.235 $X2=7.31 $Y2=0.56
r236 5 79 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=6.185
+ $Y=0.235 $X2=6.37 $Y2=0.56
r237 4 75 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=5.245
+ $Y=0.235 $X2=5.43 $Y2=0.56
r238 3 63 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.56
r239 2 51 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.56
r240 1 39 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_12%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 52 56 58 62 64 68 70 72 74 80 85 90 95 102 103 109 112 115 118 121 124 127 130
r162 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r163 128 131 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r164 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r165 125 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r166 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r167 122 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r168 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r169 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r170 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r171 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r172 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r173 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r174 103 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r175 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r176 100 130 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.945 $Y=0
+ $X2=7.755 $Y2=0
r177 100 102 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.945 $Y=0
+ $X2=8.05 $Y2=0
r178 99 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r179 99 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=3.91 $Y2=0
r180 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r181 96 118 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=3.995 $Y2=0
r182 96 98 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=4.37 $Y2=0
r183 95 121 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.745 $Y=0
+ $X2=4.935 $Y2=0
r184 95 98 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.745 $Y=0
+ $X2=4.37 $Y2=0
r185 94 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r186 94 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.99 $Y2=0
r187 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r188 91 115 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.245 $Y=0
+ $X2=3.055 $Y2=0
r189 91 93 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.245 $Y=0
+ $X2=3.45 $Y2=0
r190 90 118 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=0
+ $X2=3.995 $Y2=0
r191 90 93 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.805 $Y=0
+ $X2=3.45 $Y2=0
r192 89 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.99 $Y2=0
r193 89 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.07 $Y2=0
r194 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r195 86 112 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.115 $Y2=0
r196 86 88 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.53 $Y2=0
r197 85 115 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=3.055 $Y2=0
r198 85 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=2.53 $Y2=0
r199 84 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.07 $Y2=0
r200 84 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=1.15 $Y2=0
r201 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r202 81 109 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0
+ $X2=1.175 $Y2=0
r203 81 83 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r204 80 112 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.925 $Y=0
+ $X2=2.115 $Y2=0
r205 80 83 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.925 $Y=0
+ $X2=1.61 $Y2=0
r206 75 106 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r207 74 109 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0
+ $X2=1.175 $Y2=0
r208 72 110 0.142271 $w=4.8e-07 $l=5e-07 $layer=MET1_cond $X=0.65 $Y=0 $X2=1.15
+ $Y2=0
r209 72 107 0.119507 $w=4.8e-07 $l=4.2e-07 $layer=MET1_cond $X=0.65 $Y=0
+ $X2=0.23 $Y2=0
r210 70 74 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.65 $Y=0
+ $X2=0.985 $Y2=0
r211 70 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r212 70 75 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.65 $Y=0
+ $X2=0.425 $Y2=0
r213 66 130 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.755 $Y=0.085
+ $X2=7.755 $Y2=0
r214 66 68 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=7.755 $Y=0.085
+ $X2=7.755 $Y2=0.38
r215 65 127 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=6.815 $Y2=0
r216 64 130 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.565 $Y=0
+ $X2=7.755 $Y2=0
r217 64 65 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.565 $Y=0
+ $X2=7.005 $Y2=0
r218 60 127 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=0.085
+ $X2=6.815 $Y2=0
r219 60 62 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=6.815 $Y=0.085
+ $X2=6.815 $Y2=0.4
r220 59 124 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.065 $Y=0
+ $X2=5.875 $Y2=0
r221 58 127 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.625 $Y=0
+ $X2=6.815 $Y2=0
r222 58 59 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.625 $Y=0
+ $X2=6.065 $Y2=0
r223 54 124 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=0.085
+ $X2=5.875 $Y2=0
r224 54 56 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=5.875 $Y=0.085
+ $X2=5.875 $Y2=0.4
r225 53 121 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.125 $Y=0
+ $X2=4.935 $Y2=0
r226 52 124 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.685 $Y=0
+ $X2=5.875 $Y2=0
r227 52 53 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.685 $Y=0
+ $X2=5.125 $Y2=0
r228 48 121 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.935 $Y=0.085
+ $X2=4.935 $Y2=0
r229 48 50 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=4.935 $Y=0.085
+ $X2=4.935 $Y2=0.4
r230 44 118 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=0.085
+ $X2=3.995 $Y2=0
r231 44 46 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.995 $Y=0.085
+ $X2=3.995 $Y2=0.4
r232 40 115 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0
r233 40 42 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.4
r234 36 112 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=0.085
+ $X2=2.115 $Y2=0
r235 36 38 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.115 $Y=0.085
+ $X2=2.115 $Y2=0.4
r236 32 109 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=0.085
+ $X2=1.175 $Y2=0
r237 32 34 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.175 $Y=0.085
+ $X2=1.175 $Y2=0.4
r238 28 106 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r239 28 30 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r240 9 68 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.645
+ $Y=0.235 $X2=7.78 $Y2=0.38
r241 8 62 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.235 $X2=6.84 $Y2=0.4
r242 7 56 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=5.715
+ $Y=0.235 $X2=5.9 $Y2=0.4
r243 6 50 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.4
r244 5 46 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.4
r245 4 42 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.4
r246 3 38 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.4
r247 2 34 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.4
r248 1 30 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

