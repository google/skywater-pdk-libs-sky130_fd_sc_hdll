* File: sky130_fd_sc_hdll__inv_8.pxi.spice
* Created: Thu Aug 27 19:09:38 2020
* 
x_PM_SKY130_FD_SC_HDLL__INV_8%A N_A_c_66_n N_A_M1000_g N_A_c_75_n N_A_M1001_g
+ N_A_c_67_n N_A_M1003_g N_A_c_76_n N_A_M1002_g N_A_c_68_n N_A_M1005_g
+ N_A_c_77_n N_A_M1004_g N_A_c_69_n N_A_M1007_g N_A_c_78_n N_A_M1006_g
+ N_A_c_70_n N_A_M1009_g N_A_c_79_n N_A_M1008_g N_A_c_71_n N_A_M1012_g
+ N_A_c_80_n N_A_M1010_g N_A_c_72_n N_A_M1014_g N_A_c_81_n N_A_M1011_g
+ N_A_c_82_n N_A_M1013_g N_A_c_73_n N_A_M1015_g A A A A A A N_A_c_118_p
+ N_A_c_74_n PM_SKY130_FD_SC_HDLL__INV_8%A
x_PM_SKY130_FD_SC_HDLL__INV_8%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_M1006_s
+ N_VPWR_M1010_s N_VPWR_M1013_s N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n
+ N_VPWR_c_230_n N_VPWR_c_231_n N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n
+ N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n N_VPWR_c_239_n
+ VPWR N_VPWR_c_240_n N_VPWR_c_226_n PM_SKY130_FD_SC_HDLL__INV_8%VPWR
x_PM_SKY130_FD_SC_HDLL__INV_8%Y N_Y_M1000_d N_Y_M1005_d N_Y_M1009_d N_Y_M1014_d
+ N_Y_M1001_d N_Y_M1004_d N_Y_M1008_d N_Y_M1011_d N_Y_c_298_n N_Y_c_299_n
+ N_Y_c_315_n N_Y_c_310_n N_Y_c_316_n N_Y_c_319_n N_Y_c_300_n N_Y_c_326_n
+ N_Y_c_330_n N_Y_c_334_n N_Y_c_301_n N_Y_c_342_n N_Y_c_346_n N_Y_c_350_n
+ N_Y_c_302_n N_Y_c_358_n N_Y_c_362_n N_Y_c_364_n N_Y_c_303_n N_Y_c_311_n
+ N_Y_c_304_n N_Y_c_375_n N_Y_c_305_n N_Y_c_383_n N_Y_c_306_n N_Y_c_391_n
+ N_Y_c_307_n N_Y_c_398_n Y Y PM_SKY130_FD_SC_HDLL__INV_8%Y
x_PM_SKY130_FD_SC_HDLL__INV_8%VGND N_VGND_M1000_s N_VGND_M1003_s N_VGND_M1007_s
+ N_VGND_M1012_s N_VGND_M1015_s N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n
+ N_VGND_c_486_n N_VGND_c_487_n N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n
+ N_VGND_c_491_n N_VGND_c_492_n N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n
+ VGND N_VGND_c_496_n N_VGND_c_497_n PM_SKY130_FD_SC_HDLL__INV_8%VGND
cc_1 VNB N_A_c_66_n 0.0196767f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.995
cc_2 VNB N_A_c_67_n 0.0167606f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=0.995
cc_3 VNB N_A_c_68_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=0.995
cc_4 VNB N_A_c_69_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.045 $Y2=0.995
cc_5 VNB N_A_c_70_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=0.995
cc_6 VNB N_A_c_71_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.985 $Y2=0.995
cc_7 VNB N_A_c_72_n 0.0172f $X=-0.19 $Y=-0.24 $X2=3.455 $Y2=0.995
cc_8 VNB N_A_c_73_n 0.0201252f $X=-0.19 $Y=-0.24 $X2=3.975 $Y2=0.995
cc_9 VNB N_A_c_74_n 0.154713f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=1.202
cc_10 VNB N_VPWR_c_226_n 0.193827f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=1.202
cc_11 VNB N_Y_c_298_n 0.00180816f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=0.995
cc_12 VNB N_Y_c_299_n 0.0121685f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=0.56
cc_13 VNB N_Y_c_300_n 0.00247508f $X=-0.19 $Y=-0.24 $X2=3.455 $Y2=0.995
cc_14 VNB N_Y_c_301_n 0.00247508f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_15 VNB N_Y_c_302_n 0.00247508f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.202
cc_16 VNB N_Y_c_303_n 0.013528f $X=-0.19 $Y=-0.24 $X2=2.54 $Y2=1.202
cc_17 VNB N_Y_c_304_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=3.715 $Y2=1.16
cc_18 VNB N_Y_c_305_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=3.975 $Y2=1.202
cc_19 VNB N_Y_c_306_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.2
cc_20 VNB N_Y_c_307_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB Y 0.0229772f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.2
cc_22 VNB Y 0.0225993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_483_n 0.0145621f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.41
cc_24 VNB N_VGND_c_484_n 0.0171592f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.985
cc_25 VNB N_VGND_c_485_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.07 $Y2=1.41
cc_26 VNB N_VGND_c_486_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=0.56
cc_27 VNB N_VGND_c_487_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.54 $Y2=1.985
cc_28 VNB N_VGND_c_488_n 0.0138791f $X=-0.19 $Y=-0.24 $X2=2.985 $Y2=0.56
cc_29 VNB N_VGND_c_489_n 0.0187699f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=1.41
cc_30 VNB N_VGND_c_490_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=3.455 $Y2=0.995
cc_31 VNB N_VGND_c_491_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=3.455 $Y2=0.56
cc_32 VNB N_VGND_c_492_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=3.48 $Y2=1.41
cc_33 VNB N_VGND_c_493_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=3.48 $Y2=1.985
cc_34 VNB N_VGND_c_494_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=1.41
cc_35 VNB N_VGND_c_495_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=1.985
cc_36 VNB N_VGND_c_496_n 0.019262f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_497_n 0.239985f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=1.202
cc_38 VPB N_A_c_75_n 0.0191922f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.41
cc_39 VPB N_A_c_76_n 0.0162621f $X=-0.19 $Y=1.305 $X2=1.13 $Y2=1.41
cc_40 VPB N_A_c_77_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.41
cc_41 VPB N_A_c_78_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.07 $Y2=1.41
cc_42 VPB N_A_c_79_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=1.41
cc_43 VPB N_A_c_80_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.41
cc_44 VPB N_A_c_81_n 0.0162621f $X=-0.19 $Y=1.305 $X2=3.48 $Y2=1.41
cc_45 VPB N_A_c_82_n 0.0191964f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=1.41
cc_46 VPB N_A_c_74_n 0.0983967f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=1.202
cc_47 VPB N_VPWR_c_227_n 0.0152107f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.41
cc_48 VPB N_VPWR_c_228_n 0.0300031f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.985
cc_49 VPB N_VPWR_c_229_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.07 $Y2=1.41
cc_50 VPB N_VPWR_c_230_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.515 $Y2=0.56
cc_51 VPB N_VPWR_c_231_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=1.985
cc_52 VPB N_VPWR_c_232_n 0.0143252f $X=-0.19 $Y=1.305 $X2=2.985 $Y2=0.56
cc_53 VPB N_VPWR_c_233_n 0.0322726f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.41
cc_54 VPB N_VPWR_c_234_n 0.0206409f $X=-0.19 $Y=1.305 $X2=3.455 $Y2=0.995
cc_55 VPB N_VPWR_c_235_n 0.00324069f $X=-0.19 $Y=1.305 $X2=3.455 $Y2=0.56
cc_56 VPB N_VPWR_c_236_n 0.0206409f $X=-0.19 $Y=1.305 $X2=3.48 $Y2=1.41
cc_57 VPB N_VPWR_c_237_n 0.00324069f $X=-0.19 $Y=1.305 $X2=3.48 $Y2=1.985
cc_58 VPB N_VPWR_c_238_n 0.0206409f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=1.41
cc_59 VPB N_VPWR_c_239_n 0.00324069f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=1.985
cc_60 VPB N_VPWR_c_240_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_226_n 0.0541679f $X=-0.19 $Y=1.305 $X2=1.105 $Y2=1.202
cc_62 VPB N_Y_c_310_n 0.0156116f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=1.41
cc_63 VPB N_Y_c_311_n 0.0132603f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.202
cc_64 VPB Y 0.0109605f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.2
cc_65 VPB Y 0.0107522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 N_A_c_75_n N_VPWR_c_228_n 0.00674649f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_c_76_n N_VPWR_c_229_n 0.0052072f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A_c_77_n N_VPWR_c_229_n 0.004751f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_c_78_n N_VPWR_c_230_n 0.0052072f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_c_79_n N_VPWR_c_230_n 0.004751f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A_c_80_n N_VPWR_c_231_n 0.0052072f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_c_81_n N_VPWR_c_231_n 0.004751f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A_c_82_n N_VPWR_c_233_n 0.00739881f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_75_n N_VPWR_c_234_n 0.00597712f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_c_76_n N_VPWR_c_234_n 0.00673617f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_c_77_n N_VPWR_c_236_n 0.00597712f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_c_78_n N_VPWR_c_236_n 0.00673617f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_c_79_n N_VPWR_c_238_n 0.00597712f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_c_80_n N_VPWR_c_238_n 0.00673617f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_c_81_n N_VPWR_c_240_n 0.00597712f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_c_82_n N_VPWR_c_240_n 0.00673617f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_c_75_n N_VPWR_c_226_n 0.0110272f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_c_76_n N_VPWR_c_226_n 0.0118438f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_77_n N_VPWR_c_226_n 0.00999457f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_c_78_n N_VPWR_c_226_n 0.0118438f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_c_79_n N_VPWR_c_226_n 0.00999457f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_c_80_n N_VPWR_c_226_n 0.0118438f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_c_81_n N_VPWR_c_226_n 0.00999457f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_c_82_n N_VPWR_c_226_n 0.0128707f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_c_66_n N_Y_c_298_n 0.0124108f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_c_75_n N_Y_c_315_n 0.0131889f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_c_66_n N_Y_c_316_n 0.0109371f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_c_67_n N_Y_c_316_n 0.00674948f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_c_68_n N_Y_c_316_n 5.42233e-19 $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_c_75_n N_Y_c_319_n 0.0178402f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_c_76_n N_Y_c_319_n 0.0106251f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_c_77_n N_Y_c_319_n 6.24674e-19 $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_c_67_n N_Y_c_300_n 0.00923615f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_c_68_n N_Y_c_300_n 0.00923615f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_c_118_p N_Y_c_300_n 0.0405926f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_c_74_n N_Y_c_300_n 0.00346f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_102 N_A_c_76_n N_Y_c_326_n 0.0137916f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_77_n N_Y_c_326_n 0.0101048f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_c_118_p N_Y_c_326_n 0.0356113f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_c_74_n N_Y_c_326_n 0.00635951f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_106 N_A_c_67_n N_Y_c_330_n 5.22028e-19 $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_c_68_n N_Y_c_330_n 0.00641183f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_c_69_n N_Y_c_330_n 0.00674948f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_c_70_n N_Y_c_330_n 5.42233e-19 $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_c_76_n N_Y_c_334_n 6.48386e-19 $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_77_n N_Y_c_334_n 0.0130707f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_c_78_n N_Y_c_334_n 0.0106251f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_c_79_n N_Y_c_334_n 6.24674e-19 $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_c_69_n N_Y_c_301_n 0.00923615f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_c_70_n N_Y_c_301_n 0.00923615f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_c_118_p N_Y_c_301_n 0.0405926f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_c_74_n N_Y_c_301_n 0.00346f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_118 N_A_c_78_n N_Y_c_342_n 0.0137916f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_79_n N_Y_c_342_n 0.0101048f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_118_p N_Y_c_342_n 0.0356113f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_c_74_n N_Y_c_342_n 0.00635951f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_122 N_A_c_69_n N_Y_c_346_n 5.22028e-19 $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_c_70_n N_Y_c_346_n 0.00641183f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_c_71_n N_Y_c_346_n 0.00674948f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_72_n N_Y_c_346_n 5.42233e-19 $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_78_n N_Y_c_350_n 6.48386e-19 $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_c_79_n N_Y_c_350_n 0.0130707f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_c_80_n N_Y_c_350_n 0.0106251f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_81_n N_Y_c_350_n 6.24674e-19 $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_71_n N_Y_c_302_n 0.00923615f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_72_n N_Y_c_302_n 0.00923615f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_118_p N_Y_c_302_n 0.0405926f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_c_74_n N_Y_c_302_n 0.00346f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_134 N_A_c_80_n N_Y_c_358_n 0.0137916f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_81_n N_Y_c_358_n 0.0101048f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_c_118_p N_Y_c_358_n 0.0356113f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_74_n N_Y_c_358_n 0.00635951f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_138 N_A_c_71_n N_Y_c_362_n 5.22028e-19 $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_c_72_n N_Y_c_362_n 0.00641183f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_c_80_n N_Y_c_364_n 6.48386e-19 $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_81_n N_Y_c_364_n 0.0130707f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_82_n N_Y_c_364_n 0.0153658f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_73_n N_Y_c_303_n 0.014747f $X=3.975 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_c_118_p N_Y_c_303_n 3.32968e-19 $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_c_82_n N_Y_c_311_n 0.0173759f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_118_p N_Y_c_311_n 3.15358e-19 $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_c_66_n N_Y_c_304_n 0.00119366f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_c_67_n N_Y_c_304_n 0.00119366f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_c_118_p N_Y_c_304_n 0.031064f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_c_74_n N_Y_c_304_n 0.00358305f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_151 N_A_c_75_n N_Y_c_375_n 0.00210477f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_76_n N_Y_c_375_n 5.79575e-19 $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_118_p N_Y_c_375_n 0.0253353f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_c_74_n N_Y_c_375_n 0.00651614f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_155 N_A_c_68_n N_Y_c_305_n 0.00119366f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_c_69_n N_Y_c_305_n 0.00119366f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_c_118_p N_Y_c_305_n 0.031064f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_c_74_n N_Y_c_305_n 0.00358305f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_159 N_A_c_77_n N_Y_c_383_n 0.00210477f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_78_n N_Y_c_383_n 5.79575e-19 $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_118_p N_Y_c_383_n 0.0253353f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_c_74_n N_Y_c_383_n 0.00651614f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_163 N_A_c_70_n N_Y_c_306_n 0.00119366f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_71_n N_Y_c_306_n 0.00119366f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_118_p N_Y_c_306_n 0.031064f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_c_74_n N_Y_c_306_n 0.00358305f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_167 N_A_c_79_n N_Y_c_391_n 0.00210477f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_c_80_n N_Y_c_391_n 5.79575e-19 $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_118_p N_Y_c_391_n 0.0253353f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_c_74_n N_Y_c_391_n 0.00651614f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_171 N_A_c_72_n N_Y_c_307_n 0.00122295f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_118_p N_Y_c_307_n 0.0311977f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_c_74_n N_Y_c_307_n 0.00486271f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_174 N_A_c_81_n N_Y_c_398_n 0.00210477f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_82_n N_Y_c_398_n 5.79575e-19 $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_118_p N_Y_c_398_n 0.0253353f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_c_74_n N_Y_c_398_n 0.00631893f $X=3.95 $Y=1.202 $X2=0 $Y2=0
cc_178 N_A_c_66_n Y 0.0179374f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_75_n Y 0.0032992f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_c_118_p Y 0.015622f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_c_82_n Y 0.0032512f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_c_73_n Y 0.0178942f $X=3.975 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_c_118_p Y 0.0135527f $X=3.715 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_c_66_n N_VGND_c_484_n 0.00450113f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_c_67_n N_VGND_c_485_n 0.00376026f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_c_68_n N_VGND_c_485_n 0.00276126f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_69_n N_VGND_c_486_n 0.00376026f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_70_n N_VGND_c_486_n 0.00276126f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_71_n N_VGND_c_487_n 0.00376026f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_72_n N_VGND_c_487_n 0.00276126f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_73_n N_VGND_c_489_n 0.00455358f $X=3.975 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_c_66_n N_VGND_c_490_n 0.00422241f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_67_n N_VGND_c_490_n 0.00422241f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_68_n N_VGND_c_492_n 0.00422241f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_69_n N_VGND_c_492_n 0.00422241f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_70_n N_VGND_c_494_n 0.00422241f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_71_n N_VGND_c_494_n 0.00422241f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_c_72_n N_VGND_c_496_n 0.00422241f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_c_73_n N_VGND_c_496_n 0.00436487f $X=3.975 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_c_66_n N_VGND_c_497_n 0.0069027f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_67_n N_VGND_c_497_n 0.00607326f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_c_68_n N_VGND_c_497_n 0.0059505f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_c_69_n N_VGND_c_497_n 0.00607326f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_c_70_n N_VGND_c_497_n 0.0059505f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_c_71_n N_VGND_c_497_n 0.00607326f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_c_72_n N_VGND_c_497_n 0.00606584f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_c_73_n N_VGND_c_497_n 0.00717772f $X=3.975 $Y=0.995 $X2=0 $Y2=0
cc_208 N_VPWR_c_226_n N_Y_M1001_d 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_209 N_VPWR_c_226_n N_Y_M1004_d 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_210 N_VPWR_c_226_n N_Y_M1008_d 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_211 N_VPWR_c_226_n N_Y_M1011_d 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_212 N_VPWR_M1001_s N_Y_c_315_n 0.00234708f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_213 N_VPWR_c_228_n N_Y_c_315_n 0.00639085f $X=0.425 $Y=2 $X2=0 $Y2=0
cc_214 N_VPWR_M1001_s N_Y_c_310_n 0.0022744f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_215 N_VPWR_c_228_n N_Y_c_310_n 0.0157986f $X=0.425 $Y=2 $X2=0 $Y2=0
cc_216 N_VPWR_c_228_n N_Y_c_319_n 0.048465f $X=0.425 $Y=2 $X2=0 $Y2=0
cc_217 N_VPWR_c_229_n N_Y_c_319_n 0.0385613f $X=1.365 $Y=2 $X2=0 $Y2=0
cc_218 N_VPWR_c_234_n N_Y_c_319_n 0.0223557f $X=1.28 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_c_226_n N_Y_c_319_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_M1002_s N_Y_c_326_n 0.00325884f $X=1.22 $Y=1.485 $X2=0 $Y2=0
cc_221 N_VPWR_c_229_n N_Y_c_326_n 0.0136682f $X=1.365 $Y=2 $X2=0 $Y2=0
cc_222 N_VPWR_c_229_n N_Y_c_334_n 0.0470327f $X=1.365 $Y=2 $X2=0 $Y2=0
cc_223 N_VPWR_c_230_n N_Y_c_334_n 0.0385613f $X=2.305 $Y=2 $X2=0 $Y2=0
cc_224 N_VPWR_c_236_n N_Y_c_334_n 0.0223557f $X=2.22 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_c_226_n N_Y_c_334_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_226 N_VPWR_M1006_s N_Y_c_342_n 0.00325884f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_227 N_VPWR_c_230_n N_Y_c_342_n 0.0136682f $X=2.305 $Y=2 $X2=0 $Y2=0
cc_228 N_VPWR_c_230_n N_Y_c_350_n 0.0470327f $X=2.305 $Y=2 $X2=0 $Y2=0
cc_229 N_VPWR_c_231_n N_Y_c_350_n 0.0385613f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_230 N_VPWR_c_238_n N_Y_c_350_n 0.0223557f $X=3.16 $Y=2.72 $X2=0 $Y2=0
cc_231 N_VPWR_c_226_n N_Y_c_350_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_M1010_s N_Y_c_358_n 0.00325884f $X=3.1 $Y=1.485 $X2=0 $Y2=0
cc_233 N_VPWR_c_231_n N_Y_c_358_n 0.0136682f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_234 N_VPWR_c_231_n N_Y_c_364_n 0.0470327f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_235 N_VPWR_c_233_n N_Y_c_364_n 0.0402386f $X=4.185 $Y=2 $X2=0 $Y2=0
cc_236 N_VPWR_c_240_n N_Y_c_364_n 0.0223557f $X=4.1 $Y=2.72 $X2=0 $Y2=0
cc_237 N_VPWR_c_226_n N_Y_c_364_n 0.0140101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_238 N_VPWR_M1013_s N_Y_c_311_n 0.00471186f $X=4.04 $Y=1.485 $X2=0 $Y2=0
cc_239 N_VPWR_c_233_n N_Y_c_311_n 0.0263619f $X=4.185 $Y=2 $X2=0 $Y2=0
cc_240 N_Y_c_298_n N_VGND_M1000_s 7.48374e-19 $X=0.68 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_241 N_Y_c_299_n N_VGND_M1000_s 0.00215453f $X=0.43 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_242 N_Y_c_300_n N_VGND_M1003_s 0.0025045f $X=1.62 $Y=0.81 $X2=0 $Y2=0
cc_243 N_Y_c_301_n N_VGND_M1007_s 0.0025045f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_244 N_Y_c_302_n N_VGND_M1012_s 0.0025045f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_245 N_Y_c_303_n N_VGND_M1015_s 0.00290096f $X=4.185 $Y=0.81 $X2=0 $Y2=0
cc_246 N_Y_c_299_n N_VGND_c_483_n 0.00295616f $X=0.43 $Y=0.81 $X2=0 $Y2=0
cc_247 N_Y_c_298_n N_VGND_c_484_n 0.00570628f $X=0.68 $Y=0.81 $X2=0 $Y2=0
cc_248 N_Y_c_299_n N_VGND_c_484_n 0.0151569f $X=0.43 $Y=0.81 $X2=0 $Y2=0
cc_249 N_Y_c_316_n N_VGND_c_485_n 0.0177507f $X=0.895 $Y=0.38 $X2=0 $Y2=0
cc_250 N_Y_c_300_n N_VGND_c_485_n 0.0127393f $X=1.62 $Y=0.81 $X2=0 $Y2=0
cc_251 N_Y_c_330_n N_VGND_c_486_n 0.0177507f $X=1.835 $Y=0.38 $X2=0 $Y2=0
cc_252 N_Y_c_301_n N_VGND_c_486_n 0.0127393f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_253 N_Y_c_346_n N_VGND_c_487_n 0.0177507f $X=2.775 $Y=0.38 $X2=0 $Y2=0
cc_254 N_Y_c_302_n N_VGND_c_487_n 0.0127393f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_255 N_Y_c_303_n N_VGND_c_488_n 0.00173892f $X=4.185 $Y=0.81 $X2=0 $Y2=0
cc_256 N_Y_c_303_n N_VGND_c_489_n 0.0253066f $X=4.185 $Y=0.81 $X2=0 $Y2=0
cc_257 N_Y_c_298_n N_VGND_c_490_n 0.00203746f $X=0.68 $Y=0.81 $X2=0 $Y2=0
cc_258 N_Y_c_316_n N_VGND_c_490_n 0.0223596f $X=0.895 $Y=0.38 $X2=0 $Y2=0
cc_259 N_Y_c_300_n N_VGND_c_490_n 0.00273345f $X=1.62 $Y=0.81 $X2=0 $Y2=0
cc_260 N_Y_c_300_n N_VGND_c_492_n 0.00203746f $X=1.62 $Y=0.81 $X2=0 $Y2=0
cc_261 N_Y_c_330_n N_VGND_c_492_n 0.0223596f $X=1.835 $Y=0.38 $X2=0 $Y2=0
cc_262 N_Y_c_301_n N_VGND_c_492_n 0.00273345f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_263 N_Y_c_301_n N_VGND_c_494_n 0.00203746f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_264 N_Y_c_346_n N_VGND_c_494_n 0.0223596f $X=2.775 $Y=0.38 $X2=0 $Y2=0
cc_265 N_Y_c_302_n N_VGND_c_494_n 0.00273345f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_266 N_Y_c_302_n N_VGND_c_496_n 0.00203746f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_267 N_Y_c_362_n N_VGND_c_496_n 0.0231806f $X=3.715 $Y=0.38 $X2=0 $Y2=0
cc_268 N_Y_c_303_n N_VGND_c_496_n 0.00260993f $X=4.185 $Y=0.81 $X2=0 $Y2=0
cc_269 N_Y_M1000_d N_VGND_c_497_n 0.0025535f $X=0.71 $Y=0.235 $X2=0 $Y2=0
cc_270 N_Y_M1005_d N_VGND_c_497_n 0.0025535f $X=1.65 $Y=0.235 $X2=0 $Y2=0
cc_271 N_Y_M1009_d N_VGND_c_497_n 0.0025535f $X=2.59 $Y=0.235 $X2=0 $Y2=0
cc_272 N_Y_M1014_d N_VGND_c_497_n 0.0030386f $X=3.53 $Y=0.235 $X2=0 $Y2=0
cc_273 N_Y_c_298_n N_VGND_c_497_n 0.00420836f $X=0.68 $Y=0.81 $X2=0 $Y2=0
cc_274 N_Y_c_299_n N_VGND_c_497_n 0.00562823f $X=0.43 $Y=0.81 $X2=0 $Y2=0
cc_275 N_Y_c_316_n N_VGND_c_497_n 0.0141302f $X=0.895 $Y=0.38 $X2=0 $Y2=0
cc_276 N_Y_c_300_n N_VGND_c_497_n 0.00983903f $X=1.62 $Y=0.81 $X2=0 $Y2=0
cc_277 N_Y_c_330_n N_VGND_c_497_n 0.0141302f $X=1.835 $Y=0.38 $X2=0 $Y2=0
cc_278 N_Y_c_301_n N_VGND_c_497_n 0.00983903f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_279 N_Y_c_346_n N_VGND_c_497_n 0.0141302f $X=2.775 $Y=0.38 $X2=0 $Y2=0
cc_280 N_Y_c_302_n N_VGND_c_497_n 0.00983903f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_281 N_Y_c_362_n N_VGND_c_497_n 0.0143352f $X=3.715 $Y=0.38 $X2=0 $Y2=0
cc_282 N_Y_c_303_n N_VGND_c_497_n 0.00920694f $X=4.185 $Y=0.81 $X2=0 $Y2=0
