* File: sky130_fd_sc_hdll__nor4_4.pex.spice
* Created: Thu Aug 27 19:17:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 38 39 44
r72 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r73 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=1.75 $Y=1.202
+ $X2=1.925 $Y2=1.202
r74 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.75
+ $Y=1.16 $X2=1.75 $Y2=1.16
r75 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.75 $Y2=1.202
r76 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r77 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.43 $Y2=1.202
r78 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r79 31 44 30.368 $w=2.08e-07 $l=5.75e-07 $layer=LI1_cond $X=0.58 $Y=1.18
+ $X2=1.155 $Y2=1.18
r80 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=0.58 $Y=1.202
+ $X2=0.96 $Y2=1.202
r81 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.16 $X2=0.58 $Y2=1.16
r82 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.58 $Y2=1.202
r83 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r84 25 38 26.1429 $w=2.08e-07 $l=4.95e-07 $layer=LI1_cond $X=1.255 $Y=1.18
+ $X2=1.75 $Y2=1.18
r85 25 44 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=1.255 $Y=1.18
+ $X2=1.155 $Y2=1.18
r86 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r87 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r88 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r89 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r90 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r91 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r92 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r93 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r94 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r95 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r96 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r97 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=0.56
r98 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r99 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r100 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r101 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 27 43 48 54
r76 43 44 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.805 $Y=1.202
+ $X2=3.83 $Y2=1.202
r77 41 43 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=3.63 $Y=1.202
+ $X2=3.805 $Y2=1.202
r78 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.63
+ $Y=1.16 $X2=3.63 $Y2=1.16
r79 39 41 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=3.335 $Y=1.202
+ $X2=3.63 $Y2=1.202
r80 38 39 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.31 $Y=1.202
+ $X2=3.335 $Y2=1.202
r81 37 38 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.865 $Y=1.202
+ $X2=3.31 $Y2=1.202
r82 36 37 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.84 $Y=1.202
+ $X2=2.865 $Y2=1.202
r83 35 48 42.7792 $w=2.08e-07 $l=8.1e-07 $layer=LI1_cond $X=2.46 $Y=1.18
+ $X2=3.27 $Y2=1.18
r84 34 36 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=2.46 $Y=1.202
+ $X2=2.84 $Y2=1.202
r85 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r86 32 34 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.46 $Y2=1.202
r87 31 32 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.37 $Y=1.202
+ $X2=2.395 $Y2=1.202
r88 27 54 1.05628 $w=2.08e-07 $l=2e-08 $layer=LI1_cond $X=4.315 $Y=1.18
+ $X2=4.295 $Y2=1.18
r89 26 54 25.8788 $w=2.08e-07 $l=4.9e-07 $layer=LI1_cond $X=3.805 $Y=1.18
+ $X2=4.295 $Y2=1.18
r90 26 42 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=3.805 $Y=1.18
+ $X2=3.63 $Y2=1.18
r91 25 42 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=3.295 $Y=1.18
+ $X2=3.63 $Y2=1.18
r92 25 48 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=3.295 $Y=1.18
+ $X2=3.27 $Y2=1.18
r93 22 44 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=1.202
r94 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=0.56
r95 19 43 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.202
r96 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.985
r97 16 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.202
r98 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.985
r99 13 38 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=1.202
r100 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=0.56
r101 10 37 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.202
r102 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.985
r103 7 36 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=1.202
r104 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=0.56
r105 4 32 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.202
r106 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r107 1 31 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=1.202
r108 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%C 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 38 39 44
r76 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.205 $Y=1.202
+ $X2=6.23 $Y2=1.202
r77 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=6.03 $Y=1.202
+ $X2=6.205 $Y2=1.202
r78 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.03
+ $Y=1.16 $X2=6.03 $Y2=1.16
r79 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=5.735 $Y=1.202
+ $X2=6.03 $Y2=1.202
r80 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.71 $Y=1.202
+ $X2=5.735 $Y2=1.202
r81 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=5.265 $Y=1.202
+ $X2=5.71 $Y2=1.202
r82 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.24 $Y=1.202
+ $X2=5.265 $Y2=1.202
r83 31 44 22.1818 $w=2.08e-07 $l=4.2e-07 $layer=LI1_cond $X=4.86 $Y=1.18
+ $X2=5.28 $Y2=1.18
r84 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=4.86 $Y=1.202
+ $X2=5.24 $Y2=1.202
r85 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.86
+ $Y=1.16 $X2=4.86 $Y2=1.16
r86 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=4.795 $Y=1.202
+ $X2=4.86 $Y2=1.202
r87 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.77 $Y=1.202
+ $X2=4.795 $Y2=1.202
r88 25 38 39.3463 $w=2.08e-07 $l=7.45e-07 $layer=LI1_cond $X=5.285 $Y=1.18
+ $X2=6.03 $Y2=1.18
r89 25 44 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=5.285 $Y=1.18
+ $X2=5.28 $Y2=1.18
r90 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.23 $Y=0.995
+ $X2=6.23 $Y2=1.202
r91 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.23 $Y=0.995
+ $X2=6.23 $Y2=0.56
r92 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.205 $Y=1.41
+ $X2=6.205 $Y2=1.202
r93 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.205 $Y=1.41
+ $X2=6.205 $Y2=1.985
r94 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.735 $Y=1.41
+ $X2=5.735 $Y2=1.202
r95 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.735 $Y=1.41
+ $X2=5.735 $Y2=1.985
r96 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.71 $Y=0.995
+ $X2=5.71 $Y2=1.202
r97 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.71 $Y=0.995
+ $X2=5.71 $Y2=0.56
r98 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.202
r99 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.985
r100 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=1.202
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=0.56
r102 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.202
r103 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.985
r104 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.202
r105 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%D 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 38 39 44
r77 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.085 $Y=1.202
+ $X2=8.11 $Y2=1.202
r78 37 39 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=7.88 $Y=1.202
+ $X2=8.085 $Y2=1.202
r79 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.88
+ $Y=1.16 $X2=7.88 $Y2=1.16
r80 35 37 34.336 $w=3.72e-07 $l=2.65e-07 $layer=POLY_cond $X=7.615 $Y=1.202
+ $X2=7.88 $Y2=1.202
r81 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.59 $Y=1.202
+ $X2=7.615 $Y2=1.202
r82 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=7.145 $Y=1.202
+ $X2=7.59 $Y2=1.202
r83 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.12 $Y=1.202
+ $X2=7.145 $Y2=1.202
r84 31 44 33.5368 $w=2.08e-07 $l=6.35e-07 $layer=LI1_cond $X=6.71 $Y=1.18
+ $X2=7.345 $Y2=1.18
r85 30 32 53.1237 $w=3.72e-07 $l=4.1e-07 $layer=POLY_cond $X=6.71 $Y=1.202
+ $X2=7.12 $Y2=1.202
r86 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.71
+ $Y=1.16 $X2=6.71 $Y2=1.16
r87 28 30 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=6.675 $Y=1.202
+ $X2=6.71 $Y2=1.202
r88 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.65 $Y=1.202
+ $X2=6.675 $Y2=1.202
r89 25 38 26.671 $w=2.08e-07 $l=5.05e-07 $layer=LI1_cond $X=7.375 $Y=1.18
+ $X2=7.88 $Y2=1.18
r90 25 44 1.58442 $w=2.08e-07 $l=3e-08 $layer=LI1_cond $X=7.375 $Y=1.18
+ $X2=7.345 $Y2=1.18
r91 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.11 $Y=0.995
+ $X2=8.11 $Y2=1.202
r92 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.11 $Y=0.995
+ $X2=8.11 $Y2=0.56
r93 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.085 $Y=1.41
+ $X2=8.085 $Y2=1.202
r94 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.085 $Y=1.41
+ $X2=8.085 $Y2=1.985
r95 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.615 $Y=1.41
+ $X2=7.615 $Y2=1.202
r96 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.615 $Y=1.41
+ $X2=7.615 $Y2=1.985
r97 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.59 $Y=0.995
+ $X2=7.59 $Y2=1.202
r98 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.59 $Y=0.995
+ $X2=7.59 $Y2=0.56
r99 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.145 $Y=1.41
+ $X2=7.145 $Y2=1.202
r100 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.145 $Y=1.41
+ $X2=7.145 $Y2=1.985
r101 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.12 $Y=0.995
+ $X2=7.12 $Y2=1.202
r102 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.12 $Y=0.995
+ $X2=7.12 $Y2=0.56
r103 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.675 $Y=1.41
+ $X2=6.675 $Y2=1.202
r104 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.675 $Y=1.41
+ $X2=6.675 $Y2=1.985
r105 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.65 $Y=0.995
+ $X2=6.65 $Y2=1.202
r106 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.65 $Y=0.995
+ $X2=6.65 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 34 36 40 45 50
r62 38 40 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=4.067 $Y=2.295
+ $X2=4.067 $Y2=1.96
r63 37 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.225 $Y=2.38
+ $X2=3.1 $Y2=2.38
r64 36 38 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=3.915 $Y=2.38
+ $X2=4.067 $Y2=2.295
r65 36 37 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.915 $Y=2.38
+ $X2=3.225 $Y2=2.38
r66 32 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=2.295
+ $X2=3.1 $Y2=2.38
r67 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.1 $Y=2.295
+ $X2=3.1 $Y2=1.96
r68 31 49 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=2.38
+ $X2=2.16 $Y2=2.38
r69 30 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.975 $Y=2.38
+ $X2=3.1 $Y2=2.38
r70 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.975 $Y=2.38
+ $X2=2.285 $Y2=2.38
r71 29 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=2.295
+ $X2=2.16 $Y2=2.38
r72 28 47 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=1.625
+ $X2=2.16 $Y2=1.54
r73 28 29 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.16 $Y=1.625
+ $X2=2.16 $Y2=2.295
r74 27 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=1.54
+ $X2=1.22 $Y2=1.54
r75 26 47 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=2.16 $Y2=1.54
r76 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=1.345 $Y2=1.54
r77 22 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=1.54
r78 22 24 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=2.3
r79 21 43 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.247 $Y2=1.54
r80 20 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=1.22 $Y2=1.54
r81 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=0.405 $Y2=1.54
r82 16 43 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=1.625
+ $X2=0.247 $Y2=1.54
r83 16 18 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=0.247 $Y=1.625
+ $X2=0.247 $Y2=2.3
r84 5 40 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.895
+ $Y=1.485 $X2=4.04 $Y2=1.96
r85 4 34 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=1.96
r86 3 49 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.3
r87 3 47 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.62
r88 2 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r89 2 24 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r90 1 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r91 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%VPWR 1 2 11 13 17 19 26 27 30 33
r92 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r93 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r94 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 26 27 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r96 24 27 1.83245 $w=4.8e-07 $l=6.44e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=8.51 $Y2=2.72
r97 24 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r98 23 26 420.15 $w=1.68e-07 $l=6.44e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=8.51 $Y2=2.72
r99 23 24 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r100 21 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.69 $Y2=2.72
r101 21 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=2.07 $Y2=2.72
r102 19 31 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r103 15 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=2.72
r104 15 17 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=1.96
r105 14 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r106 13 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=1.69 $Y2=2.72
r107 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=0.875 $Y2=2.72
r108 9 30 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r109 9 11 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r110 2 17 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.96
r111 1 11 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%A_497_297# 1 2 3 4 15 19 23 28 30 32 34
r59 24 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=1.54
+ $X2=5.03 $Y2=1.54
r60 23 34 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.845 $Y=1.54
+ $X2=5.97 $Y2=1.54
r61 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.845 $Y=1.54
+ $X2=5.155 $Y2=1.54
r62 20 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.695 $Y=1.54
+ $X2=3.57 $Y2=1.54
r63 19 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=5.03 $Y2=1.54
r64 19 20 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=3.695 $Y2=1.54
r65 16 28 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=1.54
+ $X2=2.63 $Y2=1.54
r66 15 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.445 $Y=1.54
+ $X2=3.57 $Y2=1.54
r67 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.445 $Y=1.54
+ $X2=2.755 $Y2=1.54
r68 4 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.825
+ $Y=1.485 $X2=5.97 $Y2=1.62
r69 3 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.885
+ $Y=1.485 $X2=5.03 $Y2=1.62
r70 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=1.62
r71 1 28 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%A_887_297# 1 2 3 4 5 18 20 21 24 26 30 32
+ 36 38 42 44 45 46
r57 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.32 $Y=2.295
+ $X2=8.32 $Y2=1.96
r58 39 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.505 $Y=2.38
+ $X2=7.38 $Y2=2.38
r59 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.195 $Y=2.38
+ $X2=8.32 $Y2=2.295
r60 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.195 $Y=2.38
+ $X2=7.505 $Y2=2.38
r61 34 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.38 $Y=2.295
+ $X2=7.38 $Y2=2.38
r62 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.38 $Y=2.295
+ $X2=7.38 $Y2=1.96
r63 33 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.565 $Y=2.38
+ $X2=6.44 $Y2=2.38
r64 32 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.255 $Y=2.38
+ $X2=7.38 $Y2=2.38
r65 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.255 $Y=2.38
+ $X2=6.565 $Y2=2.38
r66 28 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=2.295
+ $X2=6.44 $Y2=2.38
r67 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.44 $Y=2.295
+ $X2=6.44 $Y2=1.96
r68 27 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.625 $Y=2.38
+ $X2=5.5 $Y2=2.38
r69 26 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.315 $Y=2.38
+ $X2=6.44 $Y2=2.38
r70 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.315 $Y=2.38
+ $X2=5.625 $Y2=2.38
r71 22 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=2.295
+ $X2=5.5 $Y2=2.38
r72 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.5 $Y=2.295
+ $X2=5.5 $Y2=1.96
r73 20 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.375 $Y=2.38
+ $X2=5.5 $Y2=2.38
r74 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.375 $Y=2.38
+ $X2=4.685 $Y2=2.38
r75 16 21 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.545 $Y=2.295
+ $X2=4.685 $Y2=2.38
r76 16 18 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.545 $Y=2.295
+ $X2=4.545 $Y2=1.96
r77 5 42 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.175
+ $Y=1.485 $X2=8.32 $Y2=1.96
r78 4 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.235
+ $Y=1.485 $X2=7.38 $Y2=1.96
r79 3 30 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.295
+ $Y=1.485 $X2=6.44 $Y2=1.96
r80 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.355
+ $Y=1.485 $X2=5.5 $Y2=1.96
r81 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=4.435
+ $Y=1.485 $X2=4.56 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 39 41 45 47
+ 51 53 57 59 63 65 69 73 75 79 83 85 87 88 89 90 91 92 94 95 97 99 102
r206 99 102 2.87089 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=8.495 $Y=0.815
+ $X2=8.495 $Y2=0.905
r207 99 102 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=8.495 $Y=0.92
+ $X2=8.495 $Y2=0.905
r208 98 99 22.8354 $w=2.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.495 $Y=1.455
+ $X2=8.495 $Y2=0.92
r209 86 95 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.015 $Y=0.815
+ $X2=7.825 $Y2=0.815
r210 85 99 4.30634 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=8.36 $Y=0.815
+ $X2=8.495 $Y2=0.815
r211 85 86 21.2576 $w=1.78e-07 $l=3.45e-07 $layer=LI1_cond $X=8.36 $Y=0.815
+ $X2=8.015 $Y2=0.815
r212 84 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.975 $Y=1.54
+ $X2=7.85 $Y2=1.54
r213 83 98 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=8.36 $Y=1.54
+ $X2=8.495 $Y2=1.455
r214 83 84 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.36 $Y=1.54
+ $X2=7.975 $Y2=1.54
r215 77 95 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.825 $Y=0.725
+ $X2=7.825 $Y2=0.815
r216 77 79 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.825 $Y=0.725
+ $X2=7.825 $Y2=0.39
r217 76 92 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.075 $Y=0.815
+ $X2=6.885 $Y2=0.815
r218 75 95 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.635 $Y=0.815
+ $X2=7.825 $Y2=0.815
r219 75 76 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=7.635 $Y=0.815
+ $X2=7.075 $Y2=0.815
r220 74 94 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.035 $Y=1.54
+ $X2=6.91 $Y2=1.54
r221 73 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.725 $Y=1.54
+ $X2=7.85 $Y2=1.54
r222 73 74 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.725 $Y=1.54
+ $X2=7.035 $Y2=1.54
r223 67 92 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.885 $Y=0.725
+ $X2=6.885 $Y2=0.815
r224 67 69 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.885 $Y=0.725
+ $X2=6.885 $Y2=0.39
r225 66 91 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.135 $Y=0.815
+ $X2=5.945 $Y2=0.815
r226 65 92 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.695 $Y=0.815
+ $X2=6.885 $Y2=0.815
r227 65 66 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.695 $Y=0.815
+ $X2=6.135 $Y2=0.815
r228 61 91 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.945 $Y=0.725
+ $X2=5.945 $Y2=0.815
r229 61 63 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.945 $Y=0.725
+ $X2=5.945 $Y2=0.39
r230 60 90 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.195 $Y=0.815
+ $X2=5.005 $Y2=0.815
r231 59 91 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.755 $Y=0.815
+ $X2=5.945 $Y2=0.815
r232 59 60 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.755 $Y=0.815
+ $X2=5.195 $Y2=0.815
r233 55 90 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.005 $Y=0.725
+ $X2=5.005 $Y2=0.815
r234 55 57 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.005 $Y=0.725
+ $X2=5.005 $Y2=0.39
r235 54 89 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.735 $Y=0.815
+ $X2=3.545 $Y2=0.815
r236 53 90 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.815 $Y=0.815
+ $X2=5.005 $Y2=0.815
r237 53 54 66.5455 $w=1.78e-07 $l=1.08e-06 $layer=LI1_cond $X=4.815 $Y=0.815
+ $X2=3.735 $Y2=0.815
r238 49 89 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.545 $Y2=0.815
r239 49 51 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.545 $Y2=0.39
r240 48 88 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.795 $Y=0.815
+ $X2=2.605 $Y2=0.815
r241 47 89 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=3.545 $Y2=0.815
r242 47 48 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=2.795 $Y2=0.815
r243 43 88 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.605 $Y2=0.815
r244 43 45 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.605 $Y2=0.39
r245 42 87 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=0.815
+ $X2=1.665 $Y2=0.815
r246 41 88 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=2.605 $Y2=0.815
r247 41 42 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=1.855 $Y2=0.815
r248 37 87 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.815
r249 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.39
r250 35 87 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=1.665 $Y2=0.815
r251 35 36 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=0.915 $Y2=0.815
r252 31 36 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.815
r253 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r254 10 97 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=7.705
+ $Y=1.485 $X2=7.85 $Y2=1.62
r255 9 94 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.765
+ $Y=1.485 $X2=6.91 $Y2=1.62
r256 8 79 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.665
+ $Y=0.235 $X2=7.85 $Y2=0.39
r257 7 69 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.725
+ $Y=0.235 $X2=6.91 $Y2=0.39
r258 6 63 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.785
+ $Y=0.235 $X2=5.97 $Y2=0.39
r259 5 57 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.845
+ $Y=0.235 $X2=5.03 $Y2=0.39
r260 4 51 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.235 $X2=3.57 $Y2=0.39
r261 3 45 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.235 $X2=2.63 $Y2=0.39
r262 2 39 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r263 1 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_4%VGND 1 2 3 4 5 6 7 8 9 28 30 32 36 40 44 48
+ 52 56 60 63 64 66 67 69 70 72 73 75 76 78 79 80 107 108 114 119 122
r149 121 122 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=0.235
+ $X2=4.645 $Y2=0.235
r150 117 121 3.55086 $w=6.38e-07 $l=1.9e-07 $layer=LI1_cond $X=4.37 $Y=0.235
+ $X2=4.56 $Y2=0.235
r151 117 119 15.089 $w=6.38e-07 $l=4.15e-07 $layer=LI1_cond $X=4.37 $Y=0.235
+ $X2=3.955 $Y2=0.235
r152 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r153 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r154 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r155 105 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r156 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r157 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r158 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r159 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r160 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r161 96 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r162 96 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.37 $Y2=0
r163 95 122 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=4.645 $Y2=0
r164 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r165 92 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.37 $Y2=0
r166 91 119 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.91 $Y=0
+ $X2=3.955 $Y2=0
r167 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r168 88 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r169 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r170 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r171 85 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.15 $Y2=0
r172 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r173 82 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r174 82 84 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=2.07 $Y2=0
r175 80 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r176 80 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r177 78 104 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.235 $Y=0
+ $X2=8.05 $Y2=0
r178 78 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.235 $Y=0 $X2=8.32
+ $Y2=0
r179 77 107 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.405 $Y=0
+ $X2=8.51 $Y2=0
r180 77 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=0 $X2=8.32
+ $Y2=0
r181 75 101 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.295 $Y=0
+ $X2=7.13 $Y2=0
r182 75 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.295 $Y=0 $X2=7.38
+ $Y2=0
r183 74 104 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=7.465 $Y=0
+ $X2=8.05 $Y2=0
r184 74 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.465 $Y=0 $X2=7.38
+ $Y2=0
r185 72 98 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.355 $Y=0
+ $X2=6.21 $Y2=0
r186 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.355 $Y=0 $X2=6.44
+ $Y2=0
r187 71 101 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.525 $Y=0
+ $X2=7.13 $Y2=0
r188 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.525 $Y=0 $X2=6.44
+ $Y2=0
r189 69 95 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.415 $Y=0
+ $X2=5.29 $Y2=0
r190 69 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.415 $Y=0 $X2=5.5
+ $Y2=0
r191 68 98 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.585 $Y=0
+ $X2=6.21 $Y2=0
r192 68 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.585 $Y=0 $X2=5.5
+ $Y2=0
r193 66 87 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=2.99
+ $Y2=0
r194 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.1
+ $Y2=0
r195 65 91 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=3.91 $Y2=0
r196 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.1
+ $Y2=0
r197 63 84 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r198 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.16
+ $Y2=0
r199 62 87 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.99 $Y2=0
r200 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r201 58 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.32 $Y=0.085
+ $X2=8.32 $Y2=0
r202 58 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.32 $Y=0.085
+ $X2=8.32 $Y2=0.39
r203 54 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.38 $Y=0.085
+ $X2=7.38 $Y2=0
r204 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.38 $Y=0.085
+ $X2=7.38 $Y2=0.39
r205 50 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0
r206 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0.39
r207 46 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=0.085 $X2=5.5
+ $Y2=0
r208 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.5 $Y=0.085
+ $X2=5.5 $Y2=0.39
r209 42 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0
r210 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0.39
r211 38 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r212 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.39
r213 34 114 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r214 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r215 33 111 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r216 32 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r217 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=0.365 $Y2=0
r218 28 111 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r219 28 30 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r220 9 60 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.185
+ $Y=0.235 $X2=8.32 $Y2=0.39
r221 8 56 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.195
+ $Y=0.235 $X2=7.38 $Y2=0.39
r222 7 52 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.305
+ $Y=0.235 $X2=6.44 $Y2=0.39
r223 6 48 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.315
+ $Y=0.235 $X2=5.5 $Y2=0.39
r224 5 121 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=3.905
+ $Y=0.235 $X2=4.56 $Y2=0.39
r225 4 44 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.39
r226 3 40 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r227 2 36 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
r228 1 30 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

