* File: sky130_fd_sc_hdll__nand2_2.pxi.spice
* Created: Thu Aug 27 19:12:48 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2_2%B N_B_c_40_n N_B_M1001_g N_B_c_44_n N_B_M1000_g
+ N_B_c_45_n N_B_M1003_g N_B_c_41_n N_B_M1007_g B B N_B_c_43_n
+ PM_SKY130_FD_SC_HDLL__NAND2_2%B
x_PM_SKY130_FD_SC_HDLL__NAND2_2%A N_A_c_85_n N_A_M1002_g N_A_c_89_n N_A_M1004_g
+ N_A_c_90_n N_A_M1006_g N_A_c_86_n N_A_M1005_g A A N_A_c_88_n A
+ PM_SKY130_FD_SC_HDLL__NAND2_2%A
x_PM_SKY130_FD_SC_HDLL__NAND2_2%VPWR N_VPWR_M1000_d N_VPWR_M1003_d
+ N_VPWR_M1006_d N_VPWR_c_132_n N_VPWR_c_133_n N_VPWR_c_134_n N_VPWR_c_135_n
+ N_VPWR_c_136_n N_VPWR_c_137_n VPWR N_VPWR_c_138_n N_VPWR_c_131_n
+ N_VPWR_c_140_n N_VPWR_c_141_n PM_SKY130_FD_SC_HDLL__NAND2_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2_2%Y N_Y_M1002_d N_Y_M1000_s N_Y_M1004_s
+ N_Y_c_175_n N_Y_c_179_n N_Y_c_181_n N_Y_c_171_n N_Y_c_182_n Y Y Y N_Y_c_173_n
+ Y PM_SKY130_FD_SC_HDLL__NAND2_2%Y
x_PM_SKY130_FD_SC_HDLL__NAND2_2%A_27_47# N_A_27_47#_M1001_d N_A_27_47#_M1007_d
+ N_A_27_47#_M1005_s N_A_27_47#_c_225_n N_A_27_47#_c_231_n N_A_27_47#_c_226_n
+ N_A_27_47#_c_237_n N_A_27_47#_c_227_n N_A_27_47#_c_228_n
+ PM_SKY130_FD_SC_HDLL__NAND2_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND2_2%VGND N_VGND_M1001_s N_VGND_c_267_n VGND
+ N_VGND_c_268_n N_VGND_c_269_n N_VGND_c_270_n VGND
+ PM_SKY130_FD_SC_HDLL__NAND2_2%VGND
cc_1 VNB N_B_c_40_n 0.0228251f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B_c_41_n 0.01712f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB B 0.0134006f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_4 VNB N_B_c_43_n 0.0420212f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_5 VNB N_A_c_85_n 0.0170444f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_A_c_86_n 0.020726f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_7 VNB A 0.00358166f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_8 VNB N_A_c_88_n 0.0398557f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_9 VNB N_VPWR_c_131_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_Y_c_171_n 0.00313814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB Y 0.0152231f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.2
cc_12 VNB N_Y_c_173_n 8.47837e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_225_n 0.0183571f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_14 VNB N_A_27_47#_c_226_n 0.00969418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_227_n 0.00152046f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.202
cc_16 VNB N_A_27_47#_c_228_n 0.0113357f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_17 VNB N_VGND_c_267_n 0.00469188f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_18 VNB N_VGND_c_268_n 0.0505799f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.202
cc_19 VNB N_VGND_c_269_n 0.1766f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_20 VNB N_VGND_c_270_n 0.0217561f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_21 VPB N_B_c_44_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_22 VPB N_B_c_45_n 0.016445f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_23 VPB B 0.00508358f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_24 VPB N_B_c_43_n 0.0224377f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_25 VPB N_A_c_89_n 0.0164398f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_26 VPB N_A_c_90_n 0.0196229f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_27 VPB A 0.00252951f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_28 VPB N_A_c_88_n 0.0205086f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_29 VPB N_VPWR_c_132_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_30 VPB N_VPWR_c_133_n 0.0431773f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_31 VPB N_VPWR_c_134_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_135_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.16
cc_33 VPB N_VPWR_c_136_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_34 VPB N_VPWR_c_137_n 0.0314268f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.2
cc_35 VPB N_VPWR_c_138_n 0.0164632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_131_n 0.0572499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_140_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_141_n 0.00487897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB Y 0.00686757f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.2
cc_40 N_B_c_41_n N_A_c_85_n 0.0171699f $X=0.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_41 N_B_c_45_n N_A_c_89_n 0.0235349f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_42 B A 0.0210739f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_43 N_B_c_43_n A 0.00267039f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_44 N_B_c_43_n N_A_c_88_n 0.0171699f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_45 N_B_c_44_n N_VPWR_c_133_n 0.00779021f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_46 B N_VPWR_c_133_n 0.022009f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_47 N_B_c_44_n N_VPWR_c_134_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_48 N_B_c_45_n N_VPWR_c_134_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_49 N_B_c_45_n N_VPWR_c_135_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_50 N_B_c_44_n N_VPWR_c_131_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 N_B_c_45_n N_VPWR_c_131_n 0.011869f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_52 N_B_c_44_n N_Y_c_175_n 0.00347232f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_53 N_B_c_45_n N_Y_c_175_n 5.79575e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_54 B N_Y_c_175_n 0.0253353f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_55 N_B_c_43_n N_Y_c_175_n 0.00631893f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_56 N_B_c_44_n N_Y_c_179_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_57 N_B_c_45_n N_Y_c_179_n 0.0106251f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_58 N_B_c_45_n N_Y_c_181_n 0.0159475f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_59 N_B_c_45_n N_Y_c_182_n 6.49214e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_60 N_B_c_40_n N_A_27_47#_c_225_n 0.00681792f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_61 N_B_c_41_n N_A_27_47#_c_225_n 5.31865e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_62 N_B_c_40_n N_A_27_47#_c_231_n 0.00909307f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_63 N_B_c_41_n N_A_27_47#_c_231_n 0.00722146f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_64 B N_A_27_47#_c_231_n 0.0277091f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_65 N_B_c_43_n N_A_27_47#_c_231_n 0.00462292f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_66 N_B_c_40_n N_A_27_47#_c_226_n 8.92977e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_67 B N_A_27_47#_c_226_n 0.0240047f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_68 N_B_c_41_n N_A_27_47#_c_237_n 0.00388968f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_69 N_B_c_40_n N_A_27_47#_c_227_n 5.08193e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_70 N_B_c_41_n N_A_27_47#_c_227_n 0.00808249f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_71 N_B_c_40_n N_VGND_c_267_n 0.00382269f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_72 N_B_c_41_n N_VGND_c_267_n 0.00362559f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_73 N_B_c_41_n N_VGND_c_268_n 0.0039445f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_74 N_B_c_40_n N_VGND_c_269_n 0.00701584f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_75 N_B_c_41_n N_VGND_c_269_n 0.00582805f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_76 N_B_c_40_n N_VGND_c_270_n 0.00422241f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A_c_89_n N_VPWR_c_135_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_c_89_n N_VPWR_c_136_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_c_90_n N_VPWR_c_136_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_c_90_n N_VPWR_c_137_n 0.00724735f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_c_89_n N_VPWR_c_131_n 0.0100198f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_c_90_n N_VPWR_c_131_n 0.0131262f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_c_89_n N_Y_c_179_n 6.24674e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_89_n N_Y_c_181_n 0.0100617f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_85 A N_Y_c_181_n 0.0455963f $X=1.545 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_c_85_n N_Y_c_171_n 0.00386129f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_c_86_n N_Y_c_171_n 0.00620892f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_88 A N_Y_c_171_n 0.0245375f $X=1.545 $Y=1.105 $X2=0 $Y2=0
cc_89 N_A_c_88_n N_Y_c_171_n 0.00472855f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_90 N_A_c_89_n N_Y_c_182_n 0.0133069f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_c_90_n N_Y_c_182_n 0.0154666f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_c_85_n Y 4.37287e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_c_89_n Y 3.86571e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_c_90_n Y 0.00343963f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_c_86_n Y 0.00355723f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_96 A Y 0.0196442f $X=1.545 $Y=1.105 $X2=0 $Y2=0
cc_97 N_A_c_88_n Y 0.0189648f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_98 N_A_c_86_n N_Y_c_173_n 0.00679804f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_c_89_n Y 0.00225041f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_c_90_n Y 0.0168904f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_88_n Y 0.00616252f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_102 A N_A_27_47#_c_227_n 0.0145229f $X=1.545 $Y=1.105 $X2=0 $Y2=0
cc_103 N_A_c_85_n N_A_27_47#_c_228_n 0.0115551f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_c_86_n N_A_27_47#_c_228_n 0.00993842f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_105 A N_A_27_47#_c_228_n 0.00389697f $X=1.545 $Y=1.105 $X2=0 $Y2=0
cc_106 N_A_c_85_n N_VGND_c_268_n 0.00357877f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_c_86_n N_VGND_c_268_n 0.00357877f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_c_85_n N_VGND_c_269_n 0.005504f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_c_86_n N_VGND_c_269_n 0.00680287f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_110 N_VPWR_c_131_n N_Y_M1000_s 0.00231261f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_111 N_VPWR_c_131_n N_Y_M1004_s 0.00231261f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_112 N_VPWR_c_133_n N_Y_c_175_n 0.013769f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_113 N_VPWR_c_133_n N_Y_c_179_n 0.0615942f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_114 N_VPWR_c_134_n N_Y_c_179_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_115 N_VPWR_c_135_n N_Y_c_179_n 0.0385613f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_116 N_VPWR_c_131_n N_Y_c_179_n 0.0140101f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_117 N_VPWR_M1003_d N_Y_c_181_n 0.00362938f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_118 N_VPWR_c_135_n N_Y_c_181_n 0.0136682f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_119 N_VPWR_c_135_n N_Y_c_182_n 0.0470327f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_120 N_VPWR_c_136_n N_Y_c_182_n 0.0223557f $X=2.055 $Y=2.72 $X2=0 $Y2=0
cc_121 N_VPWR_c_137_n N_Y_c_182_n 0.0397449f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_122 N_VPWR_c_131_n N_Y_c_182_n 0.0140101f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_123 N_VPWR_M1006_d Y 9.41178e-19 $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_124 N_VPWR_M1006_d Y 0.0104004f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_125 N_VPWR_c_137_n Y 0.0141199f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_126 N_Y_c_173_n N_A_27_47#_M1005_s 0.0127474f $X=2.09 $Y=0.905 $X2=0 $Y2=0
cc_127 N_Y_c_181_n N_A_27_47#_c_231_n 0.00185835f $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_128 N_Y_c_181_n N_A_27_47#_c_227_n 0.00196249f $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_129 N_Y_M1002_d N_A_27_47#_c_228_n 0.00508491f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_130 N_Y_c_171_n N_A_27_47#_c_228_n 0.0270446f $X=1.95 $Y=0.78 $X2=0 $Y2=0
cc_131 N_Y_c_173_n N_A_27_47#_c_228_n 0.0172647f $X=2.09 $Y=0.905 $X2=0 $Y2=0
cc_132 N_Y_M1002_d N_VGND_c_269_n 0.00297142f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_231_n N_VGND_M1001_s 0.00583485f $X=0.985 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_27_47#_c_225_n N_VGND_c_267_n 0.017598f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_231_n N_VGND_c_267_n 0.0131159f $X=0.985 $Y=0.8 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_237_n N_VGND_c_267_n 0.0180776f $X=1.135 $Y=0.485 $X2=0
+ $Y2=0
cc_137 N_A_27_47#_c_227_n N_VGND_c_267_n 0.00436059f $X=1.135 $Y=0.715 $X2=0
+ $Y2=0
cc_138 N_A_27_47#_c_231_n N_VGND_c_268_n 0.00203275f $X=0.985 $Y=0.8 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_237_n N_VGND_c_268_n 0.0185715f $X=1.135 $Y=0.485 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_c_228_n N_VGND_c_268_n 0.0588959f $X=2.14 $Y=0.38 $X2=0 $Y2=0
cc_141 N_A_27_47#_M1001_d N_VGND_c_269_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_M1007_d N_VGND_c_269_n 0.00215206f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_M1005_s N_VGND_c_269_n 0.00209344f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_c_225_n N_VGND_c_269_n 0.012786f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_231_n N_VGND_c_269_n 0.0100794f $X=0.985 $Y=0.8 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_237_n N_VGND_c_269_n 0.0110923f $X=1.135 $Y=0.485 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_c_228_n N_VGND_c_269_n 0.0367278f $X=2.14 $Y=0.38 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_225_n N_VGND_c_270_n 0.0216446f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_231_n N_VGND_c_270_n 0.00271675f $X=0.985 $Y=0.8 $X2=0 $Y2=0
