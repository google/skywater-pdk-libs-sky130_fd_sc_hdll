* File: sky130_fd_sc_hdll__decap_6.pex.spice
* Created: Thu Aug 27 19:04:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DECAP_6%VGND 1 7 9 12 15 23 26 29
r22 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r23 26 28 0.445255 $w=8.22e-07 $l=3e-08 $layer=LI1_cond $X=2.5 $Y=0.385 $X2=2.53
+ $Y2=0.385
r24 21 23 0.900738 $w=1.219e-06 $l=9e-08 $layer=LI1_cond $X=0.647 $Y=0.385
+ $X2=0.647 $Y2=0.475
r25 20 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r26 17 21 3.85316 $w=1.219e-06 $l=3.85e-07 $layer=LI1_cond $X=0.647 $Y=0
+ $X2=0.647 $Y2=0.385
r27 17 20 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r28 13 23 8.15669 $w=1.219e-06 $l=8.15e-07 $layer=LI1_cond $X=0.647 $Y=1.29
+ $X2=0.647 $Y2=0.475
r29 12 15 21.4725 $w=1.706e-06 $l=8.8476e-07 $layer=POLY_cond $X=1.11 $Y=1.29
+ $X2=1.38 $Y2=2.05
r30 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.11
+ $Y=1.29 $X2=1.11 $Y2=1.29
r31 9 20 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r32 9 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r33 8 21 2.26174 $w=9.4e-07 $l=6.48e-07 $layer=LI1_cond $X=1.295 $Y=0.385
+ $X2=0.647 $Y2=0.385
r34 7 26 4.05283 $w=9.4e-07 $l=2.95e-07 $layer=LI1_cond $X=2.205 $Y=0.385
+ $X2=2.5 $Y2=0.385
r35 7 8 11.8106 $w=9.38e-07 $l=9.1e-07 $layer=LI1_cond $X=2.205 $Y=0.385
+ $X2=1.295 $Y2=0.385
r36 1 26 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=2.365 $Y=0.235
+ $X2=2.5 $Y2=0.475
r37 1 23 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.235 $X2=0.26 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HDLL__DECAP_6%VPWR 1 9 10 11 12 15 17 26 29
r23 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r24 26 28 0.218638 $w=1.674e-06 $l=3e-08 $layer=LI1_cond $X=2.5 $Y=1.915
+ $X2=2.53 $Y2=1.915
r25 20 23 0.323894 $w=1.13e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=2.175
+ $X2=0.26 $Y2=2.175
r26 16 26 2.18638 $w=1.674e-06 $l=3e-07 $layer=LI1_cond $X=2.2 $Y=1.915 $X2=2.5
+ $Y2=1.915
r27 15 17 36.3375 $w=1.17e-06 $l=7.15e-07 $layer=POLY_cond $X=2.2 $Y=0.69
+ $X2=1.485 $Y2=0.69
r28 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.2 $Y=1.11
+ $X2=2.2 $Y2=1.11
r29 12 29 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.53 $Y2=2.72
r30 12 20 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r31 11 23 4.56277 $w=1.26e-06 $l=4.55e-07 $layer=LI1_cond $X=0.715 $Y=2.175
+ $X2=0.26 $Y2=2.175
r32 10 16 6.13078 $w=1.674e-06 $l=8.55175e-07 $layer=LI1_cond $X=1.465 $Y=2.175
+ $X2=2.2 $Y2=1.915
r33 10 11 7.2619 $w=1.258e-06 $l=7.5e-07 $layer=LI1_cond $X=1.465 $Y=2.175
+ $X2=0.715 $Y2=2.175
r34 9 17 6.24815 $w=8.1e-07 $l=1.05e-07 $layer=POLY_cond $X=1.38 $Y=0.51
+ $X2=1.485 $Y2=0.51
r35 1 26 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=2.365
+ $Y=1.615 $X2=2.5 $Y2=1.83
r36 1 23 300 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=2 $X=2.365
+ $Y=1.615 $X2=0.26 $Y2=1.83
.ends

