* File: sky130_fd_sc_hdll__nor4_1.pex.spice
* Created: Thu Aug 27 19:16:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4_1%D 1 3 4 6 7 8 14
c28 4 0 7.47499e-20 $X=0.52 $Y=0.995
r29 14 15 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r30 12 14 32.4423 $w=3.64e-07 $l=2.45e-07 $layer=POLY_cond $X=0.25 $Y=1.202
+ $X2=0.495 $Y2=1.202
r31 7 8 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.21 $Y=1.16 $X2=0.21
+ $Y2=0.85
r32 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r33 4 15 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r35 1 14 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_1%C 1 3 4 6 7 11
c31 1 0 1.27256e-19 $X=0.99 $Y=0.995
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.16 $X2=1.05 $Y2=1.16
r33 7 11 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.125 $Y=1.53
+ $X2=1.125 $Y2=1.16
r34 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.05 $Y2=1.16
r35 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.015 $Y2=1.985
r36 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=1.05 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_1%B 1 3 4 6 7 11
r30 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.54
+ $Y=1.16 $X2=1.54 $Y2=1.16
r31 7 11 28.215 $w=2.88e-07 $l=7.1e-07 $layer=LI1_cond $X=1.6 $Y=1.87 $X2=1.6
+ $Y2=1.16
r32 4 10 50.6531 $w=2.63e-07 $l=2.69258e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.535 $Y2=1.16
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.495 $Y2=1.985
r34 1 10 39.0634 $w=2.63e-07 $l=1.94808e-07 $layer=POLY_cond $X=1.47 $Y=0.995
+ $X2=1.535 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.47 $Y=0.995 $X2=1.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_1%A 1 3 4 6 7
r26 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.02
+ $Y=1.16 $X2=2.02 $Y2=1.16
r27 7 11 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.07 $Y=0.85 $X2=2.07
+ $Y2=1.16
r28 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.985 $Y=1.41
+ $X2=2.02 $Y2=1.16
r29 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.985 $Y=1.41
+ $X2=1.985 $Y2=1.985
r30 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.96 $Y=0.995
+ $X2=2.02 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.96 $Y=0.995 $X2=1.96
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_1%Y 1 2 3 11 12 21 26 30
c42 21 0 1.27256e-19 $X=0.73 $Y=0.55
c43 12 0 7.47499e-20 $X=1.595 $Y=0.74
r44 30 35 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=0.257 $Y=2.21
+ $X2=0.257 $Y2=2.34
r45 26 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.68 $Y=0.55
+ $X2=1.68 $Y2=0.74
r46 23 24 3.50137 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.74
+ $X2=0.665 $Y2=0.825
r47 21 23 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=0.665 $Y=0.55
+ $X2=0.665 $Y2=0.74
r48 15 30 18.7487 $w=3.33e-07 $l=5.45e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=2.21
r49 13 23 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.815 $Y=0.74 $X2=0.665
+ $Y2=0.74
r50 12 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.595 $Y=0.74
+ $X2=1.68 $Y2=0.74
r51 12 13 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.595 $Y=0.74
+ $X2=0.815 $Y2=0.74
r52 11 15 25.3134 $w=1.68e-07 $l=3.88e-07 $layer=LI1_cond $X=0.645 $Y=1.58
+ $X2=0.257 $Y2=1.58
r53 11 24 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=0.645 $Y=1.495
+ $X2=0.645 $Y2=0.825
r54 3 35 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r55 3 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r56 2 26 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=1.545
+ $Y=0.235 $X2=1.68 $Y2=0.55
r57 1 21 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_1%VPWR 1 4 6 8 10 20
r27 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r28 17 20 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r29 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r30 12 16 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r31 10 19 5.13109 $w=1.7e-07 $l=3.12e-07 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.447 $Y2=2.72
r32 10 16 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.07 $Y2=2.72
r33 8 17 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r34 8 12 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r35 4 19 3.23982 $w=4e-07 $l=1.4854e-07 $layer=LI1_cond $X=2.335 $Y=2.635
+ $X2=2.447 $Y2=2.72
r36 4 6 18.295 $w=3.98e-07 $l=6.35e-07 $layer=LI1_cond $X=2.335 $Y=2.635
+ $X2=2.335 $Y2=2
r37 1 6 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.075
+ $Y=1.485 $X2=2.22 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_1%VGND 1 2 3 10 12 16 18 20 22 31 37 40
r45 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r46 37 39 9.93665 $w=4.42e-07 $l=4.48999e-07 $layer=LI1_cond $X=2.17 $Y=0.2
+ $X2=2.53 $Y2=0
r47 35 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r48 34 37 2.76018 $w=4.42e-07 $l=1e-07 $layer=LI1_cond $X=2.07 $Y=0.2 $X2=2.17
+ $Y2=0.2
r49 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r50 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r51 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r52 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r53 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r54 23 28 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r55 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r56 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r57 22 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r58 20 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r59 20 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r60 19 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.2
+ $Y2=0
r61 18 34 6.60399 $w=4.42e-07 $l=2.30217e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=2.07 $Y2=0.2
r62 18 19 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.365
+ $Y2=0
r63 14 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0
r64 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.39
r65 10 28 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r66 10 12 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.39
r67 3 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.035
+ $Y=0.235 $X2=2.17 $Y2=0.39
r68 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.39
r69 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

