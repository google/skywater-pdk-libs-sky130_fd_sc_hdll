* NGSPICE file created from sky130_fd_sc_hdll__ebufn_8.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__ebufn_8 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR TE_B a_437_309# VPB phighvt w=940000u l=180000u
+  ad=1.9584e+12p pd=1.56e+07u as=3.2075e+12p ps=2.41e+07u
M1001 VPWR TE_B a_437_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_437_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_437_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_485_47# a_124_297# Z VNB nshort w=650000u l=150000u
+  ad=2.106e+12p pd=1.818e+07u as=8.645e+11p ps=7.86e+06u
M1005 VPWR A a_124_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 a_437_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_321_47# TE_B VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=1.417e+12p ps=1.216e+07u
M1008 a_437_309# a_124_297# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1009 a_485_47# a_321_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_485_47# a_321_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_485_47# a_124_297# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR TE_B a_437_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_124_297# A VGND VNB nshort w=650000u l=150000u
+  ad=2.08e+11p pd=1.94e+06u as=0p ps=0u
M1014 a_321_47# TE_B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1015 Z a_124_297# a_437_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR TE_B a_437_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Z a_124_297# a_437_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_321_47# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_485_47# a_321_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_437_309# a_124_297# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_437_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_321_47# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Z a_124_297# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Z a_124_297# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_485_47# a_124_297# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND A a_124_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_485_47# a_124_297# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_437_309# a_124_297# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Z a_124_297# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_437_309# a_124_297# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Z a_124_297# a_437_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND a_321_47# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_124_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_321_47# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Z a_124_297# a_437_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_485_47# a_321_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Z a_124_297# a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

