* File: sky130_fd_sc_hdll__probe_p_8.pxi.spice
* Created: Wed Sep  2 08:50:27 2020
* 
x_PM_SKY130_FD_SC_HDLL__PROBE_P_8%A N_A_c_106_n N_A_M1001_g N_A_M1002_g
+ N_A_c_107_n N_A_M1009_g N_A_M1006_g N_A_M1015_g N_A_c_108_n N_A_M1019_g A
+ N_A_c_104_n N_A_c_105_n PM_SKY130_FD_SC_HDLL__PROBE_P_8%A
x_PM_SKY130_FD_SC_HDLL__PROBE_P_8%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1006_d
+ N_A_27_47#_M1001_d N_A_27_47#_M1009_d N_A_27_47#_c_194_n N_A_27_47#_M1000_g
+ N_A_27_47#_M1004_g N_A_27_47#_M1008_g N_A_27_47#_c_195_n N_A_27_47#_M1003_g
+ N_A_27_47#_c_196_n N_A_27_47#_M1005_g N_A_27_47#_M1011_g N_A_27_47#_M1013_g
+ N_A_27_47#_c_197_n N_A_27_47#_M1007_g N_A_27_47#_c_198_n N_A_27_47#_M1010_g
+ N_A_27_47#_M1016_g N_A_27_47#_M1018_g N_A_27_47#_c_199_n N_A_27_47#_M1012_g
+ N_A_27_47#_c_200_n N_A_27_47#_M1014_g N_A_27_47#_M1020_g N_A_27_47#_M1021_g
+ N_A_27_47#_c_201_n N_A_27_47#_M1017_g N_A_27_47#_c_202_n N_A_27_47#_c_381_p
+ N_A_27_47#_c_203_n N_A_27_47#_c_204_n N_A_27_47#_c_187_n N_A_27_47#_c_188_n
+ N_A_27_47#_c_226_n N_A_27_47#_c_285_p N_A_27_47#_c_189_n N_A_27_47#_c_190_n
+ N_A_27_47#_c_191_n N_A_27_47#_c_206_n N_A_27_47#_c_192_n N_A_27_47#_c_242_n
+ N_A_27_47#_c_193_n PM_SKY130_FD_SC_HDLL__PROBE_P_8%A_27_47#
x_PM_SKY130_FD_SC_HDLL__PROBE_P_8%VPWR N_VPWR_M1001_s N_VPWR_M1019_s
+ N_VPWR_M1003_s N_VPWR_M1007_s N_VPWR_M1012_s N_VPWR_M1017_s N_VPWR_c_453_n
+ N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n
+ N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n N_VPWR_c_463_n
+ N_VPWR_c_464_n VPWR VPWR N_VPWR_c_465_n N_VPWR_c_466_n N_VPWR_c_452_n
+ N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_470_n N_VPWR_c_471_n N_VPWR_c_472_n
+ PM_SKY130_FD_SC_HDLL__PROBE_P_8%VPWR
x_PM_SKY130_FD_SC_HDLL__PROBE_P_8%A_399_297# N_A_399_297#_M1004_s
+ N_A_399_297#_M1011_s N_A_399_297#_M1016_s N_A_399_297#_M1020_s
+ N_A_399_297#_M1000_d N_A_399_297#_M1005_d N_A_399_297#_M1010_d
+ N_A_399_297#_M1014_d N_A_399_297#_c_583_n N_A_399_297#_c_584_n
+ N_A_399_297#_c_563_n N_A_399_297#_c_564_n N_A_399_297#_c_571_n
+ N_A_399_297#_c_572_n N_A_399_297#_c_622_n N_A_399_297#_c_626_n
+ N_A_399_297#_c_565_n N_A_399_297#_c_573_n N_A_399_297#_c_638_n
+ N_A_399_297#_c_642_n N_A_399_297#_c_646_n N_A_399_297#_c_649_n
+ N_A_399_297#_c_566_n N_A_399_297#_c_574_n N_A_399_297#_c_575_n
+ N_A_399_297#_c_576_n N_A_399_297#_c_577_n N_A_399_297#_c_567_n
+ N_A_399_297#_c_568_n N_A_399_297#_c_580_n N_A_399_297#_R0_pos
+ N_A_399_297#_c_569_n N_A_399_297#_c_570_n
+ PM_SKY130_FD_SC_HDLL__PROBE_P_8%A_399_297#
x_PM_SKY130_FD_SC_HDLL__PROBE_P_8%VGND N_VGND_M1002_s N_VGND_M1015_s
+ N_VGND_M1008_d N_VGND_M1013_d N_VGND_M1018_d N_VGND_M1021_d N_VGND_c_804_n
+ N_VGND_c_805_n N_VGND_c_806_n N_VGND_c_807_n N_VGND_c_808_n N_VGND_c_809_n
+ N_VGND_c_810_n N_VGND_c_811_n N_VGND_c_812_n N_VGND_c_813_n N_VGND_c_814_n
+ VGND VGND N_VGND_c_815_n N_VGND_c_816_n N_VGND_c_817_n N_VGND_c_818_n
+ N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n N_VGND_c_823_n
+ VGND VGND PM_SKY130_FD_SC_HDLL__PROBE_P_8%VGND
x_PM_SKY130_FD_SC_HDLL__PROBE_P_8%X X N_X_R0_neg
+ PM_SKY130_FD_SC_HDLL__PROBE_P_8%X
cc_1 VNB N_A_M1002_g 0.0235699f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB N_A_M1006_g 0.0178195f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_3 VNB N_A_M1015_g 0.0175958f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.56
cc_4 VNB N_A_c_104_n 0.00806404f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_5 VNB N_A_c_105_n 0.0857159f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.212
cc_6 VNB N_A_27_47#_M1004_g 0.0179864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1008_g 0.0176972f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_8 VNB N_A_27_47#_M1011_g 0.0177101f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_9 VNB N_A_27_47#_M1013_g 0.0177101f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.175
cc_10 VNB N_A_27_47#_M1016_g 0.017668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1018_g 0.0175716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_M1020_g 0.0173202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_M1021_g 0.0237845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_187_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_188_n 0.00264995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_189_n 0.00459766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_190_n 0.00158168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_191_n 0.00478392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_192_n 0.00255533f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_193_n 0.232761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_452_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_399_297#_c_563_n 0.00224216f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.212
cc_23 VNB N_A_399_297#_c_564_n 0.00156403f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.212
cc_24 VNB N_A_399_297#_c_565_n 0.00224216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_399_297#_c_566_n 0.00156403f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_399_297#_c_567_n 0.00128099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_399_297#_c_568_n 0.00329069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_399_297#_c_569_n 0.00203863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_399_297#_c_570_n 0.0108695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_804_n 0.00473987f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_31 VNB N_VGND_c_805_n 0.0042804f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_32 VNB N_VGND_c_806_n 0.0173211f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.212
cc_33 VNB N_VGND_c_807_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_34 VNB N_VGND_c_808_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.212
cc_35 VNB N_VGND_c_809_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_810_n 0.0168835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_811_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_812_n 0.0328083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_813_n 0.0175114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_814_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_815_n 0.0155708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_816_n 0.0159859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_817_n 0.310169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_818_n 0.0182824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_819_n 0.00535855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_820_n 0.00573982f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_821_n 0.00515959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_822_n 0.00515959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_823_n 0.00515959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VPB N_A_c_106_n 0.0200897f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_51 VPB N_A_c_107_n 0.0158698f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_52 VPB N_A_c_108_n 0.0157116f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_53 VPB N_A_c_105_n 0.027794f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.212
cc_54 VPB N_A_27_47#_c_194_n 0.0159578f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_55 VPB N_A_27_47#_c_195_n 0.0156957f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.212
cc_56 VPB N_A_27_47#_c_196_n 0.0157094f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_57 VPB N_A_27_47#_c_197_n 0.0157094f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.175
cc_58 VPB N_A_27_47#_c_198_n 0.0157094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_199_n 0.0156687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_200_n 0.0155986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_47#_c_201_n 0.0207627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_47#_c_202_n 0.0331497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_203_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_47#_c_204_n 0.0107029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_47#_c_190_n 0.0037956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_206_n 0.00256136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_47#_c_193_n 0.0517345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_453_n 0.00466368f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_69 VPB N_VPWR_c_454_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_455_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_71 VPB N_VPWR_c_456_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.212
cc_72 VPB N_VPWR_c_457_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.212
cc_73 VPB N_VPWR_c_458_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.212
cc_74 VPB N_VPWR_c_459_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_460_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_461_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_462_n 0.0483898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_463_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_464_n 0.00574121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_465_n 0.0178692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_466_n 0.0143948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_452_n 0.056001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_468_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_469_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_470_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_471_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_472_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_399_297#_c_571_n 0.00189903f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.212
cc_89 VPB N_A_399_297#_c_572_n 0.00181449f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.175
cc_90 VPB N_A_399_297#_c_573_n 0.00189903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_399_297#_c_574_n 0.00181449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_399_297#_c_575_n 0.00180391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_399_297#_c_576_n 7.97535e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_399_297#_c_577_n 0.0040135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_399_297#_c_567_n 9.60741e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_399_297#_c_568_n 0.00354193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_399_297#_c_580_n 7.51087e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_399_297#_c_569_n 0.00228081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_399_297#_c_570_n 0.0109971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 N_A_c_108_n N_A_27_47#_c_194_n 0.0257643f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_M1015_g N_A_27_47#_M1004_g 0.0206671f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_102 N_A_c_106_n N_A_27_47#_c_202_n 0.0109826f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_107_n N_A_27_47#_c_202_n 7.3868e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_c_106_n N_A_27_47#_c_203_n 0.0137916f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_c_107_n N_A_27_47#_c_203_n 0.0137916f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_c_104_n N_A_27_47#_c_203_n 0.0576497f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_c_105_n N_A_27_47#_c_203_n 0.00720931f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_108 N_A_c_106_n N_A_27_47#_c_204_n 0.00138874f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A_c_104_n N_A_27_47#_c_204_n 0.0231493f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_c_105_n N_A_27_47#_c_204_n 0.00628911f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_111 N_A_M1002_g N_A_27_47#_c_187_n 0.0104513f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A_M1006_g N_A_27_47#_c_187_n 0.0104513f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_113 N_A_c_104_n N_A_27_47#_c_187_n 0.0563563f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_c_105_n N_A_27_47#_c_187_n 0.0031956f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_115 N_A_M1002_g N_A_27_47#_c_188_n 3.62277e-19 $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A_c_104_n N_A_27_47#_c_188_n 0.0243677f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_c_105_n N_A_27_47#_c_188_n 0.00751272f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_118 N_A_c_106_n N_A_27_47#_c_226_n 7.39465e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_107_n N_A_27_47#_c_226_n 0.0110586f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_108_n N_A_27_47#_c_226_n 0.0106665f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_M1006_g N_A_27_47#_c_189_n 0.00130233f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_122 N_A_M1015_g N_A_27_47#_c_189_n 0.00554622f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_123 N_A_c_105_n N_A_27_47#_c_189_n 0.00352603f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_124 N_A_c_107_n N_A_27_47#_c_190_n 3.85341e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_108_n N_A_27_47#_c_190_n 0.00167292f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_104_n N_A_27_47#_c_190_n 0.00212434f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_c_105_n N_A_27_47#_c_190_n 0.00874559f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_128 N_A_c_107_n N_A_27_47#_c_206_n 0.00109264f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_108_n N_A_27_47#_c_206_n 0.0123532f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_105_n N_A_27_47#_c_206_n 0.00789391f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_131 N_A_M1006_g N_A_27_47#_c_192_n 2.0357e-19 $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_132 N_A_M1015_g N_A_27_47#_c_192_n 0.0095971f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_133 N_A_c_105_n N_A_27_47#_c_192_n 0.00236691f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_134 N_A_c_104_n N_A_27_47#_c_242_n 0.0134383f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_105_n N_A_27_47#_c_242_n 0.00572689f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_136 N_A_c_105_n N_A_27_47#_c_193_n 0.0196732f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_137 N_A_c_106_n N_VPWR_c_453_n 0.00309049f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_107_n N_VPWR_c_453_n 0.00173895f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_107_n N_VPWR_c_454_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_108_n N_VPWR_c_454_n 0.00673617f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_108_n N_VPWR_c_455_n 0.00227804f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_106_n N_VPWR_c_465_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_106_n N_VPWR_c_452_n 0.0126298f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_107_n N_VPWR_c_452_n 0.0117184f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_108_n N_VPWR_c_452_n 0.0109026f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_M1015_g N_A_399_297#_c_583_n 8.35744e-19 $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_147 N_A_c_108_n N_A_399_297#_c_584_n 0.00131703f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_M1015_g N_A_399_297#_c_564_n 3.84696e-19 $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A_c_108_n N_A_399_297#_c_572_n 3.99559e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_M1006_g N_A_399_297#_c_567_n 4.35e-19 $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A_M1015_g N_A_399_297#_c_567_n 0.00330527f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A_c_108_n N_A_399_297#_c_567_n 0.00527173f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_104_n N_A_399_297#_c_567_n 0.00108623f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_c_105_n N_A_399_297#_c_567_n 0.00491141f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_155 N_A_M1006_g N_A_399_297#_c_568_n 6.36511e-19 $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A_M1015_g N_A_399_297#_c_568_n 0.00220756f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A_c_104_n N_A_399_297#_c_568_n 0.00120253f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_c_105_n N_A_399_297#_c_568_n 0.006144f $X=1.41 $Y=1.212 $X2=0 $Y2=0
cc_159 N_A_M1002_g N_VGND_c_804_n 0.00307766f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A_M1006_g N_VGND_c_804_n 0.00165775f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_161 N_A_M1015_g N_VGND_c_805_n 0.00175184f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A_M1006_g N_VGND_c_815_n 0.00439206f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_163 N_A_M1015_g N_VGND_c_815_n 0.00439206f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_164 N_A_M1002_g N_VGND_c_817_n 0.00696186f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_165 N_A_M1006_g N_VGND_c_817_n 0.00596299f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_166 N_A_M1015_g N_VGND_c_817_n 0.00586743f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A_M1002_g N_VGND_c_818_n 0.00439206f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A_c_108_n X 0.00208546f $X=1.435 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_169 N_A_27_47#_c_203_n N_VPWR_M1001_s 0.00209407f $X=1.035 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_170 N_A_27_47#_c_206_n N_VPWR_M1019_s 0.00168556f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_203_n N_VPWR_c_453_n 0.0118222f $X=1.035 $Y=1.53 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_226_n N_VPWR_c_454_n 0.0189467f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_194_n N_VPWR_c_455_n 0.00227804f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_226_n N_VPWR_c_455_n 0.0303035f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_191_n N_VPWR_c_455_n 0.00624749f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_206_n N_VPWR_c_455_n 0.00246523f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_194_n N_VPWR_c_456_n 0.00673617f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_195_n N_VPWR_c_456_n 0.00673617f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_195_n N_VPWR_c_457_n 0.00227804f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_196_n N_VPWR_c_457_n 0.00227804f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_196_n N_VPWR_c_458_n 0.00673617f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_197_n N_VPWR_c_458_n 0.00673617f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_197_n N_VPWR_c_459_n 0.00227804f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_198_n N_VPWR_c_459_n 0.00227804f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_198_n N_VPWR_c_460_n 0.00673617f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_199_n N_VPWR_c_460_n 0.00673617f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_199_n N_VPWR_c_461_n 0.00173895f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_200_n N_VPWR_c_461_n 0.00173895f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_193_n N_VPWR_c_461_n 9.15469e-19 $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_201_n N_VPWR_c_462_n 0.00356412f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_200_n N_VPWR_c_463_n 0.00673617f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_201_n N_VPWR_c_463_n 0.00673617f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_202_n N_VPWR_c_465_n 0.0210596f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_194 N_A_27_47#_M1001_d N_VPWR_c_452_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_M1009_d N_VPWR_c_452_n 0.00228158f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_194_n N_VPWR_c_452_n 0.0109073f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_195_n N_VPWR_c_452_n 0.010882f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_196_n N_VPWR_c_452_n 0.010882f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_197_n N_VPWR_c_452_n 0.010882f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_198_n N_VPWR_c_452_n 0.010882f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_199_n N_VPWR_c_452_n 0.0116092f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_200_n N_VPWR_c_452_n 0.0117593f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_201_n N_VPWR_c_452_n 0.0128506f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_202_n N_VPWR_c_452_n 0.0124725f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_226_n N_VPWR_c_452_n 0.0123132f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_206 N_A_27_47#_M1004_g N_A_399_297#_c_583_n 0.00676782f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_M1008_g N_A_399_297#_c_583_n 0.00667323f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_M1011_g N_A_399_297#_c_583_n 8.18986e-19 $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_285_p N_A_399_297#_c_583_n 0.00463764f $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_194_n N_A_399_297#_c_584_n 0.0119593f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_195_n N_A_399_297#_c_584_n 0.0119593f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_196_n N_A_399_297#_c_584_n 0.00131703f $X=2.845 $Y=1.41
+ $X2=0 $Y2=0
cc_213 N_A_27_47#_c_226_n N_A_399_297#_c_584_n 0.00539931f $X=1.2 $Y=1.63 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_M1008_g N_A_399_297#_c_563_n 0.00865867f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_M1011_g N_A_399_297#_c_563_n 0.00865867f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_191_n N_A_399_297#_c_563_n 0.0448129f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_193_n N_A_399_297#_c_563_n 0.00426451f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_218 N_A_27_47#_M1004_g N_A_399_297#_c_564_n 0.00280547f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_M1008_g N_A_399_297#_c_564_n 9.9253e-19 $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_191_n N_A_399_297#_c_564_n 0.0264527f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_192_n N_A_399_297#_c_564_n 0.00738314f $X=1.507 $Y=0.82
+ $X2=0 $Y2=0
cc_222 N_A_27_47#_c_193_n N_A_399_297#_c_564_n 0.00208213f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_223 N_A_27_47#_c_195_n N_A_399_297#_c_571_n 0.0127878f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_196_n N_A_399_297#_c_571_n 0.0127878f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_191_n N_A_399_297#_c_571_n 0.0388326f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_193_n N_A_399_297#_c_571_n 0.00682853f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_227 N_A_27_47#_c_194_n N_A_399_297#_c_572_n 0.00393265f $X=1.905 $Y=1.41
+ $X2=0 $Y2=0
cc_228 N_A_27_47#_c_195_n N_A_399_297#_c_572_n 0.00194892f $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_229 N_A_27_47#_c_191_n N_A_399_297#_c_572_n 0.0232731f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_206_n N_A_399_297#_c_572_n 0.00741886f $X=1.507 $Y=1.53
+ $X2=0 $Y2=0
cc_231 N_A_27_47#_c_193_n N_A_399_297#_c_572_n 0.00744602f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_232 N_A_27_47#_M1008_g N_A_399_297#_c_622_n 8.18986e-19 $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_M1011_g N_A_399_297#_c_622_n 0.00667323f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_M1013_g N_A_399_297#_c_622_n 0.00667323f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_M1016_g N_A_399_297#_c_622_n 8.18986e-19 $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_195_n N_A_399_297#_c_626_n 0.00131703f $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_237 N_A_27_47#_c_196_n N_A_399_297#_c_626_n 0.0119593f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_197_n N_A_399_297#_c_626_n 0.0119593f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_198_n N_A_399_297#_c_626_n 0.00131703f $X=3.785 $Y=1.41
+ $X2=0 $Y2=0
cc_240 N_A_27_47#_M1013_g N_A_399_297#_c_565_n 0.00865867f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_M1016_g N_A_399_297#_c_565_n 0.00865867f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_191_n N_A_399_297#_c_565_n 0.0435848f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_193_n N_A_399_297#_c_565_n 0.00395902f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_244 N_A_27_47#_c_197_n N_A_399_297#_c_573_n 0.0127878f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_198_n N_A_399_297#_c_573_n 0.0127878f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_191_n N_A_399_297#_c_573_n 0.0373193f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_193_n N_A_399_297#_c_573_n 0.00571893f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_248 N_A_27_47#_M1013_g N_A_399_297#_c_638_n 8.18986e-19 $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_M1016_g N_A_399_297#_c_638_n 0.00667323f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_M1018_g N_A_399_297#_c_638_n 0.00672216f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_M1020_g N_A_399_297#_c_638_n 8.29189e-19 $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_197_n N_A_399_297#_c_642_n 0.00131703f $X=3.315 $Y=1.41
+ $X2=0 $Y2=0
cc_253 N_A_27_47#_c_198_n N_A_399_297#_c_642_n 0.0119593f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_199_n N_A_399_297#_c_642_n 0.0121815f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_200_n N_A_399_297#_c_642_n 0.00134414f $X=4.725 $Y=1.41
+ $X2=0 $Y2=0
cc_256 N_A_27_47#_M1018_g N_A_399_297#_c_646_n 5.26907e-19 $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1020_g N_A_399_297#_c_646_n 0.00682312f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1021_g N_A_399_297#_c_646_n 0.00550646f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_199_n N_A_399_297#_c_649_n 7.3868e-19 $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_200_n N_A_399_297#_c_649_n 0.0125412f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_201_n N_A_399_297#_c_649_n 0.0110847f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_M1011_g N_A_399_297#_c_566_n 0.0010041f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1013_g N_A_399_297#_c_566_n 0.0010041f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_191_n N_A_399_297#_c_566_n 0.0264527f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_193_n N_A_399_297#_c_566_n 0.00208213f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_266 N_A_27_47#_c_196_n N_A_399_297#_c_574_n 0.00196122f $X=2.845 $Y=1.41
+ $X2=0 $Y2=0
cc_267 N_A_27_47#_c_197_n N_A_399_297#_c_574_n 0.00196122f $X=3.315 $Y=1.41
+ $X2=0 $Y2=0
cc_268 N_A_27_47#_c_191_n N_A_399_297#_c_574_n 0.0232731f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_193_n N_A_399_297#_c_574_n 0.00744602f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_270 N_A_27_47#_c_191_n N_A_399_297#_c_575_n 0.00390977f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_193_n N_A_399_297#_c_575_n 0.0035502f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_193_n N_A_399_297#_c_576_n 0.021313f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_191_n N_A_399_297#_c_577_n 0.0182232f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_193_n N_A_399_297#_c_577_n 0.0162832f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_194_n N_A_399_297#_c_567_n 0.00286939f $X=1.905 $Y=1.41
+ $X2=0 $Y2=0
cc_276 N_A_27_47#_M1004_g N_A_399_297#_c_567_n 0.00244189f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_M1008_g N_A_399_297#_c_567_n 0.00195011f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_195_n N_A_399_297#_c_567_n 0.0022851f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_196_n N_A_399_297#_c_567_n 0.00227229f $X=2.845 $Y=1.41
+ $X2=0 $Y2=0
cc_280 N_A_27_47#_M1011_g N_A_399_297#_c_567_n 0.00195011f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_M1013_g N_A_399_297#_c_567_n 0.00195011f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_197_n N_A_399_297#_c_567_n 0.00227229f $X=3.315 $Y=1.41
+ $X2=0 $Y2=0
cc_283 N_A_27_47#_c_198_n N_A_399_297#_c_567_n 0.00220812f $X=3.785 $Y=1.41
+ $X2=0 $Y2=0
cc_284 N_A_27_47#_M1016_g N_A_399_297#_c_567_n 0.00169093f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_M1018_g N_A_399_297#_c_567_n 5.80122e-19 $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_226_n N_A_399_297#_c_567_n 0.00151366f $X=1.2 $Y=1.63 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_285_p N_A_399_297#_c_567_n 3.62377e-19 $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_189_n N_A_399_297#_c_567_n 0.00248095f $X=1.507 $Y=1.075
+ $X2=0 $Y2=0
cc_289 N_A_27_47#_c_190_n N_A_399_297#_c_567_n 0.00275103f $X=1.507 $Y=1.445
+ $X2=0 $Y2=0
cc_290 N_A_27_47#_c_191_n N_A_399_297#_c_567_n 0.00898621f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_206_n N_A_399_297#_c_567_n 0.00410518f $X=1.507 $Y=1.53
+ $X2=0 $Y2=0
cc_292 N_A_27_47#_c_192_n N_A_399_297#_c_567_n 0.00346878f $X=1.507 $Y=0.82
+ $X2=0 $Y2=0
cc_293 N_A_27_47#_c_242_n N_A_399_297#_c_567_n 3.47197e-19 $X=1.507 $Y=1.16
+ $X2=0 $Y2=0
cc_294 N_A_27_47#_c_193_n N_A_399_297#_c_567_n 0.00637434f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_295 N_A_27_47#_M1004_g N_A_399_297#_c_568_n 0.00181926f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_M1008_g N_A_399_297#_c_568_n 0.00180868f $X=2.35 $Y=0.56 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_M1011_g N_A_399_297#_c_568_n 0.00180868f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1013_g N_A_399_297#_c_568_n 0.00180868f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1016_g N_A_399_297#_c_568_n 0.00180868f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_M1018_g N_A_399_297#_c_568_n 0.00583367f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_199_n N_A_399_297#_c_568_n 0.00557969f $X=4.255 $Y=1.41
+ $X2=0 $Y2=0
cc_302 N_A_27_47#_c_200_n N_A_399_297#_c_568_n 5.1886e-19 $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_M1020_g N_A_399_297#_c_568_n 4.43043e-19 $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_202_n N_A_399_297#_c_568_n 6.39042e-19 $X=0.26 $Y=1.63 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_381_p N_A_399_297#_c_568_n 5.26298e-19 $X=0.31 $Y=0.42 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_226_n N_A_399_297#_c_568_n 0.00612748f $X=1.2 $Y=1.63 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_285_p N_A_399_297#_c_568_n 0.00465676f $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_206_n N_A_399_297#_c_568_n 0.0036003f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_192_n N_A_399_297#_c_568_n 0.00356332f $X=1.507 $Y=0.82
+ $X2=0 $Y2=0
cc_310 N_A_27_47#_c_193_n N_A_399_297#_c_568_n 0.00254015f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_c_191_n N_A_399_297#_c_580_n 0.00312295f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_193_n N_A_399_297#_c_580_n 0.00745114f $X=5.17 $Y=1.217
+ $X2=0 $Y2=0
cc_313 N_A_27_47#_c_198_n N_A_399_297#_c_569_n 0.00196122f $X=3.785 $Y=1.41
+ $X2=0 $Y2=0
cc_314 N_A_27_47#_M1016_g N_A_399_297#_c_569_n 0.00132485f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_M1018_g N_A_399_297#_c_569_n 0.0129266f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_199_n N_A_399_297#_c_569_n 0.0149796f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_200_n N_A_399_297#_c_569_n 0.0135468f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_M1020_g N_A_399_297#_c_569_n 0.01178f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_M1021_g N_A_399_297#_c_569_n 0.00986498f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_201_n N_A_399_297#_c_569_n 0.00677208f $X=5.195 $Y=1.41
+ $X2=0 $Y2=0
cc_321 N_A_27_47#_c_191_n N_A_399_297#_c_569_n 0.0346951f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_193_n N_A_399_297#_c_569_n 0.0753261f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_M1013_g N_A_399_297#_c_570_n 2.46205e-19 $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_M1016_g N_A_399_297#_c_570_n 0.00351582f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1018_g N_A_399_297#_c_570_n 2.47268e-19 $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_191_n N_A_399_297#_c_570_n 0.00349157f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_193_n N_A_399_297#_c_570_n 0.0101569f $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_187_n N_VGND_M1002_s 0.00213931f $X=1.065 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_329 N_A_27_47#_c_192_n N_VGND_M1015_s 0.0022207f $X=1.507 $Y=0.82 $X2=0 $Y2=0
cc_330 N_A_27_47#_c_187_n N_VGND_c_804_n 0.0161649f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_331 N_A_27_47#_M1004_g N_VGND_c_805_n 0.0016904f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_332 N_A_27_47#_c_285_p N_VGND_c_805_n 0.0126187f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_333 N_A_27_47#_c_191_n N_VGND_c_805_n 0.00749407f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A_27_47#_c_192_n N_VGND_c_805_n 0.00588718f $X=1.507 $Y=0.82 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_M1004_g N_VGND_c_806_n 0.00541359f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_336 N_A_27_47#_M1008_g N_VGND_c_806_n 0.00424416f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_337 N_A_27_47#_M1008_g N_VGND_c_807_n 0.0016763f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_338 N_A_27_47#_M1011_g N_VGND_c_807_n 0.0016763f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_339 N_A_27_47#_M1011_g N_VGND_c_808_n 0.00424416f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_340 N_A_27_47#_M1013_g N_VGND_c_808_n 0.00424416f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_341 N_A_27_47#_M1013_g N_VGND_c_809_n 0.0016763f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_342 N_A_27_47#_M1016_g N_VGND_c_809_n 0.0016763f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_343 N_A_27_47#_M1016_g N_VGND_c_810_n 0.00424416f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_344 N_A_27_47#_M1018_g N_VGND_c_810_n 0.00472104f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_345 N_A_27_47#_M1018_g N_VGND_c_811_n 0.00166854f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_346 N_A_27_47#_M1020_g N_VGND_c_811_n 0.00166854f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_347 N_A_27_47#_c_193_n N_VGND_c_811_n 7.95874e-19 $X=5.17 $Y=1.217 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_M1021_g N_VGND_c_812_n 0.00321269f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_349 N_A_27_47#_M1020_g N_VGND_c_813_n 0.00472104f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_350 N_A_27_47#_M1021_g N_VGND_c_813_n 0.00541359f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_351 N_A_27_47#_c_187_n N_VGND_c_815_n 0.00515628f $X=1.065 $Y=0.82 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_285_p N_VGND_c_815_n 0.0146703f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_353 N_A_27_47#_M1002_d N_VGND_c_817_n 0.00288496f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_M1006_d N_VGND_c_817_n 0.00212429f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_M1004_g N_VGND_c_817_n 0.00905719f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_27_47#_M1008_g N_VGND_c_817_n 0.00573509f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_27_47#_M1011_g N_VGND_c_817_n 0.00573509f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A_27_47#_M1013_g N_VGND_c_817_n 0.00573509f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A_27_47#_M1016_g N_VGND_c_817_n 0.0053659f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_27_47#_M1018_g N_VGND_c_817_n 0.00739652f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_27_47#_M1020_g N_VGND_c_817_n 0.0075548f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A_27_47#_M1021_g N_VGND_c_817_n 0.0108276f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A_27_47#_c_381_p N_VGND_c_817_n 0.0114629f $X=0.31 $Y=0.42 $X2=0 $Y2=0
cc_364 N_A_27_47#_c_187_n N_VGND_c_817_n 0.0119645f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_365 N_A_27_47#_c_285_p N_VGND_c_817_n 0.0102294f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_366 N_A_27_47#_c_192_n N_VGND_c_817_n 3.25202e-19 $X=1.507 $Y=0.82 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_381_p N_VGND_c_818_n 0.0189483f $X=0.31 $Y=0.42 $X2=0 $Y2=0
cc_368 N_A_27_47#_c_187_n N_VGND_c_818_n 0.002104f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_369 N_A_27_47#_c_194_n X 0.00208546f $X=1.905 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_370 N_A_27_47#_c_195_n X 0.00208546f $X=2.375 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_371 N_A_27_47#_c_196_n X 0.00208546f $X=2.845 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_372 N_A_27_47#_c_197_n X 0.00208546f $X=3.315 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_373 N_A_27_47#_c_198_n X 0.00208546f $X=3.785 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_374 N_A_27_47#_c_199_n X 0.00427677f $X=4.255 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_375 N_A_27_47#_c_226_n X 0.00522195f $X=1.2 $Y=1.63 $X2=-0.19 $Y2=-0.24
cc_376 N_VPWR_c_452_n N_A_399_297#_M1000_d 0.00203508f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_452_n N_A_399_297#_M1005_d 0.00203508f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_452_n N_A_399_297#_M1010_d 0.00204531f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_452_n N_A_399_297#_M1014_d 0.00232867f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_455_n N_A_399_297#_c_584_n 0.030305f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_381 N_VPWR_c_456_n N_A_399_297#_c_584_n 0.0190121f $X=2.475 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_457_n N_A_399_297#_c_584_n 0.030305f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_383 N_VPWR_c_452_n N_A_399_297#_c_584_n 0.0124581f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_384 N_VPWR_M1003_s N_A_399_297#_c_571_n 0.00156212f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_457_n N_A_399_297#_c_571_n 0.0149094f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_386 N_VPWR_c_457_n N_A_399_297#_c_626_n 0.030305f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_387 N_VPWR_c_458_n N_A_399_297#_c_626_n 0.0190121f $X=3.415 $Y=2.72 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_459_n N_A_399_297#_c_626_n 0.030305f $X=3.55 $Y=2 $X2=0 $Y2=0
cc_389 N_VPWR_c_452_n N_A_399_297#_c_626_n 0.0124581f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_390 N_VPWR_M1007_s N_A_399_297#_c_573_n 0.00156212f $X=3.405 $Y=1.485 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_459_n N_A_399_297#_c_573_n 0.0149094f $X=3.55 $Y=2 $X2=0 $Y2=0
cc_392 N_VPWR_c_459_n N_A_399_297#_c_642_n 0.030305f $X=3.55 $Y=2 $X2=0 $Y2=0
cc_393 N_VPWR_c_460_n N_A_399_297#_c_642_n 0.0190121f $X=4.355 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_452_n N_A_399_297#_c_642_n 0.0124581f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_463_n N_A_399_297#_c_649_n 0.0190121f $X=5.295 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_452_n N_A_399_297#_c_649_n 0.0124581f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_461_n N_A_399_297#_c_576_n 0.00125602f $X=4.49 $Y=2 $X2=0 $Y2=0
cc_398 N_VPWR_c_455_n N_A_399_297#_c_567_n 0.00434171f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_399 N_VPWR_c_457_n N_A_399_297#_c_567_n 0.00397614f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_400 N_VPWR_c_459_n N_A_399_297#_c_567_n 0.00394775f $X=3.55 $Y=2 $X2=0 $Y2=0
cc_401 N_VPWR_c_452_n N_A_399_297#_c_567_n 0.0465657f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_453_n N_A_399_297#_c_568_n 2.77994e-19 $X=0.73 $Y=2 $X2=0 $Y2=0
cc_403 N_VPWR_c_455_n N_A_399_297#_c_568_n 2.82168e-19 $X=1.67 $Y=2 $X2=0 $Y2=0
cc_404 N_VPWR_c_457_n N_A_399_297#_c_568_n 2.82168e-19 $X=2.61 $Y=2 $X2=0 $Y2=0
cc_405 N_VPWR_c_459_n N_A_399_297#_c_568_n 2.82168e-19 $X=3.55 $Y=2 $X2=0 $Y2=0
cc_406 N_VPWR_c_461_n N_A_399_297#_c_568_n 6.38767e-19 $X=4.49 $Y=2 $X2=0 $Y2=0
cc_407 N_VPWR_c_462_n N_A_399_297#_c_568_n 2.81286e-19 $X=5.43 $Y=1.66 $X2=0
+ $Y2=0
cc_408 N_VPWR_M1012_s N_A_399_297#_c_569_n 0.00218233f $X=4.345 $Y=1.485 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_461_n N_A_399_297#_c_569_n 0.0123277f $X=4.49 $Y=2 $X2=0 $Y2=0
cc_410 N_VPWR_c_462_n N_VGND_c_812_n 0.00782513f $X=5.43 $Y=1.66 $X2=0 $Y2=0
cc_411 N_VPWR_M1019_s X 2.64944e-19 $X=1.525 $Y=1.485 $X2=-0.19 $Y2=-0.24
cc_412 N_VPWR_M1003_s X 2.64944e-19 $X=2.465 $Y=1.485 $X2=-0.19 $Y2=-0.24
cc_413 N_VPWR_M1007_s X 2.64944e-19 $X=3.405 $Y=1.485 $X2=-0.19 $Y2=-0.24
cc_414 N_VPWR_c_453_n X 5.32599e-19 $X=0.73 $Y=2 $X2=-0.19 $Y2=-0.24
cc_415 N_VPWR_c_455_n X 0.00447217f $X=1.67 $Y=2 $X2=-0.19 $Y2=-0.24
cc_416 N_VPWR_c_457_n X 0.00447217f $X=2.61 $Y=2 $X2=-0.19 $Y2=-0.24
cc_417 N_VPWR_c_459_n X 0.00447217f $X=3.55 $Y=2 $X2=-0.19 $Y2=-0.24
cc_418 N_VPWR_c_461_n X 0.00122421f $X=4.49 $Y=2 $X2=-0.19 $Y2=-0.24
cc_419 N_VPWR_c_452_n X 0.0375576f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_420 N_A_399_297#_c_567_n N_VGND_M1015_s 0.00417198f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_421 N_A_399_297#_c_568_n N_VGND_M1015_s 0.00132928f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_422 N_A_399_297#_c_563_n N_VGND_M1008_d 0.00204876f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_423 N_A_399_297#_c_567_n N_VGND_M1008_d 0.00417198f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_424 N_A_399_297#_c_568_n N_VGND_M1008_d 0.0019335f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_425 N_A_399_297#_c_565_n N_VGND_M1013_d 0.00204876f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_426 N_A_399_297#_c_567_n N_VGND_M1013_d 0.00417198f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_427 N_A_399_297#_c_568_n N_VGND_M1013_d 0.0019335f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_428 N_A_399_297#_c_569_n N_VGND_M1018_d 0.00282836f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_429 N_A_399_297#_c_583_n N_VGND_c_805_n 0.0117379f $X=2.14 $Y=0.42 $X2=0
+ $Y2=0
cc_430 N_A_399_297#_c_567_n N_VGND_c_805_n 0.0026606f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_431 N_A_399_297#_c_568_n N_VGND_c_805_n 0.00519536f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_432 N_A_399_297#_c_583_n N_VGND_c_806_n 0.0188551f $X=2.14 $Y=0.42 $X2=0
+ $Y2=0
cc_433 N_A_399_297#_c_563_n N_VGND_c_806_n 0.00289562f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_434 N_A_399_297#_c_583_n N_VGND_c_807_n 0.0117367f $X=2.14 $Y=0.42 $X2=0
+ $Y2=0
cc_435 N_A_399_297#_c_563_n N_VGND_c_807_n 0.021547f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_436 N_A_399_297#_c_622_n N_VGND_c_807_n 0.0117367f $X=3.08 $Y=0.42 $X2=0
+ $Y2=0
cc_437 N_A_399_297#_c_567_n N_VGND_c_807_n 0.00215981f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_438 N_A_399_297#_c_568_n N_VGND_c_807_n 0.00445215f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_439 N_A_399_297#_c_563_n N_VGND_c_808_n 0.00289562f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_440 N_A_399_297#_c_622_n N_VGND_c_808_n 0.0188551f $X=3.08 $Y=0.42 $X2=0
+ $Y2=0
cc_441 N_A_399_297#_c_565_n N_VGND_c_808_n 0.00289562f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_442 N_A_399_297#_c_622_n N_VGND_c_809_n 0.0117367f $X=3.08 $Y=0.42 $X2=0
+ $Y2=0
cc_443 N_A_399_297#_c_565_n N_VGND_c_809_n 0.021547f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_444 N_A_399_297#_c_638_n N_VGND_c_809_n 0.0117367f $X=4.02 $Y=0.42 $X2=0
+ $Y2=0
cc_445 N_A_399_297#_c_567_n N_VGND_c_809_n 0.00215981f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_446 N_A_399_297#_c_568_n N_VGND_c_809_n 0.00445215f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_447 N_A_399_297#_c_565_n N_VGND_c_810_n 0.00289562f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_448 N_A_399_297#_c_638_n N_VGND_c_810_n 0.0188551f $X=4.02 $Y=0.42 $X2=0
+ $Y2=0
cc_449 N_A_399_297#_c_569_n N_VGND_c_810_n 0.0015162f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_450 N_A_399_297#_c_576_n N_VGND_c_811_n 0.00113651f $X=5.005 $Y=1.19 $X2=0
+ $Y2=0
cc_451 N_A_399_297#_c_569_n N_VGND_c_811_n 0.0214341f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_452 N_A_399_297#_c_568_n N_VGND_c_812_n 3.21297e-19 $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_453 N_A_399_297#_c_646_n N_VGND_c_813_n 0.0189039f $X=4.96 $Y=0.42 $X2=0
+ $Y2=0
cc_454 N_A_399_297#_c_569_n N_VGND_c_813_n 0.0013974f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_455 N_A_399_297#_M1004_s N_VGND_c_817_n 0.00187087f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_A_399_297#_M1011_s N_VGND_c_817_n 0.00187087f $X=2.945 $Y=0.235 $X2=0
+ $Y2=0
cc_457 N_A_399_297#_M1016_s N_VGND_c_817_n 0.00144642f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_458 N_A_399_297#_M1020_s N_VGND_c_817_n 0.00215201f $X=4.825 $Y=0.235 $X2=0
+ $Y2=0
cc_459 N_A_399_297#_c_583_n N_VGND_c_817_n 0.0122069f $X=2.14 $Y=0.42 $X2=0
+ $Y2=0
cc_460 N_A_399_297#_c_563_n N_VGND_c_817_n 0.00852807f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_461 N_A_399_297#_c_622_n N_VGND_c_817_n 0.0122069f $X=3.08 $Y=0.42 $X2=0
+ $Y2=0
cc_462 N_A_399_297#_c_565_n N_VGND_c_817_n 0.00852807f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_463 N_A_399_297#_c_638_n N_VGND_c_817_n 0.0122069f $X=4.02 $Y=0.42 $X2=0
+ $Y2=0
cc_464 N_A_399_297#_c_646_n N_VGND_c_817_n 0.0122217f $X=4.96 $Y=0.42 $X2=0
+ $Y2=0
cc_465 N_A_399_297#_c_567_n N_VGND_c_817_n 0.051254f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_466 N_A_399_297#_c_568_n N_VGND_c_817_n 0.0528267f $X=3.56 $Y=1.27 $X2=0
+ $Y2=0
cc_467 N_A_399_297#_c_580_n N_VGND_c_817_n 0.0119699f $X=3.985 $Y=1.19 $X2=0
+ $Y2=0
cc_468 N_A_399_297#_c_569_n N_VGND_c_817_n 0.0070103f $X=4.96 $Y=1.175 $X2=0
+ $Y2=0
cc_469 N_A_399_297#_c_584_n X 0.00499989f $X=2.14 $Y=1.755 $X2=-0.19 $Y2=-0.24
cc_470 N_A_399_297#_c_626_n X 0.00499989f $X=3.08 $Y=1.755 $X2=-0.19 $Y2=-0.24
cc_471 N_A_399_297#_c_642_n X 0.0047356f $X=4.02 $Y=1.755 $X2=-0.19 $Y2=-0.24
