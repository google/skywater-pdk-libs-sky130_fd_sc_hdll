* File: sky130_fd_sc_hdll__or3_4.pex.spice
* Created: Wed Sep  2 08:48:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR3_4%C 1 3 4 6 7 12
c28 7 0 1.65414e-19 $X=0.23 $Y=1.19
r29 12 13 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r30 10 12 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r31 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r32 4 13 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r34 1 12 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_4%B 1 3 4 6 7 9 13 14
c38 7 0 1.47946e-20 $X=0.83 $Y=1.2
c39 1 0 1.65414e-19 $X=0.965 $Y=1.41
r40 13 14 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.712 $Y=1.53
+ $X2=0.712 $Y2=1.87
r41 12 13 10.0532 $w=2.33e-07 $l=2.05e-07 $layer=LI1_cond $X=0.712 $Y=1.325
+ $X2=0.712 $Y2=1.53
r42 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r43 7 12 6.82498 $w=2.5e-07 $l=1.74284e-07 $layer=LI1_cond $X=0.83 $Y=1.2
+ $X2=0.712 $Y2=1.325
r44 7 9 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=0.83 $Y=1.2 $X2=0.94
+ $Y2=1.2
r45 4 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.965 $Y2=1.16
r46 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.56
r47 1 10 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.16
r48 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_4%A 1 3 4 6 7 16
r36 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.16 $X2=1.49 $Y2=1.16
r37 7 16 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=1.2 $X2=1.615
+ $Y2=1.2
r38 7 11 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=1.61 $Y=1.2 $X2=1.49
+ $Y2=1.2
r39 4 10 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.505 $Y2=1.16
r40 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r41 1 10 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.505 $Y2=1.16
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_4%A_27_47# 1 2 3 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 36 38 40 42 43 44 48 51 52 54 55 57 59 62 67 69 79
r158 79 80 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=3.845 $Y=1.202
+ $X2=3.87 $Y2=1.202
r159 76 77 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=3.375 $Y=1.202
+ $X2=3.4 $Y2=1.202
r160 75 76 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=2.93 $Y=1.202
+ $X2=3.375 $Y2=1.202
r161 74 75 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.905 $Y=1.202
+ $X2=2.93 $Y2=1.202
r162 73 74 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=2.46 $Y=1.202
+ $X2=2.905 $Y2=1.202
r163 72 73 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.435 $Y=1.202
+ $X2=2.46 $Y2=1.202
r164 70 72 29.0521 $w=3.65e-07 $l=2.2e-07 $layer=POLY_cond $X=2.215 $Y=1.202
+ $X2=2.435 $Y2=1.202
r165 69 70 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.215
+ $Y=1.16 $X2=2.215 $Y2=1.16
r166 63 79 15.8466 $w=3.65e-07 $l=1.2e-07 $layer=POLY_cond $X=3.725 $Y=1.202
+ $X2=3.845 $Y2=1.202
r167 63 77 42.9178 $w=3.65e-07 $l=3.25e-07 $layer=POLY_cond $X=3.725 $Y=1.202
+ $X2=3.4 $Y2=1.202
r168 62 63 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.725
+ $Y=1.16 $X2=3.725 $Y2=1.16
r169 60 69 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.24 $Y=1.16
+ $X2=2.13 $Y2=1.16
r170 60 62 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=2.24 $Y=1.16
+ $X2=3.725 $Y2=1.16
r171 58 69 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=1.245
+ $X2=2.13 $Y2=1.16
r172 58 59 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=2.13 $Y=1.245
+ $X2=2.13 $Y2=1.495
r173 57 69 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=1.075
+ $X2=2.13 $Y2=1.16
r174 56 57 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=2.13 $Y=0.905
+ $X2=2.13 $Y2=1.075
r175 54 59 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.02 $Y=1.58
+ $X2=2.13 $Y2=1.495
r176 54 55 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.02 $Y=1.58
+ $X2=1.365 $Y2=1.58
r177 53 67 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0.815
+ $X2=1.175 $Y2=0.815
r178 52 56 6.90553 $w=1.8e-07 $l=1.48324e-07 $layer=LI1_cond $X=2.02 $Y=0.815
+ $X2=2.13 $Y2=0.905
r179 52 53 40.3586 $w=1.78e-07 $l=6.55e-07 $layer=LI1_cond $X=2.02 $Y=0.815
+ $X2=1.365 $Y2=0.815
r180 50 55 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=1.232 $Y=1.665
+ $X2=1.365 $Y2=1.58
r181 50 51 27.3977 $w=2.63e-07 $l=6.3e-07 $layer=LI1_cond $X=1.232 $Y=1.665
+ $X2=1.232 $Y2=2.295
r182 46 67 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.175 $Y=0.725
+ $X2=1.175 $Y2=0.815
r183 46 48 9.85642 $w=3.78e-07 $l=3.25e-07 $layer=LI1_cond $X=1.175 $Y=0.725
+ $X2=1.175 $Y2=0.4
r184 45 66 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.255 $Y2=2.38
r185 44 51 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=1.1 $Y=2.38
+ $X2=1.232 $Y2=2.295
r186 44 45 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.1 $Y=2.38
+ $X2=0.425 $Y2=2.38
r187 42 67 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0.815
+ $X2=1.175 $Y2=0.815
r188 42 43 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.815
+ $X2=0.425 $Y2=0.815
r189 38 66 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=2.295
+ $X2=0.255 $Y2=2.38
r190 38 40 21.5236 $w=3.38e-07 $l=6.35e-07 $layer=LI1_cond $X=0.255 $Y=2.295
+ $X2=0.255 $Y2=1.66
r191 34 43 7.6914 $w=1.8e-07 $l=2.10238e-07 $layer=LI1_cond $X=0.255 $Y=0.725
+ $X2=0.425 $Y2=0.815
r192 34 36 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=0.255 $Y=0.725
+ $X2=0.255 $Y2=0.4
r193 31 80 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.87 $Y=0.995
+ $X2=3.87 $Y2=1.202
r194 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.87 $Y=0.995
+ $X2=3.87 $Y2=0.56
r195 28 79 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.845 $Y=1.41
+ $X2=3.845 $Y2=1.202
r196 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.845 $Y=1.41
+ $X2=3.845 $Y2=1.985
r197 25 77 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.4 $Y=0.995
+ $X2=3.4 $Y2=1.202
r198 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.4 $Y=0.995
+ $X2=3.4 $Y2=0.56
r199 22 76 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.375 $Y=1.41
+ $X2=3.375 $Y2=1.202
r200 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.375 $Y=1.41
+ $X2=3.375 $Y2=1.985
r201 19 75 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=1.202
r202 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=0.56
r203 16 74 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.905 $Y=1.41
+ $X2=2.905 $Y2=1.202
r204 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.905 $Y=1.41
+ $X2=2.905 $Y2=1.985
r205 13 73 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.46 $Y=0.995
+ $X2=2.46 $Y2=1.202
r206 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.46 $Y=0.995
+ $X2=2.46 $Y2=0.56
r207 10 72 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.435 $Y=1.41
+ $X2=2.435 $Y2=1.202
r208 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.435 $Y=1.41
+ $X2=2.435 $Y2=1.985
r209 3 66 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r210 3 40 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r211 2 48 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.4
r212 1 36 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_4%VPWR 1 2 3 12 16 20 23 24 26 27 28 30 43 44
+ 47
r55 48 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 47 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r57 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r59 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r60 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r61 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r62 38 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r64 35 47 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=1.935 $Y2=2.72
r65 35 37 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=2.99 $Y2=2.72
r66 30 47 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=1.935 $Y2=2.72
r67 30 32 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 28 50 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r69 28 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 26 40 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.955 $Y=2.72
+ $X2=3.91 $Y2=2.72
r71 26 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.955 $Y=2.72
+ $X2=4.08 $Y2=2.72
r72 25 43 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=2.72
+ $X2=4.37 $Y2=2.72
r73 25 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.205 $Y=2.72
+ $X2=4.08 $Y2=2.72
r74 23 37 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.015 $Y=2.72
+ $X2=2.99 $Y2=2.72
r75 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.015 $Y=2.72
+ $X2=3.14 $Y2=2.72
r76 22 40 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=3.91 $Y2=2.72
r77 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=3.14 $Y2=2.72
r78 18 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=2.635
+ $X2=4.08 $Y2=2.72
r79 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.08 $Y=2.635
+ $X2=4.08 $Y2=1.96
r80 14 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=2.635
+ $X2=3.14 $Y2=2.72
r81 14 16 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.14 $Y=2.635
+ $X2=3.14 $Y2=1.96
r82 10 47 2.86223 $w=7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.935 $Y=2.635
+ $X2=1.935 $Y2=2.72
r83 10 12 10.8501 $w=6.98e-07 $l=6.35e-07 $layer=LI1_cond $X=1.935 $Y=2.635
+ $X2=1.935 $Y2=2
r84 3 20 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.935
+ $Y=1.485 $X2=4.08 $Y2=1.96
r85 2 16 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.995
+ $Y=1.485 $X2=3.14 $Y2=1.96
r86 1 12 150 $w=1.7e-07 $l=8.96242e-07 $layer=licon1_PDIFF $count=4 $X=1.525
+ $Y=1.485 $X2=2.2 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41
+ 42 44 47
r76 44 47 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.285 $Y=0.82
+ $X2=4.285 $Y2=0.905
r77 44 47 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=4.285 $Y=0.92
+ $X2=4.285 $Y2=0.905
r78 43 44 17.7951 $w=3.38e-07 $l=5.25e-07 $layer=LI1_cond $X=4.285 $Y=1.445
+ $X2=4.285 $Y2=0.92
r79 40 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.775 $Y=0.82
+ $X2=3.585 $Y2=0.82
r80 39 44 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.115 $Y=0.82
+ $X2=4.285 $Y2=0.82
r81 39 40 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.115 $Y=0.82
+ $X2=3.775 $Y2=0.82
r82 38 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.735 $Y=1.53
+ $X2=3.61 $Y2=1.53
r83 37 43 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.115 $Y=1.53
+ $X2=4.285 $Y2=1.445
r84 37 38 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.115 $Y=1.53
+ $X2=3.735 $Y2=1.53
r85 33 35 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=3.61 $Y=1.62
+ $X2=3.61 $Y2=2.3
r86 31 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=1.615
+ $X2=3.61 $Y2=1.53
r87 31 33 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.61 $Y=1.615
+ $X2=3.61 $Y2=1.62
r88 27 41 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=0.735
+ $X2=3.585 $Y2=0.82
r89 27 29 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=3.585 $Y=0.735
+ $X2=3.585 $Y2=0.39
r90 25 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.395 $Y=0.82
+ $X2=3.585 $Y2=0.82
r91 25 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.395 $Y=0.82
+ $X2=2.835 $Y2=0.82
r92 23 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.485 $Y=1.53
+ $X2=3.61 $Y2=1.53
r93 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.485 $Y=1.53
+ $X2=2.795 $Y2=1.53
r94 19 21 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.67 $Y=1.62
+ $X2=2.67 $Y2=2.3
r95 17 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.67 $Y=1.615
+ $X2=2.795 $Y2=1.53
r96 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.67 $Y=1.615
+ $X2=2.67 $Y2=1.62
r97 13 26 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.645 $Y=0.735
+ $X2=2.835 $Y2=0.82
r98 13 15 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=2.645 $Y=0.735
+ $X2=2.645 $Y2=0.39
r99 4 35 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.465
+ $Y=1.485 $X2=3.61 $Y2=2.3
r100 4 33 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.465
+ $Y=1.485 $X2=3.61 $Y2=1.62
r101 3 21 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.485 $X2=2.67 $Y2=2.3
r102 3 19 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.485 $X2=2.67 $Y2=1.62
r103 2 29 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.475
+ $Y=0.235 $X2=3.61 $Y2=0.39
r104 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.535
+ $Y=0.235 $X2=2.67 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_4%VGND 1 2 3 4 17 23 27 30 31 33 34 35 45 46
+ 49 54 60 62
r73 59 60 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0.235
+ $X2=2.285 $Y2=0.235
r74 56 59 2.42953 $w=6.38e-07 $l=1.3e-07 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.2 $Y2=0.235
r75 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r76 53 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r77 52 56 8.59681 $w=6.38e-07 $l=4.6e-07 $layer=LI1_cond $X=1.61 $Y=0.235
+ $X2=2.07 $Y2=0.235
r78 52 54 7.80044 $w=6.38e-07 $l=2.5e-08 $layer=LI1_cond $X=1.61 $Y=0.235
+ $X2=1.585 $Y2=0.235
r79 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r80 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r81 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r82 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r83 43 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r84 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r85 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r86 40 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r87 39 60 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.285
+ $Y2=0
r88 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r89 35 50 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r90 35 62 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r91 33 42 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.91
+ $Y2=0
r92 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=0 $X2=4.08
+ $Y2=0
r93 32 45 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=4.37
+ $Y2=0
r94 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=0 $X2=4.08
+ $Y2=0
r95 30 39 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=0 $X2=2.99
+ $Y2=0
r96 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0 $X2=3.14
+ $Y2=0
r97 29 42 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.91
+ $Y2=0
r98 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.14
+ $Y2=0
r99 25 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=0.085
+ $X2=4.08 $Y2=0
r100 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.08 $Y=0.085
+ $X2=4.08 $Y2=0.39
r101 21 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r102 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.39
r103 20 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r104 20 54 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.815 $Y=0
+ $X2=1.585 $Y2=0
r105 15 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r106 15 17 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.39
r107 4 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.945
+ $Y=0.235 $X2=4.08 $Y2=0.39
r108 3 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.005
+ $Y=0.235 $X2=3.14 $Y2=0.39
r109 2 59 91 $w=1.7e-07 $l=7.88701e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.235 $X2=2.2 $Y2=0.39
r110 1 17 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

