# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a221oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.145000 1.075000 8.755000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.585000 1.075000  6.965000 1.445000 ;
        RECT 6.585000 1.445000  9.135000 1.615000 ;
        RECT 8.965000 1.075000 10.400000 1.275000 ;
        RECT 8.965000 1.275000  9.135000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.335000 0.995000 5.885000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 0.995000 4.165000 1.325000 ;
        RECT 3.945000 1.325000 4.165000 1.445000 ;
        RECT 3.945000 1.445000 6.410000 1.615000 ;
        RECT 6.065000 1.075000 6.410000 1.445000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.435000 1.275000 ;
    END
  END C1
  PIN VGND
    ANTENNADIFFAREA  1.485250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.160000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.893000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 1.855000 0.905000 ;
        RECT 0.625000 1.445000 1.855000 1.615000 ;
        RECT 0.625000 1.615000 0.875000 2.125000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 1.565000 1.615000 1.815000 2.125000 ;
        RECT 1.655000 0.905000 1.855000 1.095000 ;
        RECT 1.655000 1.095000 3.595000 1.275000 ;
        RECT 1.655000 1.275000 1.855000 1.445000 ;
        RECT 3.375000 0.645000 6.280000 0.735000 ;
        RECT 3.375000 0.735000 8.585000 0.820000 ;
        RECT 3.375000 0.820000 3.595000 1.095000 ;
        RECT 6.110000 0.820000 7.130000 0.905000 ;
        RECT 6.960000 0.645000 8.585000 0.735000 ;
    END
  END Y
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.770000 2.910000 ;
    END
  END VPB
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.090000  1.445000  0.405000 2.295000 ;
      RECT  0.090000  2.295000  2.325000 2.465000 ;
      RECT  0.115000  0.085000  0.365000 0.895000 ;
      RECT  1.095000  1.785000  1.345000 2.295000 ;
      RECT  1.135000  0.085000  1.305000 0.555000 ;
      RECT  2.075000  0.085000  2.245000 0.645000 ;
      RECT  2.075000  0.645000  3.205000 0.925000 ;
      RECT  2.075000  1.445000  3.330000 1.615000 ;
      RECT  2.075000  1.615000  2.325000 2.295000 ;
      RECT  2.435000  0.255000  6.185000 0.425000 ;
      RECT  2.435000  0.425000  2.860000 0.475000 ;
      RECT  2.565000  1.795000  2.815000 2.215000 ;
      RECT  2.565000  2.215000  6.655000 2.465000 ;
      RECT  3.035000  0.595000  3.205000 0.645000 ;
      RECT  3.035000  1.615000  3.330000 1.835000 ;
      RECT  3.035000  1.835000  6.185000 2.045000 ;
      RECT  3.335000  0.425000  6.185000 0.475000 ;
      RECT  6.405000  1.785000  9.525000 2.045000 ;
      RECT  6.405000  2.045000  6.655000 2.215000 ;
      RECT  6.455000  0.085000  6.625000 0.555000 ;
      RECT  6.795000  0.255000  9.055000 0.475000 ;
      RECT  6.825000  2.215000  9.085000 2.635000 ;
      RECT  8.805000  0.475000  9.055000 0.725000 ;
      RECT  8.805000  0.725000  9.995000 0.905000 ;
      RECT  9.275000  0.085000  9.445000 0.555000 ;
      RECT  9.275000  2.045000  9.445000 2.465000 ;
      RECT  9.355000  1.445000 10.425000 1.615000 ;
      RECT  9.355000  1.615000  9.525000 1.785000 ;
      RECT  9.615000  0.255000  9.995000 0.725000 ;
      RECT  9.745000  1.795000  9.915000 2.635000 ;
      RECT 10.165000  0.085000 10.335000 0.905000 ;
      RECT 10.175000  1.615000 10.425000 2.465000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a221oi_4
END LIBRARY
