* File: sky130_fd_sc_hdll__or3_4.spice
* Created: Wed Sep  2 08:48:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or3_4.pex.spice"
.subckt sky130_fd_sc_hdll__or3_4  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_C_M1010_g N_A_27_47#_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_47#_M1001_d N_B_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_27_47#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2925 AS=0.08775 PD=1.55 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1003_d N_A_27_47#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2925 AS=0.104 PD=1.55 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_27_47#_M1007_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1007_d N_A_27_47#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_27_47#_M1011_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.20475 AS=0.104 PD=1.93 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 A_117_297# N_C_M1005_g N_A_27_47#_M1005_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=17.7103 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90003.6 A=0.18 P=2.36 MULT=1
MM1000 A_211_297# N_B_M1000_g A_117_297# VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=17.7103 NRS=17.7103 M=1 R=5.55556 SA=90000.6
+ SB=90003.2 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g A_211_297# VPB PHIGHVT L=0.18 W=1 AD=0.41
+ AS=0.145 PD=1.82 PS=1.29 NRD=13.7703 NRS=17.7103 M=1 R=5.55556 SA=90001.1
+ SB=90002.7 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1012_d N_A_27_47#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.41 AS=0.145 PD=1.82 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_27_47#_M1004_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1004_d N_A_27_47#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A_27_47#_M1013_g N_X_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.37 AS=0.145 PD=2.74 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.3 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
c_76 VPB 0 1.47946e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__or3_4.pxi.spice"
*
.ends
*
*
