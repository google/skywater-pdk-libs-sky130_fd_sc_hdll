* File: sky130_fd_sc_hdll__o211ai_1.pxi.spice
* Created: Thu Aug 27 19:18:31 2020
* 
x_PM_SKY130_FD_SC_HDLL__O211AI_1%A1 N_A1_c_40_n N_A1_M1005_g N_A1_c_41_n
+ N_A1_M1000_g A1 PM_SKY130_FD_SC_HDLL__O211AI_1%A1
x_PM_SKY130_FD_SC_HDLL__O211AI_1%A2 N_A2_c_63_n N_A2_M1002_g N_A2_c_64_n
+ N_A2_M1001_g N_A2_c_65_n A2 PM_SKY130_FD_SC_HDLL__O211AI_1%A2
x_PM_SKY130_FD_SC_HDLL__O211AI_1%B1 N_B1_c_99_n N_B1_M1007_g N_B1_c_100_n
+ N_B1_M1003_g B1 B1 PM_SKY130_FD_SC_HDLL__O211AI_1%B1
x_PM_SKY130_FD_SC_HDLL__O211AI_1%C1 N_C1_c_129_n N_C1_M1004_g N_C1_c_130_n
+ N_C1_M1006_g C1 N_C1_c_132_n PM_SKY130_FD_SC_HDLL__O211AI_1%C1
x_PM_SKY130_FD_SC_HDLL__O211AI_1%VPWR N_VPWR_M1005_s N_VPWR_M1003_d
+ N_VPWR_c_156_n N_VPWR_c_157_n N_VPWR_c_158_n VPWR N_VPWR_c_159_n
+ N_VPWR_c_160_n N_VPWR_c_155_n N_VPWR_c_162_n
+ PM_SKY130_FD_SC_HDLL__O211AI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O211AI_1%Y N_Y_M1004_d N_Y_M1002_d N_Y_M1006_d
+ N_Y_c_203_n N_Y_c_193_n N_Y_c_197_n N_Y_c_198_n N_Y_c_195_n N_Y_c_194_n Y
+ N_Y_c_206_n PM_SKY130_FD_SC_HDLL__O211AI_1%Y
x_PM_SKY130_FD_SC_HDLL__O211AI_1%A_27_47# N_A_27_47#_M1000_s N_A_27_47#_M1001_d
+ N_A_27_47#_c_237_n N_A_27_47#_c_239_n N_A_27_47#_c_238_n N_A_27_47#_c_242_n
+ PM_SKY130_FD_SC_HDLL__O211AI_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O211AI_1%VGND N_VGND_M1000_d N_VGND_c_263_n VGND
+ N_VGND_c_264_n N_VGND_c_265_n N_VGND_c_266_n N_VGND_c_267_n
+ PM_SKY130_FD_SC_HDLL__O211AI_1%VGND
cc_1 VNB N_A1_c_40_n 0.0326818f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_2 VNB N_A1_c_41_n 0.0224994f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_3 VNB A1 0.0125518f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A2_c_63_n 0.019402f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_5 VNB N_A2_c_64_n 0.017224f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_6 VNB N_A2_c_65_n 0.00450877f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_7 VNB N_B1_c_99_n 0.0175975f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_8 VNB N_B1_c_100_n 0.0243505f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_9 VNB B1 0.0104129f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_10 VNB N_C1_c_129_n 0.0208602f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_11 VNB N_C1_c_130_n 0.0319886f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_12 VNB N_VPWR_c_155_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_Y_c_193_n 0.0246328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_194_n 0.0240081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_237_n 0.0140519f $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.16
cc_16 VNB N_A_27_47#_c_238_n 0.00921527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_263_n 0.00276073f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.56
cc_18 VNB N_VGND_c_264_n 0.0155904f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_19 VNB N_VGND_c_265_n 0.0476646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_266_n 0.162188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_267_n 0.0050671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_A1_c_40_n 0.0351367f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_23 VPB A1 0.00184586f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_24 VPB N_A2_c_63_n 0.0243996f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_25 VPB N_A2_c_65_n 7.56831e-19 $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_26 VPB A2 5.99582e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_B1_c_100_n 0.0270128f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_28 VPB B1 0.00108009f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_29 VPB N_C1_c_130_n 0.0342144f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_30 VPB N_C1_c_132_n 0.00148865f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_31 VPB N_VPWR_c_156_n 0.0109759f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_VPWR_c_157_n 0.0435899f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.16
cc_33 VPB N_VPWR_c_158_n 0.00285982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_159_n 0.0298338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_160_n 0.0238665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_155_n 0.0435986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_162_n 0.00512961f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_Y_c_195_n 0.0275968f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_Y_c_194_n 0.0214741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 N_A1_c_40_n N_A2_c_63_n 0.0962299f $X=0.5 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_41 N_A1_c_41_n N_A2_c_64_n 0.0221742f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_42 N_A1_c_40_n N_A2_c_65_n 0.00935108f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_43 A1 N_A2_c_65_n 0.0256264f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_44 N_A1_c_40_n A2 0.0257471f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_45 N_A1_c_40_n N_VPWR_c_157_n 0.00986695f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_46 A1 N_VPWR_c_157_n 0.0231627f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_47 N_A1_c_40_n N_VPWR_c_159_n 0.00672576f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_48 N_A1_c_40_n N_VPWR_c_155_n 0.012411f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_49 N_A1_c_40_n N_Y_c_197_n 4.32038e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_50 N_A1_c_40_n N_Y_c_198_n 5.35664e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_51 N_A1_c_41_n N_A_27_47#_c_239_n 0.0174439f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_52 N_A1_c_40_n N_A_27_47#_c_238_n 0.00518572f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_53 A1 N_A_27_47#_c_238_n 0.0247373f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A1_c_41_n N_A_27_47#_c_242_n 3.68761e-19 $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_55 N_A1_c_41_n N_VGND_c_263_n 0.00811875f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_56 N_A1_c_41_n N_VGND_c_264_n 0.00337001f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_57 N_A1_c_41_n N_VGND_c_266_n 0.00498987f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_58 N_A2_c_64_n N_B1_c_99_n 0.0127704f $X=1.005 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_59 N_A2_c_63_n N_B1_c_100_n 0.0352137f $X=0.91 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A2_c_65_n N_B1_c_100_n 0.00130741f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_61 A2 N_B1_c_100_n 8.39578e-19 $X=0.6 $Y=1.445 $X2=0 $Y2=0
cc_62 N_A2_c_63_n B1 0.0010105f $X=0.91 $Y=1.41 $X2=0 $Y2=0
cc_63 N_A2_c_65_n B1 0.0146841f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_64 A2 B1 0.00623952f $X=0.6 $Y=1.445 $X2=0 $Y2=0
cc_65 N_A2_c_63_n N_VPWR_c_158_n 9.22834e-19 $X=0.91 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A2_c_63_n N_VPWR_c_159_n 0.00691519f $X=0.91 $Y=1.41 $X2=0 $Y2=0
cc_67 A2 N_VPWR_c_159_n 0.00589613f $X=0.6 $Y=1.445 $X2=0 $Y2=0
cc_68 N_A2_c_63_n N_VPWR_c_155_n 0.0124552f $X=0.91 $Y=1.41 $X2=0 $Y2=0
cc_69 A2 N_VPWR_c_155_n 0.00859471f $X=0.6 $Y=1.445 $X2=0 $Y2=0
cc_70 A2 A_118_297# 0.00169349f $X=0.6 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_71 N_A2_c_63_n N_Y_c_197_n 0.00766773f $X=0.91 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A2_c_65_n N_Y_c_197_n 0.0030046f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_73 A2 N_Y_c_197_n 0.0482352f $X=0.6 $Y=1.445 $X2=0 $Y2=0
cc_74 N_A2_c_63_n N_Y_c_198_n 0.0061869f $X=0.91 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A2_c_63_n N_A_27_47#_c_239_n 0.00301656f $X=0.91 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A2_c_64_n N_A_27_47#_c_239_n 0.011183f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A2_c_65_n N_A_27_47#_c_239_n 0.0340359f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A2_c_64_n N_A_27_47#_c_242_n 0.00591749f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A2_c_65_n N_A_27_47#_c_242_n 6.6737e-19 $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A2_c_64_n N_VGND_c_263_n 0.00308386f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A2_c_64_n N_VGND_c_265_n 0.00419334f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A2_c_64_n N_VGND_c_266_n 0.00577133f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_83 N_B1_c_99_n N_C1_c_129_n 0.0275931f $X=1.445 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_84 N_B1_c_100_n N_C1_c_130_n 0.0590798f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_85 B1 N_C1_c_130_n 0.00438568f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_86 N_B1_c_100_n N_C1_c_132_n 5.98806e-19 $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_87 B1 N_C1_c_132_n 0.0468546f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_88 B1 N_VPWR_M1003_d 0.00261369f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_89 N_B1_c_100_n N_VPWR_c_158_n 0.00781145f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B1_c_100_n N_VPWR_c_159_n 0.00458874f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B1_c_100_n N_VPWR_c_155_n 0.00551952f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_92 N_B1_c_100_n N_Y_c_203_n 0.0177197f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_93 B1 N_Y_c_203_n 0.0161659f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_94 N_B1_c_100_n N_Y_c_195_n 8.72769e-19 $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B1_c_99_n N_Y_c_206_n 0.004805f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_96 B1 N_Y_c_206_n 0.00179418f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_97 N_B1_c_99_n N_A_27_47#_c_242_n 0.0128654f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_98 B1 N_A_27_47#_c_242_n 0.00230436f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B1_c_99_n N_VGND_c_265_n 0.00465454f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B1_c_99_n N_VGND_c_266_n 0.00820049f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_101 N_C1_c_130_n N_VPWR_c_158_n 0.00423652f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_102 N_C1_c_130_n N_VPWR_c_160_n 0.00513711f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_103 N_C1_c_130_n N_VPWR_c_155_n 0.00802261f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_104 N_C1_c_132_n N_Y_M1006_d 0.00291874f $X=2.105 $Y=1.16 $X2=0 $Y2=0
cc_105 N_C1_c_130_n N_Y_c_203_n 0.0145001f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_106 N_C1_c_132_n N_Y_c_203_n 0.0107344f $X=2.105 $Y=1.16 $X2=0 $Y2=0
cc_107 N_C1_c_130_n N_Y_c_195_n 0.0243597f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_108 N_C1_c_132_n N_Y_c_195_n 0.0106628f $X=2.105 $Y=1.16 $X2=0 $Y2=0
cc_109 N_C1_c_129_n N_Y_c_194_n 0.00473798f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_110 N_C1_c_130_n N_Y_c_194_n 0.0157224f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_111 N_C1_c_132_n N_Y_c_194_n 0.0469185f $X=2.105 $Y=1.16 $X2=0 $Y2=0
cc_112 N_C1_c_129_n N_Y_c_206_n 0.0313023f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_113 N_C1_c_130_n N_Y_c_206_n 0.00636655f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_114 N_C1_c_132_n N_Y_c_206_n 0.0243681f $X=2.105 $Y=1.16 $X2=0 $Y2=0
cc_115 N_C1_c_129_n N_A_27_47#_c_242_n 5.26337e-19 $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_116 N_C1_c_129_n N_VGND_c_265_n 0.00357877f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C1_c_129_n N_VGND_c_266_n 0.00673322f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_118 N_VPWR_c_155_n A_118_297# 0.00218212f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_119 N_VPWR_c_155_n N_Y_M1002_d 0.00327804f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_120 N_VPWR_c_155_n N_Y_M1006_d 0.00439666f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_121 N_VPWR_M1003_d N_Y_c_203_n 0.00818614f $X=1.56 $Y=1.485 $X2=0 $Y2=0
cc_122 N_VPWR_c_158_n N_Y_c_203_n 0.0148805f $X=1.705 $Y=2.36 $X2=0 $Y2=0
cc_123 N_VPWR_c_159_n N_Y_c_203_n 0.00291265f $X=1.54 $Y=2.72 $X2=0 $Y2=0
cc_124 N_VPWR_c_160_n N_Y_c_203_n 0.00288861f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_125 N_VPWR_c_155_n N_Y_c_203_n 0.0116345f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_126 N_VPWR_c_159_n N_Y_c_198_n 0.0186279f $X=1.54 $Y=2.72 $X2=0 $Y2=0
cc_127 N_VPWR_c_155_n N_Y_c_198_n 0.0124148f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_128 N_VPWR_c_160_n N_Y_c_195_n 0.0400427f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_129 N_VPWR_c_155_n N_Y_c_195_n 0.0229723f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_130 N_Y_c_206_n N_A_27_47#_c_242_n 0.0327308f $X=2.44 $Y=0.54 $X2=0 $Y2=0
cc_131 N_Y_c_193_n N_VGND_c_265_n 0.0165941f $X=2.557 $Y=0.825 $X2=0 $Y2=0
cc_132 N_Y_c_206_n N_VGND_c_265_n 0.0451177f $X=2.44 $Y=0.54 $X2=0 $Y2=0
cc_133 N_Y_M1004_d N_VGND_c_266_n 0.00472496f $X=2.045 $Y=0.235 $X2=0 $Y2=0
cc_134 N_Y_c_193_n N_VGND_c_266_n 0.00905026f $X=2.557 $Y=0.825 $X2=0 $Y2=0
cc_135 N_Y_c_206_n N_VGND_c_266_n 0.0267029f $X=2.44 $Y=0.54 $X2=0 $Y2=0
cc_136 N_Y_c_206_n A_304_47# 0.0115248f $X=2.44 $Y=0.54 $X2=-0.19 $Y2=-0.24
cc_137 N_A_27_47#_c_239_n N_VGND_M1000_d 0.00438654f $X=1.07 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_138 N_A_27_47#_c_239_n N_VGND_c_263_n 0.0186469f $X=1.07 $Y=0.72 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_237_n N_VGND_c_264_n 0.0208826f $X=0.26 $Y=0.485 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_239_n N_VGND_c_264_n 0.00258359f $X=1.07 $Y=0.72 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_239_n N_VGND_c_265_n 0.00273188f $X=1.07 $Y=0.72 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_242_n N_VGND_c_265_n 0.0221228f $X=1.235 $Y=0.38 $X2=0 $Y2=0
cc_143 N_A_27_47#_M1000_s N_VGND_c_266_n 0.00271217f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_M1001_d N_VGND_c_266_n 0.00231261f $X=1.08 $Y=0.235 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_c_237_n N_VGND_c_266_n 0.0116156f $X=0.26 $Y=0.485 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_239_n N_VGND_c_266_n 0.0100606f $X=1.07 $Y=0.72 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_242_n N_VGND_c_266_n 0.0139443f $X=1.235 $Y=0.38 $X2=0 $Y2=0
cc_148 N_VGND_c_266_n A_304_47# 0.0101281f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
