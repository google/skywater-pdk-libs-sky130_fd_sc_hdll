* File: sky130_fd_sc_hdll__or2b_4.spice
* Created: Wed Sep  2 08:48:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or2b_4.pex.spice"
.subckt sky130_fd_sc_hdll__or2b_4  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_B_N_M1000_g N_A_27_53#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.17116 AS=0.1302 PD=1.13832 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_229_297#_M1004_d N_A_27_53#_M1004_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.26489 PD=0.92 PS=1.76168 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.9 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_229_297#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.08775 PD=1.04 PS=0.92 NRD=21.228 NRS=0 M=1 R=4.33333
+ SA=75001.3 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1008_d N_A_229_297#_M1008_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12675 PD=0.97 PS=1.04 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1008_d N_A_229_297#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.3
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1010_d N_A_229_297#_M1010_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1013 N_X_M1010_d N_A_229_297#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.2145 PD=1.02 PS=1.96 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.3
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_53#_M1001_d N_B_N_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1218 AS=0.1134 PD=1.42 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1005 A_319_297# N_A_27_53#_M1005_g N_A_229_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.115 AS=0.27 PD=1.23 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_319_297# VPB PHIGHVT L=0.18 W=1 AD=0.18
+ AS=0.115 PD=1.36 PS=1.23 NRD=13.7703 NRS=11.8003 M=1 R=5.55556 SA=90000.6
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1007_d N_A_229_297#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.18 AS=0.145 PD=1.36 PS=1.29 NRD=1.9503 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_229_297#_M1006_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1006_d N_A_229_297#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_229_297#_M1012_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.305 AS=0.145 PD=2.61 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX15_noxref noxref_11 A A PROBETYPE=1
*
.include "sky130_fd_sc_hdll__or2b_4.pxi.spice"
*
.ends
*
*
