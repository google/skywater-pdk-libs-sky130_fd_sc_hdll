* File: sky130_fd_sc_hdll__or4bb_4.spice
* Created: Wed Sep  2 08:50:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or4bb_4.pex.spice"
.subckt sky130_fd_sc_hdll__or4bb_4  VNB VPB C_N D_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C_N_M1008_g N_A_27_410#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07245 AS=0.1302 PD=0.765 PS=1.46 NRD=5.712 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_224_297#_M1004_d N_D_N_M1004_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.07245 PD=1.36 PS=0.765 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_335_297#_M1011_d N_A_224_297#_M1011_g N_VGND_M1011_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.13 AS=0.2015 PD=1.05 PS=1.92 NRD=13.836 NRS=8.304 M=1
+ R=4.33333 SA=75000.2 SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_27_410#_M1012_g N_A_335_297#_M1011_d VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.13 PD=0.97 PS=1.05 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.8 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1005 N_A_335_297#_M1005_d N_B_M1005_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.3
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_335_297#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1365 AS=0.08775 PD=1.07 PS=0.92 NRD=24.912 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_335_297#_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.1365 PD=0.97 PS=1.07 NRD=8.304 NRS=0.912 M=1 R=4.33333
+ SA=75002.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1013 N_X_M1006_d N_A_335_297#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1015 N_X_M1015_d N_A_335_297#_M1015_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1019 N_X_M1015_d N_A_335_297#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_VPWR_M1014_d N_C_N_M1014_g N_A_27_410#_M1014_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.126812 AS=0.1134 PD=1.34 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1017 N_A_224_297#_M1017_d N_D_N_M1017_g N_VPWR_M1014_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.126812 PD=1.38 PS=1.34 NRD=2.3443 NRS=115.816 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1001 A_425_297# N_A_224_297#_M1001_g N_A_335_297#_M1001_s VPB PHIGHVT L=0.18
+ W=1 AD=0.175 AS=0.27 PD=1.35 PS=2.54 NRD=23.6203 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.6 A=0.18 P=2.36 MULT=1
MM1010 A_531_297# N_A_27_410#_M1010_g A_425_297# VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.175 PD=1.29 PS=1.35 NRD=17.7103 NRS=23.6203 M=1 R=5.55556 SA=90000.7
+ SB=90003.1 A=0.18 P=2.36 MULT=1
MM1009 A_625_297# N_B_M1009_g A_531_297# VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=17.7103 NRS=17.7103 M=1 R=5.55556 SA=90001.2
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g A_625_297# VPB PHIGHVT L=0.18 W=1 AD=0.195
+ AS=0.145 PD=1.39 PS=1.29 NRD=9.8303 NRS=17.7103 M=1 R=5.55556 SA=90001.6
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1000 N_X_M1000_d N_A_335_297#_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.195 PD=1.29 PS=1.39 NRD=0.9653 NRS=11.8003 M=1 R=5.55556
+ SA=90002.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1007 N_X_M1000_d N_A_335_297#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1016 N_X_M1016_d N_A_335_297#_M1016_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1018 N_X_M1016_d N_A_335_297#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.335 P=15.97
*
.include "sky130_fd_sc_hdll__or4bb_4.pxi.spice"
*
.ends
*
*
