* File: sky130_fd_sc_hdll__nand2_12.pxi.spice
* Created: Wed Sep  2 08:36:22 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2_12%B N_B_c_132_n N_B_M1003_g N_B_c_146_n
+ N_B_M1000_g N_B_c_147_n N_B_M1001_g N_B_c_133_n N_B_M1011_g N_B_c_134_n
+ N_B_M1013_g N_B_c_148_n N_B_M1004_g N_B_c_149_n N_B_M1005_g N_B_c_135_n
+ N_B_M1016_g N_B_c_136_n N_B_M1021_g N_B_c_150_n N_B_M1012_g N_B_c_151_n
+ N_B_M1015_g N_B_c_137_n N_B_M1026_g N_B_c_138_n N_B_M1031_g N_B_c_152_n
+ N_B_M1022_g N_B_c_153_n N_B_M1025_g N_B_c_139_n N_B_M1036_g N_B_c_140_n
+ N_B_M1040_g N_B_c_154_n N_B_M1029_g N_B_c_155_n N_B_M1033_g N_B_c_141_n
+ N_B_M1042_g N_B_c_142_n N_B_M1043_g N_B_c_156_n N_B_M1038_g N_B_c_157_n
+ N_B_M1041_g N_B_c_143_n N_B_M1044_g B N_B_c_144_n N_B_c_145_n
+ PM_SKY130_FD_SC_HDLL__NAND2_12%B
x_PM_SKY130_FD_SC_HDLL__NAND2_12%A N_A_c_384_n N_A_M1007_g N_A_c_397_n
+ N_A_M1002_g N_A_c_385_n N_A_M1008_g N_A_c_398_n N_A_M1006_g N_A_c_386_n
+ N_A_M1009_g N_A_c_399_n N_A_M1010_g N_A_c_400_n N_A_M1017_g N_A_c_387_n
+ N_A_M1014_g N_A_c_388_n N_A_M1018_g N_A_c_401_n N_A_M1020_g N_A_c_402_n
+ N_A_M1023_g N_A_c_389_n N_A_M1019_g N_A_c_390_n N_A_M1024_g N_A_c_403_n
+ N_A_M1030_g N_A_c_391_n N_A_M1027_g N_A_c_404_n N_A_M1035_g N_A_c_392_n
+ N_A_M1028_g N_A_c_405_n N_A_M1037_g N_A_c_406_n N_A_M1039_g N_A_c_393_n
+ N_A_M1032_g N_A_c_394_n N_A_M1034_g N_A_c_407_n N_A_M1046_g N_A_c_408_n
+ N_A_M1047_g N_A_c_395_n N_A_M1045_g A N_A_c_465_p N_A_c_396_n
+ PM_SKY130_FD_SC_HDLL__NAND2_12%A
x_PM_SKY130_FD_SC_HDLL__NAND2_12%VPWR N_VPWR_M1000_d N_VPWR_M1001_d
+ N_VPWR_M1005_d N_VPWR_M1015_d N_VPWR_M1025_d N_VPWR_M1033_d N_VPWR_M1041_d
+ N_VPWR_M1006_d N_VPWR_M1017_d N_VPWR_M1023_d N_VPWR_M1035_d N_VPWR_M1039_d
+ N_VPWR_M1047_d N_VPWR_c_580_n N_VPWR_c_581_n N_VPWR_c_582_n N_VPWR_c_583_n
+ N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_588_n
+ N_VPWR_c_589_n N_VPWR_c_590_n N_VPWR_c_591_n N_VPWR_c_592_n N_VPWR_c_593_n
+ N_VPWR_c_594_n N_VPWR_c_595_n N_VPWR_c_596_n N_VPWR_c_597_n N_VPWR_c_598_n
+ N_VPWR_c_599_n N_VPWR_c_600_n N_VPWR_c_601_n N_VPWR_c_602_n N_VPWR_c_603_n
+ N_VPWR_c_604_n N_VPWR_c_605_n N_VPWR_c_606_n N_VPWR_c_607_n N_VPWR_c_608_n
+ N_VPWR_c_609_n N_VPWR_c_610_n N_VPWR_c_611_n N_VPWR_c_612_n VPWR
+ N_VPWR_c_613_n N_VPWR_c_579_n N_VPWR_c_615_n N_VPWR_c_616_n N_VPWR_c_617_n
+ N_VPWR_c_618_n N_VPWR_c_619_n PM_SKY130_FD_SC_HDLL__NAND2_12%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2_12%Y N_Y_M1007_d N_Y_M1009_d N_Y_M1018_d
+ N_Y_M1024_d N_Y_M1028_d N_Y_M1034_d N_Y_M1000_s N_Y_M1004_s N_Y_M1012_s
+ N_Y_M1022_s N_Y_M1029_s N_Y_M1038_s N_Y_M1002_s N_Y_M1010_s N_Y_M1020_s
+ N_Y_M1030_s N_Y_M1037_s N_Y_M1046_s N_Y_c_760_n N_Y_c_764_n N_Y_c_767_n
+ N_Y_c_771_n N_Y_c_775_n N_Y_c_779_n N_Y_c_783_n N_Y_c_787_n N_Y_c_791_n
+ N_Y_c_795_n N_Y_c_799_n N_Y_c_803_n N_Y_c_806_n N_Y_c_834_n N_Y_c_808_n
+ N_Y_c_838_n N_Y_c_850_n N_Y_c_854_n N_Y_c_858_n N_Y_c_862_n N_Y_c_866_n
+ N_Y_c_870_n N_Y_c_874_n N_Y_c_878_n N_Y_c_882_n N_Y_c_886_n N_Y_c_997_p
+ N_Y_c_757_n N_Y_c_809_n N_Y_c_813_n N_Y_c_817_n N_Y_c_821_n N_Y_c_825_n
+ N_Y_c_892_n N_Y_c_895_n N_Y_c_899_n N_Y_c_903_n N_Y_c_907_n N_Y_c_911_n
+ N_Y_c_754_n N_Y_c_755_n Y N_Y_c_756_n Y PM_SKY130_FD_SC_HDLL__NAND2_12%Y
x_PM_SKY130_FD_SC_HDLL__NAND2_12%A_27_47# N_A_27_47#_M1003_d N_A_27_47#_M1011_d
+ N_A_27_47#_M1016_d N_A_27_47#_M1026_d N_A_27_47#_M1036_d N_A_27_47#_M1042_d
+ N_A_27_47#_M1044_d N_A_27_47#_M1008_s N_A_27_47#_M1014_s N_A_27_47#_M1019_s
+ N_A_27_47#_M1027_s N_A_27_47#_M1032_s N_A_27_47#_M1045_s N_A_27_47#_c_1006_n
+ N_A_27_47#_c_1018_n N_A_27_47#_c_1007_n N_A_27_47#_c_1025_n
+ N_A_27_47#_c_1029_n N_A_27_47#_c_1033_n N_A_27_47#_c_1037_n
+ N_A_27_47#_c_1041_n N_A_27_47#_c_1045_n N_A_27_47#_c_1049_n
+ N_A_27_47#_c_1053_n N_A_27_47#_c_1057_n N_A_27_47#_c_1061_n
+ N_A_27_47#_c_1065_n N_A_27_47#_c_1008_n N_A_27_47#_c_1089_n
+ N_A_27_47#_c_1009_n N_A_27_47#_c_1010_n N_A_27_47#_c_1011_n
+ N_A_27_47#_c_1012_n N_A_27_47#_c_1013_n N_A_27_47#_c_1014_n
+ N_A_27_47#_c_1015_n PM_SKY130_FD_SC_HDLL__NAND2_12%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND2_12%VGND N_VGND_M1003_s N_VGND_M1013_s
+ N_VGND_M1021_s N_VGND_M1031_s N_VGND_M1040_s N_VGND_M1043_s N_VGND_c_1182_n
+ N_VGND_c_1183_n N_VGND_c_1184_n N_VGND_c_1185_n N_VGND_c_1186_n
+ N_VGND_c_1187_n N_VGND_c_1188_n N_VGND_c_1189_n N_VGND_c_1190_n
+ N_VGND_c_1191_n N_VGND_c_1192_n N_VGND_c_1193_n VGND N_VGND_c_1194_n
+ N_VGND_c_1195_n N_VGND_c_1196_n N_VGND_c_1197_n N_VGND_c_1198_n
+ N_VGND_c_1199_n N_VGND_c_1200_n N_VGND_c_1201_n
+ PM_SKY130_FD_SC_HDLL__NAND2_12%VGND
cc_1 VNB N_B_c_132_n 0.0228251f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B_c_133_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_B_c_134_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_4 VNB N_B_c_135_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_B_c_136_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.995
cc_6 VNB N_B_c_137_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.995
cc_7 VNB N_B_c_138_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.995
cc_8 VNB N_B_c_139_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.995
cc_9 VNB N_B_c_140_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=0.995
cc_10 VNB N_B_c_141_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=4.75 $Y2=0.995
cc_11 VNB N_B_c_142_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.995
cc_12 VNB N_B_c_143_n 0.0171127f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=0.995
cc_13 VNB N_B_c_144_n 0.0120453f $X=-0.19 $Y=-0.24 $X2=5.6 $Y2=1.16
cc_14 VNB N_B_c_145_n 0.232215f $X=-0.19 $Y=-0.24 $X2=5.665 $Y2=1.202
cc_15 VNB N_A_c_384_n 0.0162568f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_16 VNB N_A_c_385_n 0.0168735f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_17 VNB N_A_c_386_n 0.0173555f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_18 VNB N_A_c_387_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_19 VNB N_A_c_388_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.995
cc_20 VNB N_A_c_389_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.995
cc_21 VNB N_A_c_390_n 0.0164369f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.995
cc_22 VNB N_A_c_391_n 0.0169186f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_23 VNB N_A_c_392_n 0.0173608f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=0.995
cc_24 VNB N_A_c_393_n 0.0168753f $X=-0.19 $Y=-0.24 $X2=4.75 $Y2=0.995
cc_25 VNB N_A_c_394_n 0.0168204f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.995
cc_26 VNB N_A_c_395_n 0.0228463f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=0.995
cc_27 VNB N_A_c_396_n 0.232169f $X=-0.19 $Y=-0.24 $X2=5.665 $Y2=1.202
cc_28 VNB N_VPWR_c_579_n 0.497461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_754_n 0.00209731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_755_n 0.0101903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_756_n 0.00106016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_1006_n 0.0182048f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.985
cc_33 VNB N_A_27_47#_c_1007_n 0.0120628f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.985
cc_34 VNB N_A_27_47#_c_1008_n 0.00257277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.202
cc_35 VNB N_A_27_47#_c_1009_n 0.00914706f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=1.202
cc_36 VNB N_A_27_47#_c_1010_n 0.0204013f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.202
cc_37 VNB N_A_27_47#_c_1011_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=1.202
cc_38 VNB N_A_27_47#_c_1012_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=4.255 $Y2=1.202
cc_39 VNB N_A_27_47#_c_1013_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=4.725 $Y2=1.202
cc_40 VNB N_A_27_47#_c_1014_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=4.75 $Y2=1.202
cc_41 VNB N_A_27_47#_c_1015_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=1.202
cc_42 VNB N_VGND_c_1182_n 0.00466649f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_43 VNB N_VGND_c_1183_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_44 VNB N_VGND_c_1184_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.56
cc_45 VNB N_VGND_c_1185_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.985
cc_46 VNB N_VGND_c_1186_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.985
cc_47 VNB N_VGND_c_1187_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.56
cc_48 VNB N_VGND_c_1188_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.56
cc_49 VNB N_VGND_c_1189_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.985
cc_50 VNB N_VGND_c_1190_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.985
cc_51 VNB N_VGND_c_1191_n 0.00466098f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=0.995
cc_52 VNB N_VGND_c_1192_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=4.255 $Y2=1.41
cc_53 VNB N_VGND_c_1193_n 0.00515836f $X=-0.19 $Y=-0.24 $X2=4.255 $Y2=1.985
cc_54 VNB N_VGND_c_1194_n 0.0171658f $X=-0.19 $Y=-0.24 $X2=4.725 $Y2=1.985
cc_55 VNB N_VGND_c_1195_n 0.147159f $X=-0.19 $Y=-0.24 $X2=5.665 $Y2=1.985
cc_56 VNB N_VGND_c_1196_n 0.549424f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=0.995
cc_57 VNB N_VGND_c_1197_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.105
cc_58 VNB N_VGND_c_1198_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_59 VNB N_VGND_c_1199_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_60 VNB N_VGND_c_1200_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.202
cc_61 VNB N_VGND_c_1201_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_62 VPB N_B_c_146_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_63 VPB N_B_c_147_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_64 VPB N_B_c_148_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_65 VPB N_B_c_149_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_66 VPB N_B_c_150_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_67 VPB N_B_c_151_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_68 VPB N_B_c_152_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_69 VPB N_B_c_153_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_70 VPB N_B_c_154_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.41
cc_71 VPB N_B_c_155_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.725 $Y2=1.41
cc_72 VPB N_B_c_156_n 0.0162635f $X=-0.19 $Y=1.305 $X2=5.195 $Y2=1.41
cc_73 VPB N_B_c_157_n 0.0164324f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.41
cc_74 VPB N_B_c_144_n 9.19116e-19 $X=-0.19 $Y=1.305 $X2=5.6 $Y2=1.16
cc_75 VPB N_B_c_145_n 0.153595f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.202
cc_76 VPB N_A_c_397_n 0.0160834f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_77 VPB N_A_c_398_n 0.0162386f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_78 VPB N_A_c_399_n 0.016261f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_79 VPB N_A_c_400_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_80 VPB N_A_c_401_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_81 VPB N_A_c_402_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_82 VPB N_A_c_403_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_83 VPB N_A_c_404_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.995
cc_84 VPB N_A_c_405_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.41
cc_85 VPB N_A_c_406_n 0.0162606f $X=-0.19 $Y=1.305 $X2=4.725 $Y2=1.41
cc_86 VPB N_A_c_407_n 0.016238f $X=-0.19 $Y=1.305 $X2=5.195 $Y2=1.41
cc_87 VPB N_A_c_408_n 0.0207627f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.41
cc_88 VPB N_A_c_396_n 0.153211f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.202
cc_89 VPB N_VPWR_c_580_n 0.0113525f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_90 VPB N_VPWR_c_581_n 0.0410822f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.985
cc_91 VPB N_VPWR_c_582_n 0.0041373f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.56
cc_92 VPB N_VPWR_c_583_n 0.017949f $X=-0.19 $Y=1.305 $X2=4.23 $Y2=0.56
cc_93 VPB N_VPWR_c_584_n 0.0041373f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.985
cc_94 VPB N_VPWR_c_585_n 0.017949f $X=-0.19 $Y=1.305 $X2=4.725 $Y2=1.985
cc_95 VPB N_VPWR_c_586_n 0.0041373f $X=-0.19 $Y=1.305 $X2=4.75 $Y2=0.56
cc_96 VPB N_VPWR_c_587_n 0.017949f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=0.56
cc_97 VPB N_VPWR_c_588_n 0.0041373f $X=-0.19 $Y=1.305 $X2=5.195 $Y2=1.985
cc_98 VPB N_VPWR_c_589_n 0.017949f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.985
cc_99 VPB N_VPWR_c_590_n 0.0041373f $X=-0.19 $Y=1.305 $X2=5.69 $Y2=0.56
cc_100 VPB N_VPWR_c_591_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_101 VPB N_VPWR_c_592_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_102 VPB N_VPWR_c_593_n 0.0041373f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_103 VPB N_VPWR_c_594_n 0.0041373f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.202
cc_104 VPB N_VPWR_c_595_n 0.0041373f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.202
cc_105 VPB N_VPWR_c_596_n 0.0041373f $X=-0.19 $Y=1.305 $X2=4.725 $Y2=1.202
cc_106 VPB N_VPWR_c_597_n 0.0410822f $X=-0.19 $Y=1.305 $X2=5.6 $Y2=1.202
cc_107 VPB N_VPWR_c_598_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_108 VPB N_VPWR_c_599_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_600_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_601_n 0.00516083f $X=-0.19 $Y=1.305 $X2=5.6 $Y2=1.19
cc_111 VPB N_VPWR_c_602_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_603_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_604_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_605_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_606_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_607_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_608_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_609_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_610_n 0.0112126f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_611_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_612_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_613_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_579_n 0.0533504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_615_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_616_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_617_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_618_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_619_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_Y_c_757_n 0.0015125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_Y_c_755_n 0.00103664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB Y 0.00161879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 N_B_c_143_n N_A_c_384_n 0.0164694f $X=5.69 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_133 N_B_c_157_n N_A_c_397_n 0.0230419f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B_c_144_n N_A_c_396_n 0.00120069f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_135 N_B_c_145_n N_A_c_396_n 0.0164694f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_136 N_B_c_146_n N_VPWR_c_581_n 0.00354866f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B_c_144_n N_VPWR_c_581_n 0.00274043f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_138 N_B_c_145_n N_VPWR_c_581_n 0.00123428f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_139 N_B_c_147_n N_VPWR_c_582_n 0.00173895f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B_c_148_n N_VPWR_c_582_n 0.00173895f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B_c_148_n N_VPWR_c_583_n 0.00673617f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B_c_149_n N_VPWR_c_583_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B_c_149_n N_VPWR_c_584_n 0.00173895f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B_c_150_n N_VPWR_c_584_n 0.00173895f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B_c_150_n N_VPWR_c_585_n 0.00673617f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B_c_151_n N_VPWR_c_585_n 0.00673617f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B_c_151_n N_VPWR_c_586_n 0.00173895f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B_c_152_n N_VPWR_c_586_n 0.00173895f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B_c_152_n N_VPWR_c_587_n 0.00673617f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B_c_153_n N_VPWR_c_587_n 0.00673617f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B_c_153_n N_VPWR_c_588_n 0.00173895f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B_c_154_n N_VPWR_c_588_n 0.00173895f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_153 N_B_c_154_n N_VPWR_c_589_n 0.00673617f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_154 N_B_c_155_n N_VPWR_c_589_n 0.00673617f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B_c_155_n N_VPWR_c_590_n 0.00173895f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_156 N_B_c_156_n N_VPWR_c_590_n 0.00173895f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_157 N_B_c_157_n N_VPWR_c_591_n 0.00173895f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_158 N_B_c_156_n N_VPWR_c_598_n 0.00673617f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_159 N_B_c_157_n N_VPWR_c_598_n 0.00673617f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_160 N_B_c_146_n N_VPWR_c_613_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_161 N_B_c_147_n N_VPWR_c_613_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_162 N_B_c_146_n N_VPWR_c_579_n 0.0126298f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_163 N_B_c_147_n N_VPWR_c_579_n 0.0117184f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_164 N_B_c_148_n N_VPWR_c_579_n 0.0117184f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B_c_149_n N_VPWR_c_579_n 0.0117184f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B_c_150_n N_VPWR_c_579_n 0.0117184f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_167 N_B_c_151_n N_VPWR_c_579_n 0.0117184f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_168 N_B_c_152_n N_VPWR_c_579_n 0.0117184f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B_c_153_n N_VPWR_c_579_n 0.0117184f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B_c_154_n N_VPWR_c_579_n 0.0117184f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_171 N_B_c_155_n N_VPWR_c_579_n 0.0117184f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B_c_156_n N_VPWR_c_579_n 0.0117184f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_173 N_B_c_157_n N_VPWR_c_579_n 0.0117436f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B_c_146_n N_Y_c_760_n 0.00215964f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B_c_147_n N_Y_c_760_n 5.79575e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_176 N_B_c_144_n N_Y_c_760_n 0.0215641f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B_c_145_n N_Y_c_760_n 0.00631893f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_178 N_B_c_146_n N_Y_c_764_n 0.00897418f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B_c_147_n N_Y_c_764_n 0.0100233f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B_c_148_n N_Y_c_764_n 5.91934e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_181 N_B_c_147_n N_Y_c_767_n 0.0137916f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B_c_148_n N_Y_c_767_n 0.0137916f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B_c_144_n N_Y_c_767_n 0.0393642f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_184 N_B_c_145_n N_Y_c_767_n 0.00655651f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_185 N_B_c_147_n N_Y_c_771_n 5.91934e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B_c_148_n N_Y_c_771_n 0.0100233f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_187 N_B_c_149_n N_Y_c_771_n 0.0100233f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B_c_150_n N_Y_c_771_n 5.91934e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_189 N_B_c_149_n N_Y_c_775_n 0.0137916f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_190 N_B_c_150_n N_Y_c_775_n 0.0137916f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B_c_144_n N_Y_c_775_n 0.0393642f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_192 N_B_c_145_n N_Y_c_775_n 0.00655651f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_193 N_B_c_149_n N_Y_c_779_n 5.91934e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B_c_150_n N_Y_c_779_n 0.0100233f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_195 N_B_c_151_n N_Y_c_779_n 0.0100233f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B_c_152_n N_Y_c_779_n 5.91934e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B_c_151_n N_Y_c_783_n 0.0137916f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B_c_152_n N_Y_c_783_n 0.0137916f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B_c_144_n N_Y_c_783_n 0.0393642f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B_c_145_n N_Y_c_783_n 0.00655651f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_201 N_B_c_151_n N_Y_c_787_n 5.91934e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_152_n N_Y_c_787_n 0.0100233f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B_c_153_n N_Y_c_787_n 0.0100233f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_154_n N_Y_c_787_n 5.91934e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B_c_153_n N_Y_c_791_n 0.0137916f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B_c_154_n N_Y_c_791_n 0.0137916f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B_c_144_n N_Y_c_791_n 0.0393642f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B_c_145_n N_Y_c_791_n 0.00655651f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_209 N_B_c_153_n N_Y_c_795_n 5.91934e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B_c_154_n N_Y_c_795_n 0.0100233f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B_c_155_n N_Y_c_795_n 0.0100233f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_212 N_B_c_156_n N_Y_c_795_n 5.91934e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_213 N_B_c_155_n N_Y_c_799_n 0.0137916f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B_c_156_n N_Y_c_799_n 0.0137916f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_215 N_B_c_144_n N_Y_c_799_n 0.0393642f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_216 N_B_c_145_n N_Y_c_799_n 0.00655651f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_217 N_B_c_155_n N_Y_c_803_n 5.91934e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B_c_156_n N_Y_c_803_n 0.0100233f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B_c_157_n N_Y_c_803_n 0.0100233f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_220 N_B_c_157_n N_Y_c_806_n 0.0137485f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_221 N_B_c_144_n N_Y_c_806_n 0.0115742f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B_c_157_n N_Y_c_808_n 5.91934e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B_c_148_n N_Y_c_809_n 5.79575e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_224 N_B_c_149_n N_Y_c_809_n 5.79575e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B_c_144_n N_Y_c_809_n 0.0215641f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_226 N_B_c_145_n N_Y_c_809_n 0.00631893f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_227 N_B_c_150_n N_Y_c_813_n 5.79575e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_228 N_B_c_151_n N_Y_c_813_n 5.79575e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B_c_144_n N_Y_c_813_n 0.0215641f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_230 N_B_c_145_n N_Y_c_813_n 0.00631893f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_231 N_B_c_152_n N_Y_c_817_n 5.79575e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_232 N_B_c_153_n N_Y_c_817_n 5.79575e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_233 N_B_c_144_n N_Y_c_817_n 0.0215641f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_234 N_B_c_145_n N_Y_c_817_n 0.00631893f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_235 N_B_c_154_n N_Y_c_821_n 5.79575e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_236 N_B_c_155_n N_Y_c_821_n 5.79575e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B_c_144_n N_Y_c_821_n 0.0215641f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_238 N_B_c_145_n N_Y_c_821_n 0.00631893f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_239 N_B_c_156_n N_Y_c_825_n 5.79575e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_240 N_B_c_157_n N_Y_c_825_n 5.79575e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_241 N_B_c_144_n N_Y_c_825_n 0.0215641f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_242 N_B_c_145_n N_Y_c_825_n 0.00631893f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_243 N_B_c_157_n Y 5.27102e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B_c_144_n Y 0.0145331f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_245 N_B_c_145_n Y 8.80121e-19 $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_246 N_B_c_143_n N_Y_c_756_n 8.84206e-19 $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_247 N_B_c_132_n N_A_27_47#_c_1006_n 0.00661134f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B_c_133_n N_A_27_47#_c_1006_n 5.22294e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B_c_132_n N_A_27_47#_c_1018_n 0.00899636f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B_c_133_n N_A_27_47#_c_1018_n 0.00899636f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B_c_144_n N_A_27_47#_c_1018_n 0.0395582f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_252 N_B_c_145_n N_A_27_47#_c_1018_n 0.00457246f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_253 N_B_c_132_n N_A_27_47#_c_1007_n 8.68782e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_254 N_B_c_144_n N_A_27_47#_c_1007_n 0.00463142f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B_c_145_n N_A_27_47#_c_1007_n 0.00130673f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_256 N_B_c_132_n N_A_27_47#_c_1025_n 5.22365e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_257 N_B_c_133_n N_A_27_47#_c_1025_n 0.00661134f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B_c_134_n N_A_27_47#_c_1025_n 0.00661134f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_259 N_B_c_135_n N_A_27_47#_c_1025_n 5.22365e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_260 N_B_c_134_n N_A_27_47#_c_1029_n 0.00899636f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_261 N_B_c_135_n N_A_27_47#_c_1029_n 0.00899636f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_262 N_B_c_144_n N_A_27_47#_c_1029_n 0.0395582f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B_c_145_n N_A_27_47#_c_1029_n 0.00457246f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_264 N_B_c_134_n N_A_27_47#_c_1033_n 5.22365e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_265 N_B_c_135_n N_A_27_47#_c_1033_n 0.00661134f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_266 N_B_c_136_n N_A_27_47#_c_1033_n 0.00661134f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_267 N_B_c_137_n N_A_27_47#_c_1033_n 5.22365e-19 $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_268 N_B_c_136_n N_A_27_47#_c_1037_n 0.00899636f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B_c_137_n N_A_27_47#_c_1037_n 0.00899636f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B_c_144_n N_A_27_47#_c_1037_n 0.0395582f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_271 N_B_c_145_n N_A_27_47#_c_1037_n 0.00457246f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_272 N_B_c_136_n N_A_27_47#_c_1041_n 5.22365e-19 $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_273 N_B_c_137_n N_A_27_47#_c_1041_n 0.00661134f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_274 N_B_c_138_n N_A_27_47#_c_1041_n 0.00661134f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_275 N_B_c_139_n N_A_27_47#_c_1041_n 5.22365e-19 $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_276 N_B_c_138_n N_A_27_47#_c_1045_n 0.00899636f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_277 N_B_c_139_n N_A_27_47#_c_1045_n 0.00899636f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B_c_144_n N_A_27_47#_c_1045_n 0.0395582f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_279 N_B_c_145_n N_A_27_47#_c_1045_n 0.00457246f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_280 N_B_c_138_n N_A_27_47#_c_1049_n 5.22365e-19 $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_281 N_B_c_139_n N_A_27_47#_c_1049_n 0.00661134f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B_c_140_n N_A_27_47#_c_1049_n 0.00661134f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B_c_141_n N_A_27_47#_c_1049_n 5.22365e-19 $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B_c_140_n N_A_27_47#_c_1053_n 0.00899636f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B_c_141_n N_A_27_47#_c_1053_n 0.00899636f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B_c_144_n N_A_27_47#_c_1053_n 0.0395582f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_287 N_B_c_145_n N_A_27_47#_c_1053_n 0.00457246f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_288 N_B_c_140_n N_A_27_47#_c_1057_n 5.22365e-19 $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B_c_141_n N_A_27_47#_c_1057_n 0.00661134f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B_c_142_n N_A_27_47#_c_1057_n 0.00661134f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B_c_143_n N_A_27_47#_c_1057_n 5.22365e-19 $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B_c_142_n N_A_27_47#_c_1061_n 0.00899636f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B_c_143_n N_A_27_47#_c_1061_n 0.00899636f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B_c_144_n N_A_27_47#_c_1061_n 0.0395582f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_295 N_B_c_145_n N_A_27_47#_c_1061_n 0.00457246f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_296 N_B_c_143_n N_A_27_47#_c_1065_n 0.00248145f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B_c_142_n N_A_27_47#_c_1008_n 4.7541e-19 $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_298 N_B_c_143_n N_A_27_47#_c_1008_n 0.00502046f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B_c_144_n N_A_27_47#_c_1008_n 0.00230426f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_300 N_B_c_133_n N_A_27_47#_c_1011_n 8.68782e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B_c_134_n N_A_27_47#_c_1011_n 8.68782e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B_c_144_n N_A_27_47#_c_1011_n 0.0214029f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_303 N_B_c_145_n N_A_27_47#_c_1011_n 0.00224547f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_304 N_B_c_135_n N_A_27_47#_c_1012_n 8.68782e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_305 N_B_c_136_n N_A_27_47#_c_1012_n 8.68782e-19 $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B_c_144_n N_A_27_47#_c_1012_n 0.0214029f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_307 N_B_c_145_n N_A_27_47#_c_1012_n 0.00224547f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_308 N_B_c_137_n N_A_27_47#_c_1013_n 8.68782e-19 $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_309 N_B_c_138_n N_A_27_47#_c_1013_n 8.68782e-19 $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_310 N_B_c_144_n N_A_27_47#_c_1013_n 0.0214029f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_311 N_B_c_145_n N_A_27_47#_c_1013_n 0.00224547f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_312 N_B_c_139_n N_A_27_47#_c_1014_n 8.68782e-19 $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_313 N_B_c_140_n N_A_27_47#_c_1014_n 8.68782e-19 $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_314 N_B_c_144_n N_A_27_47#_c_1014_n 0.0214029f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_315 N_B_c_145_n N_A_27_47#_c_1014_n 0.00224547f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_316 N_B_c_141_n N_A_27_47#_c_1015_n 8.68782e-19 $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B_c_142_n N_A_27_47#_c_1015_n 8.68782e-19 $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B_c_144_n N_A_27_47#_c_1015_n 0.0214029f $X=5.6 $Y=1.16 $X2=0 $Y2=0
cc_319 N_B_c_145_n N_A_27_47#_c_1015_n 0.00224547f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_320 N_B_c_132_n N_VGND_c_1182_n 0.00296353f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_321 N_B_c_133_n N_VGND_c_1182_n 0.00166854f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_322 N_B_c_133_n N_VGND_c_1183_n 0.00422241f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_323 N_B_c_134_n N_VGND_c_1183_n 0.00422241f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_324 N_B_c_134_n N_VGND_c_1184_n 0.00166854f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_325 N_B_c_135_n N_VGND_c_1184_n 0.00166854f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_326 N_B_c_135_n N_VGND_c_1185_n 0.00422241f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_327 N_B_c_136_n N_VGND_c_1185_n 0.00422241f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_328 N_B_c_136_n N_VGND_c_1186_n 0.00166854f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B_c_137_n N_VGND_c_1186_n 0.00166854f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_330 N_B_c_137_n N_VGND_c_1187_n 0.00422241f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_331 N_B_c_138_n N_VGND_c_1187_n 0.00422241f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_332 N_B_c_138_n N_VGND_c_1188_n 0.00166854f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_333 N_B_c_139_n N_VGND_c_1188_n 0.00166854f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_334 N_B_c_139_n N_VGND_c_1189_n 0.00422241f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_335 N_B_c_140_n N_VGND_c_1189_n 0.00422241f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_336 N_B_c_140_n N_VGND_c_1190_n 0.00166854f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_337 N_B_c_141_n N_VGND_c_1190_n 0.00166854f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_338 N_B_c_142_n N_VGND_c_1191_n 0.00166854f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_339 N_B_c_143_n N_VGND_c_1191_n 0.00296353f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_340 N_B_c_141_n N_VGND_c_1192_n 0.00422241f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_341 N_B_c_142_n N_VGND_c_1192_n 0.00422241f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_342 N_B_c_132_n N_VGND_c_1194_n 0.00422241f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_343 N_B_c_143_n N_VGND_c_1195_n 0.00420723f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_344 N_B_c_132_n N_VGND_c_1196_n 0.00689308f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_345 N_B_c_133_n N_VGND_c_1196_n 0.00593887f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_346 N_B_c_134_n N_VGND_c_1196_n 0.00593887f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_347 N_B_c_135_n N_VGND_c_1196_n 0.00593887f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_348 N_B_c_136_n N_VGND_c_1196_n 0.00593887f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_349 N_B_c_137_n N_VGND_c_1196_n 0.00593887f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_350 N_B_c_138_n N_VGND_c_1196_n 0.00593887f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_351 N_B_c_139_n N_VGND_c_1196_n 0.00593887f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_352 N_B_c_140_n N_VGND_c_1196_n 0.00593887f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_353 N_B_c_141_n N_VGND_c_1196_n 0.00593887f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_354 N_B_c_142_n N_VGND_c_1196_n 0.00593887f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_355 N_B_c_143_n N_VGND_c_1196_n 0.00597515f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_356 N_A_c_397_n N_VPWR_c_591_n 0.00173895f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_357 N_A_c_398_n N_VPWR_c_592_n 0.00173895f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_358 N_A_c_399_n N_VPWR_c_592_n 0.00173895f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_359 N_A_c_400_n N_VPWR_c_593_n 0.00173895f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_360 N_A_c_401_n N_VPWR_c_593_n 0.00173895f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_361 N_A_c_402_n N_VPWR_c_594_n 0.00173895f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_362 N_A_c_403_n N_VPWR_c_594_n 0.00173895f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_363 N_A_c_404_n N_VPWR_c_595_n 0.00173895f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_364 N_A_c_405_n N_VPWR_c_595_n 0.00173895f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_365 N_A_c_406_n N_VPWR_c_596_n 0.00173895f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_366 N_A_c_407_n N_VPWR_c_596_n 0.00173895f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_367 N_A_c_408_n N_VPWR_c_597_n 0.00354866f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_368 N_A_c_397_n N_VPWR_c_600_n 0.00673617f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_369 N_A_c_398_n N_VPWR_c_600_n 0.00673617f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_370 N_A_c_399_n N_VPWR_c_602_n 0.00673617f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_371 N_A_c_400_n N_VPWR_c_602_n 0.00673617f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_372 N_A_c_401_n N_VPWR_c_604_n 0.00673617f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_373 N_A_c_402_n N_VPWR_c_604_n 0.00673617f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_374 N_A_c_403_n N_VPWR_c_606_n 0.00673617f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_375 N_A_c_404_n N_VPWR_c_606_n 0.00673617f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_376 N_A_c_405_n N_VPWR_c_608_n 0.00673617f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_377 N_A_c_406_n N_VPWR_c_608_n 0.00673617f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_378 N_A_c_407_n N_VPWR_c_611_n 0.00673617f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_379 N_A_c_408_n N_VPWR_c_611_n 0.00673617f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_380 N_A_c_397_n N_VPWR_c_579_n 0.0117436f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_381 N_A_c_398_n N_VPWR_c_579_n 0.0117184f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_382 N_A_c_399_n N_VPWR_c_579_n 0.0117184f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_383 N_A_c_400_n N_VPWR_c_579_n 0.0117184f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_384 N_A_c_401_n N_VPWR_c_579_n 0.0117184f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_385 N_A_c_402_n N_VPWR_c_579_n 0.0117184f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_386 N_A_c_403_n N_VPWR_c_579_n 0.0117184f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_387 N_A_c_404_n N_VPWR_c_579_n 0.0117184f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_388 N_A_c_405_n N_VPWR_c_579_n 0.0117184f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_389 N_A_c_406_n N_VPWR_c_579_n 0.0117184f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_390 N_A_c_407_n N_VPWR_c_579_n 0.0117184f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_391 N_A_c_408_n N_VPWR_c_579_n 0.0127482f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_392 N_A_c_397_n N_Y_c_803_n 5.91934e-19 $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_393 N_A_c_384_n N_Y_c_834_n 0.00303037f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_394 N_A_c_397_n N_Y_c_808_n 0.0100233f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_395 N_A_c_398_n N_Y_c_808_n 0.0100233f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_396 N_A_c_399_n N_Y_c_808_n 5.91934e-19 $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_397 N_A_c_385_n N_Y_c_838_n 0.0124451f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_398 N_A_c_386_n N_Y_c_838_n 0.0109111f $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_399 N_A_c_387_n N_Y_c_838_n 0.0104739f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_400 N_A_c_388_n N_Y_c_838_n 0.0104739f $X=7.99 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A_c_389_n N_Y_c_838_n 0.0104739f $X=8.51 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A_c_390_n N_Y_c_838_n 0.0104739f $X=8.93 $Y=0.995 $X2=0 $Y2=0
cc_403 N_A_c_391_n N_Y_c_838_n 0.0109111f $X=9.4 $Y=0.995 $X2=0 $Y2=0
cc_404 N_A_c_392_n N_Y_c_838_n 0.0109111f $X=9.87 $Y=0.995 $X2=0 $Y2=0
cc_405 N_A_c_393_n N_Y_c_838_n 0.0104739f $X=10.39 $Y=0.995 $X2=0 $Y2=0
cc_406 N_A_c_394_n N_Y_c_838_n 0.0123979f $X=10.81 $Y=0.995 $X2=0 $Y2=0
cc_407 N_A_c_465_p N_Y_c_838_n 0.263367f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_408 N_A_c_396_n N_Y_c_838_n 0.0306126f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_409 N_A_c_398_n N_Y_c_850_n 0.014973f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_410 N_A_c_399_n N_Y_c_850_n 0.0137916f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_411 N_A_c_465_p N_Y_c_850_n 0.0330732f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_412 N_A_c_396_n N_Y_c_850_n 0.00635951f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_413 N_A_c_398_n N_Y_c_854_n 5.91934e-19 $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_414 N_A_c_399_n N_Y_c_854_n 0.0100233f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_415 N_A_c_400_n N_Y_c_854_n 0.0100233f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_416 N_A_c_401_n N_Y_c_854_n 5.91934e-19 $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_417 N_A_c_400_n N_Y_c_858_n 0.0137916f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_418 N_A_c_401_n N_Y_c_858_n 0.0137916f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_419 N_A_c_465_p N_Y_c_858_n 0.0393642f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_420 N_A_c_396_n N_Y_c_858_n 0.00655651f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_421 N_A_c_400_n N_Y_c_862_n 5.91934e-19 $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_422 N_A_c_401_n N_Y_c_862_n 0.0100233f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_423 N_A_c_402_n N_Y_c_862_n 0.0100233f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_424 N_A_c_403_n N_Y_c_862_n 5.91934e-19 $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_425 N_A_c_402_n N_Y_c_866_n 0.0137916f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_426 N_A_c_403_n N_Y_c_866_n 0.0137916f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_427 N_A_c_465_p N_Y_c_866_n 0.0393642f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_428 N_A_c_396_n N_Y_c_866_n 0.00655651f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_429 N_A_c_402_n N_Y_c_870_n 5.91934e-19 $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_430 N_A_c_403_n N_Y_c_870_n 0.0100233f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_431 N_A_c_404_n N_Y_c_870_n 0.0100233f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_432 N_A_c_405_n N_Y_c_870_n 5.91934e-19 $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_433 N_A_c_404_n N_Y_c_874_n 0.0137916f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_434 N_A_c_405_n N_Y_c_874_n 0.0137916f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_435 N_A_c_465_p N_Y_c_874_n 0.0393642f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_436 N_A_c_396_n N_Y_c_874_n 0.00635951f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_437 N_A_c_404_n N_Y_c_878_n 5.91934e-19 $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_438 N_A_c_405_n N_Y_c_878_n 0.0100233f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_439 N_A_c_406_n N_Y_c_878_n 0.0100233f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_440 N_A_c_407_n N_Y_c_878_n 5.91934e-19 $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_441 N_A_c_406_n N_Y_c_882_n 0.0137916f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_442 N_A_c_407_n N_Y_c_882_n 0.0159022f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_443 N_A_c_465_p N_Y_c_882_n 0.0263345f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_444 N_A_c_396_n N_Y_c_882_n 0.00655651f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_445 N_A_c_406_n N_Y_c_886_n 5.91934e-19 $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_446 N_A_c_407_n N_Y_c_886_n 0.0100233f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_447 N_A_c_408_n N_Y_c_886_n 0.00897418f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_448 N_A_c_407_n N_Y_c_757_n 0.0019905f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_449 N_A_c_408_n N_Y_c_757_n 0.00423504f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_450 N_A_c_396_n N_Y_c_757_n 0.00694896f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_451 N_A_c_397_n N_Y_c_892_n 0.0130984f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_452 N_A_c_398_n N_Y_c_892_n 8.15944e-19 $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_453 N_A_c_396_n N_Y_c_892_n 0.00123735f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_454 N_A_c_399_n N_Y_c_895_n 5.79575e-19 $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_455 N_A_c_400_n N_Y_c_895_n 5.79575e-19 $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_456 N_A_c_465_p N_Y_c_895_n 0.0215641f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_457 N_A_c_396_n N_Y_c_895_n 0.00631893f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_458 N_A_c_401_n N_Y_c_899_n 5.79575e-19 $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_459 N_A_c_402_n N_Y_c_899_n 5.79575e-19 $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_460 N_A_c_465_p N_Y_c_899_n 0.0215641f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_461 N_A_c_396_n N_Y_c_899_n 0.00631893f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_462 N_A_c_403_n N_Y_c_903_n 5.79575e-19 $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_463 N_A_c_404_n N_Y_c_903_n 5.79575e-19 $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_464 N_A_c_465_p N_Y_c_903_n 0.0215641f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_465 N_A_c_396_n N_Y_c_903_n 0.00651614f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_466 N_A_c_405_n N_Y_c_907_n 5.79575e-19 $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_467 N_A_c_406_n N_Y_c_907_n 5.79575e-19 $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_468 N_A_c_465_p N_Y_c_907_n 0.0215641f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_469 N_A_c_396_n N_Y_c_907_n 0.00631893f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_470 N_A_c_407_n N_Y_c_911_n 8.15944e-19 $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_471 N_A_c_408_n N_Y_c_911_n 0.00188422f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_472 N_A_c_394_n N_Y_c_754_n 0.00286869f $X=10.81 $Y=0.995 $X2=0 $Y2=0
cc_473 N_A_c_395_n N_Y_c_754_n 0.0031043f $X=11.33 $Y=0.995 $X2=0 $Y2=0
cc_474 N_A_c_396_n N_Y_c_754_n 0.0106358f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_475 N_A_c_465_p N_Y_c_755_n 0.0151436f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_476 N_A_c_396_n N_Y_c_755_n 0.0384565f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_477 N_A_c_397_n Y 0.00326841f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_478 N_A_c_398_n Y 0.00234191f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_479 N_A_c_465_p Y 0.0216953f $X=10.53 $Y=1.16 $X2=0 $Y2=0
cc_480 N_A_c_396_n Y 0.0307267f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_481 N_A_c_384_n N_Y_c_756_n 0.00315482f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_482 N_A_c_385_n N_Y_c_756_n 0.00297134f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_483 N_A_c_396_n N_Y_c_756_n 0.00830622f $X=11.305 $Y=1.202 $X2=0 $Y2=0
cc_484 N_A_c_384_n N_A_27_47#_c_1089_n 0.0108171f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_485 N_A_c_385_n N_A_27_47#_c_1089_n 0.00903374f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_486 N_A_c_386_n N_A_27_47#_c_1089_n 0.00935436f $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_487 N_A_c_387_n N_A_27_47#_c_1089_n 0.00935436f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_488 N_A_c_388_n N_A_27_47#_c_1089_n 0.00935436f $X=7.99 $Y=0.995 $X2=0 $Y2=0
cc_489 N_A_c_389_n N_A_27_47#_c_1089_n 0.00935436f $X=8.51 $Y=0.995 $X2=0 $Y2=0
cc_490 N_A_c_390_n N_A_27_47#_c_1089_n 0.00903374f $X=8.93 $Y=0.995 $X2=0 $Y2=0
cc_491 N_A_c_391_n N_A_27_47#_c_1089_n 0.00903374f $X=9.4 $Y=0.995 $X2=0 $Y2=0
cc_492 N_A_c_392_n N_A_27_47#_c_1089_n 0.00935436f $X=9.87 $Y=0.995 $X2=0 $Y2=0
cc_493 N_A_c_393_n N_A_27_47#_c_1089_n 0.00935436f $X=10.39 $Y=0.995 $X2=0 $Y2=0
cc_494 N_A_c_394_n N_A_27_47#_c_1089_n 0.00935436f $X=10.81 $Y=0.995 $X2=0 $Y2=0
cc_495 N_A_c_395_n N_A_27_47#_c_1089_n 0.0113632f $X=11.33 $Y=0.995 $X2=0 $Y2=0
cc_496 N_A_c_396_n N_A_27_47#_c_1089_n 0.00110461f $X=11.305 $Y=1.202 $X2=0
+ $Y2=0
cc_497 N_A_c_384_n N_VGND_c_1195_n 0.00357877f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_498 N_A_c_385_n N_VGND_c_1195_n 0.00357877f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_499 N_A_c_386_n N_VGND_c_1195_n 0.00357877f $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_500 N_A_c_387_n N_VGND_c_1195_n 0.00357877f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_501 N_A_c_388_n N_VGND_c_1195_n 0.00357877f $X=7.99 $Y=0.995 $X2=0 $Y2=0
cc_502 N_A_c_389_n N_VGND_c_1195_n 0.00357877f $X=8.51 $Y=0.995 $X2=0 $Y2=0
cc_503 N_A_c_390_n N_VGND_c_1195_n 0.00357877f $X=8.93 $Y=0.995 $X2=0 $Y2=0
cc_504 N_A_c_391_n N_VGND_c_1195_n 0.00357877f $X=9.4 $Y=0.995 $X2=0 $Y2=0
cc_505 N_A_c_392_n N_VGND_c_1195_n 0.00357877f $X=9.87 $Y=0.995 $X2=0 $Y2=0
cc_506 N_A_c_393_n N_VGND_c_1195_n 0.00357877f $X=10.39 $Y=0.995 $X2=0 $Y2=0
cc_507 N_A_c_394_n N_VGND_c_1195_n 0.00357877f $X=10.81 $Y=0.995 $X2=0 $Y2=0
cc_508 N_A_c_395_n N_VGND_c_1195_n 0.00357877f $X=11.33 $Y=0.995 $X2=0 $Y2=0
cc_509 N_A_c_384_n N_VGND_c_1196_n 0.00538422f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_510 N_A_c_385_n N_VGND_c_1196_n 0.00548399f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_511 N_A_c_386_n N_VGND_c_1196_n 0.00560377f $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_512 N_A_c_387_n N_VGND_c_1196_n 0.0054768f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_513 N_A_c_388_n N_VGND_c_1196_n 0.0054768f $X=7.99 $Y=0.995 $X2=0 $Y2=0
cc_514 N_A_c_389_n N_VGND_c_1196_n 0.0054768f $X=8.51 $Y=0.995 $X2=0 $Y2=0
cc_515 N_A_c_390_n N_VGND_c_1196_n 0.00535702f $X=8.93 $Y=0.995 $X2=0 $Y2=0
cc_516 N_A_c_391_n N_VGND_c_1196_n 0.00548399f $X=9.4 $Y=0.995 $X2=0 $Y2=0
cc_517 N_A_c_392_n N_VGND_c_1196_n 0.00560377f $X=9.87 $Y=0.995 $X2=0 $Y2=0
cc_518 N_A_c_393_n N_VGND_c_1196_n 0.0054768f $X=10.39 $Y=0.995 $X2=0 $Y2=0
cc_519 N_A_c_394_n N_VGND_c_1196_n 0.0054768f $X=10.81 $Y=0.995 $X2=0 $Y2=0
cc_520 N_A_c_395_n N_VGND_c_1196_n 0.00655303f $X=11.33 $Y=0.995 $X2=0 $Y2=0
cc_521 N_VPWR_c_579_n N_Y_M1000_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_522 N_VPWR_c_579_n N_Y_M1004_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_523 N_VPWR_c_579_n N_Y_M1012_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_524 N_VPWR_c_579_n N_Y_M1022_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_525 N_VPWR_c_579_n N_Y_M1029_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_526 N_VPWR_c_579_n N_Y_M1038_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_527 N_VPWR_c_579_n N_Y_M1002_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_528 N_VPWR_c_579_n N_Y_M1010_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_529 N_VPWR_c_579_n N_Y_M1020_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_530 N_VPWR_c_579_n N_Y_M1030_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_531 N_VPWR_c_579_n N_Y_M1037_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_532 N_VPWR_c_579_n N_Y_M1046_s 0.00231261f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_533 N_VPWR_c_613_n N_Y_c_764_n 0.0189467f $X=1.065 $Y=2.72 $X2=0 $Y2=0
cc_534 N_VPWR_c_579_n N_Y_c_764_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_535 N_VPWR_M1001_d N_Y_c_767_n 0.00334388f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_536 N_VPWR_c_582_n N_Y_c_767_n 0.0143191f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_537 N_VPWR_c_583_n N_Y_c_771_n 0.0189467f $X=2.005 $Y=2.72 $X2=0 $Y2=0
cc_538 N_VPWR_c_579_n N_Y_c_771_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_539 N_VPWR_M1005_d N_Y_c_775_n 0.00334388f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_540 N_VPWR_c_584_n N_Y_c_775_n 0.0143191f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_541 N_VPWR_c_585_n N_Y_c_779_n 0.0189467f $X=2.945 $Y=2.72 $X2=0 $Y2=0
cc_542 N_VPWR_c_579_n N_Y_c_779_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_543 N_VPWR_M1015_d N_Y_c_783_n 0.00334388f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_544 N_VPWR_c_586_n N_Y_c_783_n 0.0143191f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_545 N_VPWR_c_587_n N_Y_c_787_n 0.0189467f $X=3.885 $Y=2.72 $X2=0 $Y2=0
cc_546 N_VPWR_c_579_n N_Y_c_787_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_547 N_VPWR_M1025_d N_Y_c_791_n 0.00334388f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_548 N_VPWR_c_588_n N_Y_c_791_n 0.0143191f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_549 N_VPWR_c_589_n N_Y_c_795_n 0.0189467f $X=4.825 $Y=2.72 $X2=0 $Y2=0
cc_550 N_VPWR_c_579_n N_Y_c_795_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_551 N_VPWR_M1033_d N_Y_c_799_n 0.00334388f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_552 N_VPWR_c_590_n N_Y_c_799_n 0.0143191f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_553 N_VPWR_c_598_n N_Y_c_803_n 0.0189467f $X=5.765 $Y=2.72 $X2=0 $Y2=0
cc_554 N_VPWR_c_579_n N_Y_c_803_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_555 N_VPWR_M1041_d N_Y_c_806_n 0.00534233f $X=5.755 $Y=1.485 $X2=0 $Y2=0
cc_556 N_VPWR_c_591_n N_Y_c_806_n 0.0143191f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_557 N_VPWR_c_600_n N_Y_c_808_n 0.0189467f $X=6.705 $Y=2.72 $X2=0 $Y2=0
cc_558 N_VPWR_c_579_n N_Y_c_808_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_559 N_VPWR_M1006_d N_Y_c_850_n 0.00334388f $X=6.695 $Y=1.485 $X2=0 $Y2=0
cc_560 N_VPWR_c_592_n N_Y_c_850_n 0.0143191f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_561 N_VPWR_c_602_n N_Y_c_854_n 0.0189467f $X=7.645 $Y=2.72 $X2=0 $Y2=0
cc_562 N_VPWR_c_579_n N_Y_c_854_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_563 N_VPWR_M1017_d N_Y_c_858_n 0.00334388f $X=7.635 $Y=1.485 $X2=0 $Y2=0
cc_564 N_VPWR_c_593_n N_Y_c_858_n 0.0143191f $X=7.78 $Y=2 $X2=0 $Y2=0
cc_565 N_VPWR_c_604_n N_Y_c_862_n 0.0189467f $X=8.585 $Y=2.72 $X2=0 $Y2=0
cc_566 N_VPWR_c_579_n N_Y_c_862_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_567 N_VPWR_M1023_d N_Y_c_866_n 0.00334388f $X=8.575 $Y=1.485 $X2=0 $Y2=0
cc_568 N_VPWR_c_594_n N_Y_c_866_n 0.0143191f $X=8.72 $Y=2 $X2=0 $Y2=0
cc_569 N_VPWR_c_606_n N_Y_c_870_n 0.0189467f $X=9.525 $Y=2.72 $X2=0 $Y2=0
cc_570 N_VPWR_c_579_n N_Y_c_870_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_571 N_VPWR_M1035_d N_Y_c_874_n 0.00334388f $X=9.515 $Y=1.485 $X2=0 $Y2=0
cc_572 N_VPWR_c_595_n N_Y_c_874_n 0.0143191f $X=9.66 $Y=2 $X2=0 $Y2=0
cc_573 N_VPWR_c_608_n N_Y_c_878_n 0.0189467f $X=10.465 $Y=2.72 $X2=0 $Y2=0
cc_574 N_VPWR_c_579_n N_Y_c_878_n 0.0123132f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_575 N_VPWR_M1039_d N_Y_c_882_n 0.00334388f $X=10.455 $Y=1.485 $X2=0 $Y2=0
cc_576 N_VPWR_c_596_n N_Y_c_882_n 0.0143191f $X=10.6 $Y=2 $X2=0 $Y2=0
cc_577 N_VPWR_c_611_n N_Y_c_886_n 0.0189467f $X=11.405 $Y=2.72 $X2=0 $Y2=0
cc_578 N_VPWR_c_579_n N_Y_c_886_n 0.0123027f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_579 N_VPWR_c_581_n N_A_27_47#_c_1007_n 0.0071931f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_580 N_VPWR_c_597_n N_A_27_47#_c_1010_n 0.00739919f $X=11.54 $Y=1.66 $X2=0
+ $Y2=0
cc_581 N_Y_c_838_n N_A_27_47#_M1008_s 0.00401355f $X=10.965 $Y=0.76 $X2=0 $Y2=0
cc_582 N_Y_c_838_n N_A_27_47#_M1014_s 0.00307883f $X=10.965 $Y=0.76 $X2=0 $Y2=0
cc_583 N_Y_c_838_n N_A_27_47#_M1019_s 0.00307883f $X=10.965 $Y=0.76 $X2=0 $Y2=0
cc_584 N_Y_c_838_n N_A_27_47#_M1027_s 0.00401355f $X=10.965 $Y=0.76 $X2=0 $Y2=0
cc_585 N_Y_c_838_n N_A_27_47#_M1032_s 0.00307883f $X=10.965 $Y=0.76 $X2=0 $Y2=0
cc_586 N_Y_c_806_n N_A_27_47#_c_1008_n 0.00507137f $X=6.045 $Y=1.58 $X2=0 $Y2=0
cc_587 N_Y_M1007_d N_A_27_47#_c_1089_n 0.00399738f $X=6.185 $Y=0.235 $X2=0 $Y2=0
cc_588 N_Y_M1009_d N_A_27_47#_c_1089_n 0.00507102f $X=7.125 $Y=0.235 $X2=0 $Y2=0
cc_589 N_Y_M1018_d N_A_27_47#_c_1089_n 0.00507102f $X=8.065 $Y=0.235 $X2=0 $Y2=0
cc_590 N_Y_M1024_d N_A_27_47#_c_1089_n 0.00400219f $X=9.005 $Y=0.235 $X2=0 $Y2=0
cc_591 N_Y_M1028_d N_A_27_47#_c_1089_n 0.00507102f $X=9.945 $Y=0.235 $X2=0 $Y2=0
cc_592 N_Y_M1034_d N_A_27_47#_c_1089_n 0.00506571f $X=10.885 $Y=0.235 $X2=0
+ $Y2=0
cc_593 N_Y_c_834_n N_A_27_47#_c_1089_n 0.0182216f $X=6.305 $Y=0.885 $X2=0 $Y2=0
cc_594 N_Y_c_838_n N_A_27_47#_c_1089_n 0.235458f $X=10.965 $Y=0.76 $X2=0 $Y2=0
cc_595 N_Y_c_997_p N_A_27_47#_c_1089_n 0.018174f $X=11.1 $Y=0.885 $X2=0 $Y2=0
cc_596 N_Y_c_755_n N_A_27_47#_c_1089_n 0.00458386f $X=11.2 $Y=1.325 $X2=0 $Y2=0
cc_597 Y N_A_27_47#_c_1089_n 0.00297886f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_598 N_Y_M1007_d N_VGND_c_1196_n 0.00256987f $X=6.185 $Y=0.235 $X2=0 $Y2=0
cc_599 N_Y_M1009_d N_VGND_c_1196_n 0.00297142f $X=7.125 $Y=0.235 $X2=0 $Y2=0
cc_600 N_Y_M1018_d N_VGND_c_1196_n 0.00297142f $X=8.065 $Y=0.235 $X2=0 $Y2=0
cc_601 N_Y_M1024_d N_VGND_c_1196_n 0.00256987f $X=9.005 $Y=0.235 $X2=0 $Y2=0
cc_602 N_Y_M1028_d N_VGND_c_1196_n 0.00297142f $X=9.945 $Y=0.235 $X2=0 $Y2=0
cc_603 N_Y_M1034_d N_VGND_c_1196_n 0.00297142f $X=10.885 $Y=0.235 $X2=0 $Y2=0
cc_604 N_A_27_47#_c_1018_n N_VGND_M1003_s 0.00500594f $X=1.035 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_605 N_A_27_47#_c_1029_n N_VGND_M1013_s 0.00500594f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_606 N_A_27_47#_c_1037_n N_VGND_M1021_s 0.00500594f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_607 N_A_27_47#_c_1045_n N_VGND_M1031_s 0.00500594f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_608 N_A_27_47#_c_1053_n N_VGND_M1040_s 0.00500594f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_609 N_A_27_47#_c_1061_n N_VGND_M1043_s 0.00500594f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_610 N_A_27_47#_c_1018_n N_VGND_c_1182_n 0.0199861f $X=1.035 $Y=0.8 $X2=0
+ $Y2=0
cc_611 N_A_27_47#_c_1018_n N_VGND_c_1183_n 0.0020257f $X=1.035 $Y=0.8 $X2=0
+ $Y2=0
cc_612 N_A_27_47#_c_1025_n N_VGND_c_1183_n 0.0188215f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_613 N_A_27_47#_c_1029_n N_VGND_c_1183_n 0.0020257f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_614 N_A_27_47#_c_1029_n N_VGND_c_1184_n 0.0199861f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_615 N_A_27_47#_c_1029_n N_VGND_c_1185_n 0.0020257f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_616 N_A_27_47#_c_1033_n N_VGND_c_1185_n 0.0188215f $X=2.14 $Y=0.38 $X2=0
+ $Y2=0
cc_617 N_A_27_47#_c_1037_n N_VGND_c_1185_n 0.0020257f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_618 N_A_27_47#_c_1037_n N_VGND_c_1186_n 0.0199861f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_619 N_A_27_47#_c_1037_n N_VGND_c_1187_n 0.0020257f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_620 N_A_27_47#_c_1041_n N_VGND_c_1187_n 0.0188215f $X=3.08 $Y=0.38 $X2=0
+ $Y2=0
cc_621 N_A_27_47#_c_1045_n N_VGND_c_1187_n 0.0020257f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_622 N_A_27_47#_c_1045_n N_VGND_c_1188_n 0.0199861f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_623 N_A_27_47#_c_1045_n N_VGND_c_1189_n 0.0020257f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_624 N_A_27_47#_c_1049_n N_VGND_c_1189_n 0.0188215f $X=4.02 $Y=0.38 $X2=0
+ $Y2=0
cc_625 N_A_27_47#_c_1053_n N_VGND_c_1189_n 0.0020257f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_626 N_A_27_47#_c_1053_n N_VGND_c_1190_n 0.0199861f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_627 N_A_27_47#_c_1061_n N_VGND_c_1191_n 0.0199861f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_628 N_A_27_47#_c_1053_n N_VGND_c_1192_n 0.0020257f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_629 N_A_27_47#_c_1057_n N_VGND_c_1192_n 0.0188215f $X=4.96 $Y=0.38 $X2=0
+ $Y2=0
cc_630 N_A_27_47#_c_1061_n N_VGND_c_1192_n 0.0020257f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_631 N_A_27_47#_c_1006_n N_VGND_c_1194_n 0.0212882f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_632 N_A_27_47#_c_1018_n N_VGND_c_1194_n 0.0020257f $X=1.035 $Y=0.8 $X2=0
+ $Y2=0
cc_633 N_A_27_47#_c_1061_n N_VGND_c_1195_n 0.0020257f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_634 N_A_27_47#_c_1065_n N_VGND_c_1195_n 0.0151813f $X=5.86 $Y=0.465 $X2=0
+ $Y2=0
cc_635 N_A_27_47#_c_1089_n N_VGND_c_1195_n 0.308632f $X=11.455 $Y=0.36 $X2=0
+ $Y2=0
cc_636 N_A_27_47#_c_1009_n N_VGND_c_1195_n 0.0172955f $X=11.58 $Y=0.465 $X2=0
+ $Y2=0
cc_637 N_A_27_47#_M1003_d N_VGND_c_1196_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_638 N_A_27_47#_M1011_d N_VGND_c_1196_n 0.00215201f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_639 N_A_27_47#_M1016_d N_VGND_c_1196_n 0.00215201f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_640 N_A_27_47#_M1026_d N_VGND_c_1196_n 0.00215201f $X=2.945 $Y=0.235 $X2=0
+ $Y2=0
cc_641 N_A_27_47#_M1036_d N_VGND_c_1196_n 0.00215201f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_642 N_A_27_47#_M1042_d N_VGND_c_1196_n 0.00215201f $X=4.825 $Y=0.235 $X2=0
+ $Y2=0
cc_643 N_A_27_47#_M1044_d N_VGND_c_1196_n 0.00215206f $X=5.765 $Y=0.235 $X2=0
+ $Y2=0
cc_644 N_A_27_47#_M1008_s N_VGND_c_1196_n 0.00255381f $X=6.655 $Y=0.235 $X2=0
+ $Y2=0
cc_645 N_A_27_47#_M1014_s N_VGND_c_1196_n 0.00215227f $X=7.645 $Y=0.235 $X2=0
+ $Y2=0
cc_646 N_A_27_47#_M1019_s N_VGND_c_1196_n 0.00215227f $X=8.585 $Y=0.235 $X2=0
+ $Y2=0
cc_647 N_A_27_47#_M1027_s N_VGND_c_1196_n 0.00255381f $X=9.475 $Y=0.235 $X2=0
+ $Y2=0
cc_648 N_A_27_47#_M1032_s N_VGND_c_1196_n 0.00215227f $X=10.465 $Y=0.235 $X2=0
+ $Y2=0
cc_649 N_A_27_47#_M1045_s N_VGND_c_1196_n 0.00209324f $X=11.405 $Y=0.235 $X2=0
+ $Y2=0
cc_650 N_A_27_47#_c_1006_n N_VGND_c_1196_n 0.0125939f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_651 N_A_27_47#_c_1018_n N_VGND_c_1196_n 0.00880092f $X=1.035 $Y=0.8 $X2=0
+ $Y2=0
cc_652 N_A_27_47#_c_1025_n N_VGND_c_1196_n 0.0121968f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_653 N_A_27_47#_c_1029_n N_VGND_c_1196_n 0.00880092f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_654 N_A_27_47#_c_1033_n N_VGND_c_1196_n 0.0121968f $X=2.14 $Y=0.38 $X2=0
+ $Y2=0
cc_655 N_A_27_47#_c_1037_n N_VGND_c_1196_n 0.00880092f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_656 N_A_27_47#_c_1041_n N_VGND_c_1196_n 0.0121968f $X=3.08 $Y=0.38 $X2=0
+ $Y2=0
cc_657 N_A_27_47#_c_1045_n N_VGND_c_1196_n 0.00880092f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_658 N_A_27_47#_c_1049_n N_VGND_c_1196_n 0.0121968f $X=4.02 $Y=0.38 $X2=0
+ $Y2=0
cc_659 N_A_27_47#_c_1053_n N_VGND_c_1196_n 0.00880092f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_660 N_A_27_47#_c_1057_n N_VGND_c_1196_n 0.0121968f $X=4.96 $Y=0.38 $X2=0
+ $Y2=0
cc_661 N_A_27_47#_c_1061_n N_VGND_c_1196_n 0.00880092f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_662 N_A_27_47#_c_1065_n N_VGND_c_1196_n 0.0093992f $X=5.86 $Y=0.465 $X2=0
+ $Y2=0
cc_663 N_A_27_47#_c_1089_n N_VGND_c_1196_n 0.195611f $X=11.455 $Y=0.36 $X2=0
+ $Y2=0
cc_664 N_A_27_47#_c_1009_n N_VGND_c_1196_n 0.00960883f $X=11.58 $Y=0.465 $X2=0
+ $Y2=0
