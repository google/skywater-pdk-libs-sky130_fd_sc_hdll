* File: sky130_fd_sc_hdll__clkbuf_4.spice
* Created: Wed Sep  2 08:25:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkbuf_4.pex.spice"
.subckt sky130_fd_sc_hdll__clkbuf_4  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_27_47#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.1323 PD=0.75 PS=1.47 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.0693 PD=0.755 PS=0.75 NRD=15.708 NRS=14.28 M=1 R=2.8
+ SA=75000.7 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1001_d N_A_27_47#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.0693 PD=0.755 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_27_47#_M1005_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07875 AS=0.0693 PD=0.795 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1005_d N_A_27_47#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07875 AS=0.1239 PD=0.795 PS=1.43 NRD=12.852 NRS=1.428 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_27_47#_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.275 PD=1.35 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1003_d N_A_27_47#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=5.55556
+ SA=90000.7 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_27_47#_M1006_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.2
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1006_d N_A_27_47#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.7
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_27_47#_M1008_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.31 AS=0.15 PD=2.62 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_34 VNB 0 1.0084e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hdll__clkbuf_4.pxi.spice"
*
.ends
*
*
