* File: sky130_fd_sc_hdll__nor2_1.pxi.spice
* Created: Thu Aug 27 19:15:22 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR2_1%B N_B_c_28_n N_B_M1002_g N_B_c_29_n N_B_M1003_g B
+ PM_SKY130_FD_SC_HDLL__NOR2_1%B
x_PM_SKY130_FD_SC_HDLL__NOR2_1%A N_A_c_53_n N_A_M1001_g N_A_c_56_n N_A_M1000_g A
+ N_A_c_55_n PM_SKY130_FD_SC_HDLL__NOR2_1%A
x_PM_SKY130_FD_SC_HDLL__NOR2_1%Y N_Y_M1003_d N_Y_M1002_s N_Y_c_84_n N_Y_c_86_n
+ N_Y_c_79_n N_Y_c_82_n N_Y_c_80_n Y PM_SKY130_FD_SC_HDLL__NOR2_1%Y
x_PM_SKY130_FD_SC_HDLL__NOR2_1%VPWR N_VPWR_M1000_d N_VPWR_c_115_n N_VPWR_c_116_n
+ VPWR N_VPWR_c_117_n N_VPWR_c_114_n PM_SKY130_FD_SC_HDLL__NOR2_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR2_1%VGND N_VGND_M1003_s N_VGND_M1001_d N_VGND_c_132_n
+ N_VGND_c_133_n N_VGND_c_134_n N_VGND_c_135_n VGND N_VGND_c_136_n
+ N_VGND_c_137_n PM_SKY130_FD_SC_HDLL__NOR2_1%VGND
cc_1 VNB N_B_c_28_n 0.0435152f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_B_c_29_n 0.0218571f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB B 0.00935867f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_c_53_n 0.0218621f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB A 0.00879043f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_6 VNB N_A_c_55_n 0.043526f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_7 VNB N_Y_c_79_n 0.00749827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_Y_c_80_n 0.00378006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_VPWR_c_114_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_132_n 0.0101633f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_11 VNB N_VGND_c_133_n 0.0308989f $X=-0.19 $Y=-0.24 $X2=0.352 $Y2=1.16
cc_12 VNB N_VGND_c_134_n 0.0204605f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_13 VNB N_VGND_c_135_n 0.012224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_136_n 0.0190531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_137_n 0.128576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VPB N_B_c_28_n 0.0380561f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_17 VPB B 0.00121238f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_18 VPB N_A_c_56_n 0.0212438f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_19 VPB A 8.98319e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_20 VPB N_A_c_55_n 0.019432f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_21 VPB N_Y_c_79_n 0.00328455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_22 VPB N_Y_c_82_n 0.00741865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_23 VPB Y 0.0306411f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_115_n 0.018843f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_25 VPB N_VPWR_c_116_n 0.00664889f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_26 VPB N_VPWR_c_117_n 0.0346282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_114_n 0.0467325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 N_B_c_29_n N_A_c_53_n 0.0143924f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_29 N_B_c_28_n N_A_c_56_n 0.0498365f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_30 N_B_c_28_n N_A_c_55_n 0.0143924f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_31 N_B_c_28_n N_Y_c_84_n 0.0165114f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_32 B N_Y_c_84_n 6.64606e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_33 N_B_c_29_n N_Y_c_86_n 0.00710219f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_34 N_B_c_28_n N_Y_c_79_n 0.00192074f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_35 N_B_c_29_n N_Y_c_79_n 0.00903215f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_36 B N_Y_c_79_n 0.018812f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_37 N_B_c_28_n N_Y_c_82_n 0.00707562f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_38 B N_Y_c_82_n 0.0242077f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_39 N_B_c_29_n N_Y_c_80_n 0.0049136f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_40 N_B_c_28_n Y 0.0147792f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_41 N_B_c_28_n N_VPWR_c_117_n 0.00674013f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_42 N_B_c_28_n N_VPWR_c_114_n 0.0129574f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_43 N_B_c_28_n N_VGND_c_133_n 0.00597918f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_44 N_B_c_29_n N_VGND_c_133_n 0.00639232f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_45 B N_VGND_c_133_n 0.0188825f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_46 N_B_c_29_n N_VGND_c_136_n 0.00465454f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_47 N_B_c_29_n N_VGND_c_137_n 0.00880113f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_48 N_A_c_56_n N_Y_c_84_n 0.00179985f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_49 N_A_c_53_n N_Y_c_86_n 0.00517661f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_50 N_A_c_53_n N_Y_c_79_n 0.00837433f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_51 N_A_c_56_n N_Y_c_79_n 0.00191836f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_52 A N_Y_c_79_n 0.0132871f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_53 N_A_c_53_n N_Y_c_80_n 0.00365727f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A_c_56_n Y 0.00364275f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_55 N_A_c_56_n N_VPWR_c_116_n 0.0263505f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_56 A N_VPWR_c_116_n 0.0226811f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_57 N_A_c_55_n N_VPWR_c_116_n 0.00603357f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_58 N_A_c_56_n N_VPWR_c_117_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A_c_56_n N_VPWR_c_114_n 0.013896f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_c_53_n N_VGND_c_135_n 0.00493561f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_61 A N_VGND_c_135_n 0.0261605f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_62 N_A_c_55_n N_VGND_c_135_n 0.00789559f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_63 N_A_c_53_n N_VGND_c_136_n 0.00541359f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_64 N_A_c_53_n N_VGND_c_137_n 0.0108548f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_65 N_Y_c_84_n A_117_297# 0.00798242f $X=0.605 $Y=1.58 $X2=-0.19 $Y2=-0.24
cc_66 N_Y_c_84_n N_VPWR_c_116_n 0.00894521f $X=0.605 $Y=1.58 $X2=0 $Y2=0
cc_67 Y N_VPWR_c_117_n 0.0192237f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_68 N_Y_M1002_s N_VPWR_c_114_n 0.00218082f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_69 Y N_VPWR_c_114_n 0.012382f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_70 N_Y_c_86_n N_VGND_c_133_n 0.0489875f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_71 N_Y_c_86_n N_VGND_c_135_n 0.0249f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_72 N_Y_c_86_n N_VGND_c_136_n 0.0222708f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_73 N_Y_M1003_d N_VGND_c_137_n 0.00215201f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_74 N_Y_c_86_n N_VGND_c_137_n 0.0139062f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_75 A_117_297# N_VPWR_c_114_n 0.0123962f $X=0.585 $Y=1.485 $X2=0.15 $Y2=2.125
cc_76 N_VPWR_c_116_n N_VGND_c_135_n 0.00659342f $X=1.2 $Y=1.66 $X2=0 $Y2=0
