* File: sky130_fd_sc_hdll__a21oi_1.spice
* Created: Thu Aug 27 18:53:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21oi_1.pex.spice"
.subckt sky130_fd_sc_hdll__a21oi_1  VNB VPB B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_B1_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.20475 PD=0.98 PS=1.93 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.2
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1002 A_219_47# N_A1_M1002_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.65 AD=0.095875
+ AS=0.10725 PD=0.945 PS=0.98 NRD=17.076 NRS=9.228 M=1 R=4.33333 SA=75000.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_219_47# VNB NSHORT L=0.15 W=0.65 AD=0.20475
+ AS=0.095875 PD=1.93 PS=0.945 NRD=9.228 NRS=17.076 M=1 R=4.33333 SA=75001.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_121_297#_M1000_d N_B1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_121_297#_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1575 AS=0.15 PD=1.315 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1004 N_A_121_297#_M1004_d N_A2_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.1575 PD=2.55 PS=1.315 NRD=1.9503 NRS=4.9053 M=1 R=5.55556
+ SA=90001.2 SB=90000.2 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hdll__a21oi_1.pxi.spice"
*
.ends
*
*
