* File: sky130_fd_sc_hdll__a21bo_4.pxi.spice
* Created: Wed Sep  2 08:16:37 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21BO_4%B1_N N_B1_N_c_85_n N_B1_N_M1003_g N_B1_N_c_86_n
+ N_B1_N_M1013_g B1_N B1_N PM_SKY130_FD_SC_HDLL__A21BO_4%B1_N
x_PM_SKY130_FD_SC_HDLL__A21BO_4%A_209_21# N_A_209_21#_M1010_s
+ N_A_209_21#_M1011_d N_A_209_21#_M1005_s N_A_209_21#_c_116_n
+ N_A_209_21#_M1001_g N_A_209_21#_c_124_n N_A_209_21#_M1000_g
+ N_A_209_21#_c_117_n N_A_209_21#_M1004_g N_A_209_21#_c_125_n
+ N_A_209_21#_M1006_g N_A_209_21#_c_118_n N_A_209_21#_M1007_g
+ N_A_209_21#_c_126_n N_A_209_21#_M1012_g N_A_209_21#_c_119_n
+ N_A_209_21#_M1009_g N_A_209_21#_c_127_n N_A_209_21#_M1018_g
+ N_A_209_21#_c_195_p N_A_209_21#_c_120_n N_A_209_21#_c_138_p
+ N_A_209_21#_c_196_p N_A_209_21#_c_232_p N_A_209_21#_c_121_n
+ N_A_209_21#_c_142_p N_A_209_21#_c_122_n N_A_209_21#_c_173_p
+ N_A_209_21#_c_123_n PM_SKY130_FD_SC_HDLL__A21BO_4%A_209_21#
x_PM_SKY130_FD_SC_HDLL__A21BO_4%A_36_47# N_A_36_47#_M1013_s N_A_36_47#_M1003_s
+ N_A_36_47#_c_263_n N_A_36_47#_M1005_g N_A_36_47#_c_257_n N_A_36_47#_M1010_g
+ N_A_36_47#_c_264_n N_A_36_47#_M1019_g N_A_36_47#_c_258_n N_A_36_47#_M1016_g
+ N_A_36_47#_c_259_n N_A_36_47#_c_266_n N_A_36_47#_c_267_n N_A_36_47#_c_268_n
+ N_A_36_47#_c_260_n N_A_36_47#_c_261_n N_A_36_47#_c_270_n N_A_36_47#_c_262_n
+ PM_SKY130_FD_SC_HDLL__A21BO_4%A_36_47#
x_PM_SKY130_FD_SC_HDLL__A21BO_4%A2 N_A2_c_361_n N_A2_M1002_g N_A2_c_362_n
+ N_A2_M1015_g N_A2_c_363_n N_A2_M1017_g N_A2_c_364_n N_A2_M1008_g N_A2_c_365_n
+ N_A2_c_387_p N_A2_c_408_p N_A2_c_366_n A2 N_A2_c_368_n A2 N_A2_c_411_p
+ PM_SKY130_FD_SC_HDLL__A21BO_4%A2
x_PM_SKY130_FD_SC_HDLL__A21BO_4%A1 N_A1_c_442_n N_A1_M1011_g N_A1_c_445_n
+ N_A1_M1014_g N_A1_c_446_n N_A1_M1020_g N_A1_c_443_n N_A1_M1021_g A1
+ N_A1_c_444_n PM_SKY130_FD_SC_HDLL__A21BO_4%A1
x_PM_SKY130_FD_SC_HDLL__A21BO_4%VPWR N_VPWR_M1003_d N_VPWR_M1006_s
+ N_VPWR_M1018_s N_VPWR_M1002_d N_VPWR_M1020_d N_VPWR_c_490_n N_VPWR_c_491_n
+ N_VPWR_c_492_n N_VPWR_c_493_n VPWR N_VPWR_c_494_n N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_489_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n
+ N_VPWR_c_501_n PM_SKY130_FD_SC_HDLL__A21BO_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A21BO_4%X N_X_M1001_d N_X_M1007_d N_X_M1000_d
+ N_X_M1012_d N_X_c_593_n N_X_c_599_n N_X_c_589_n X N_X_c_614_n X
+ PM_SKY130_FD_SC_HDLL__A21BO_4%X
x_PM_SKY130_FD_SC_HDLL__A21BO_4%A_647_297# N_A_647_297#_M1005_d
+ N_A_647_297#_M1019_d N_A_647_297#_M1014_s N_A_647_297#_M1008_s
+ N_A_647_297#_c_638_n N_A_647_297#_c_640_n N_A_647_297#_c_675_n
+ N_A_647_297#_c_635_n N_A_647_297#_c_636_n N_A_647_297#_c_637_n
+ N_A_647_297#_c_666_n PM_SKY130_FD_SC_HDLL__A21BO_4%A_647_297#
x_PM_SKY130_FD_SC_HDLL__A21BO_4%VGND N_VGND_M1013_d N_VGND_M1004_s
+ N_VGND_M1009_s N_VGND_M1016_d N_VGND_M1017_s N_VGND_c_690_n N_VGND_c_691_n
+ N_VGND_c_692_n N_VGND_c_693_n N_VGND_c_694_n VGND N_VGND_c_695_n
+ N_VGND_c_696_n N_VGND_c_697_n N_VGND_c_698_n N_VGND_c_699_n N_VGND_c_700_n
+ N_VGND_c_701_n PM_SKY130_FD_SC_HDLL__A21BO_4%VGND
cc_1 VNB N_B1_N_c_85_n 0.0303545f $X=-0.19 $Y=-0.24 $X2=0.665 $Y2=1.41
cc_2 VNB N_B1_N_c_86_n 0.0193875f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=0.995
cc_3 VNB B1_N 0.00539178f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.105
cc_4 VNB N_A_209_21#_c_116_n 0.0161856f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_5 VNB N_A_209_21#_c_117_n 0.0164758f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_209_21#_c_118_n 0.0169445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_209_21#_c_119_n 0.0199397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_209_21#_c_120_n 0.00270467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_209_21#_c_121_n 0.00200356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_209_21#_c_122_n 0.0127551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_209_21#_c_123_n 0.0867889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_36_47#_c_257_n 0.0203971f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_13 VNB N_A_36_47#_c_258_n 0.0174864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_36_47#_c_259_n 0.0227203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_36_47#_c_260_n 0.00563558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_36_47#_c_261_n 0.0244955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_36_47#_c_262_n 0.0505713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_361_n 0.0214769f $X=-0.19 $Y=-0.24 $X2=0.665 $Y2=1.41
cc_19 VNB N_A2_c_362_n 0.016891f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=0.995
cc_20 VNB N_A2_c_363_n 0.0222254f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.105
cc_21 VNB N_A2_c_364_n 0.0315997f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_22 VNB N_A2_c_365_n 4.45289e-19 $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.19
cc_23 VNB N_A2_c_366_n 0.0106746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB A2 0.0103411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A2_c_368_n 0.00551268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A1_c_442_n 0.0167836f $X=-0.19 $Y=-0.24 $X2=0.665 $Y2=1.41
cc_27 VNB N_A1_c_443_n 0.0171772f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_28 VNB N_A1_c_444_n 0.0378066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_489_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_690_n 0.00508428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_691_n 0.0106171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_692_n 0.0330065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_693_n 0.00547506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_694_n 0.0136657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_695_n 0.0174728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_696_n 0.0451341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_697_n 0.0245781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_698_n 0.0191309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_699_n 0.0223596f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_700_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_701_n 0.314954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VPB N_B1_N_c_85_n 0.029797f $X=-0.19 $Y=1.305 $X2=0.665 $Y2=1.41
cc_43 VPB B1_N 0.00284034f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.105
cc_44 VPB N_A_209_21#_c_124_n 0.0156286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_209_21#_c_125_n 0.0156811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_209_21#_c_126_n 0.0162804f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_209_21#_c_127_n 0.0182602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_209_21#_c_121_n 0.00239987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_209_21#_c_122_n 0.00105623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_209_21#_c_123_n 0.0525047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_36_47#_c_263_n 0.0196006f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.105
cc_52 VPB N_A_36_47#_c_264_n 0.0164022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_36_47#_c_259_n 0.0241587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_36_47#_c_266_n 0.00348512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_36_47#_c_267_n 0.00584684f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_36_47#_c_268_n 0.0126124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_36_47#_c_260_n 0.00142271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_36_47#_c_270_n 0.0323602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_36_47#_c_262_n 0.0307875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A2_c_361_n 0.0255632f $X=-0.19 $Y=1.305 $X2=0.665 $Y2=1.41
cc_61 VPB N_A2_c_364_n 0.032768f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_62 VPB N_A2_c_365_n 0.0015339f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.19
cc_63 VPB A2 0.00168688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A1_c_445_n 0.0162041f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=0.995
cc_65 VPB N_A1_c_446_n 0.0159226f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.105
cc_66 VPB A1 0.00282525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A1_c_444_n 0.0203032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_490_n 0.00538384f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_491_n 0.01367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_492_n 0.0115737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_493_n 0.013534f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_494_n 0.0386589f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_495_n 0.013126f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_496_n 0.0169235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_489_n 0.0535609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_498_n 0.00547506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_499_n 0.0183862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_500_n 0.00547137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_501_n 0.00547137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB X 5.07614e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_647_297#_c_635_n 0.00333169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_647_297#_c_636_n 0.00767904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_647_297#_c_637_n 0.0210132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 N_B1_N_c_86_n N_A_209_21#_c_116_n 0.0246057f $X=0.69 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B1_N_c_85_n N_A_209_21#_c_124_n 0.037019f $X=0.665 $Y=1.41 $X2=0 $Y2=0
cc_86 B1_N N_A_209_21#_c_124_n 8.06251e-19 $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_87 N_B1_N_c_85_n N_A_209_21#_c_123_n 0.0237476f $X=0.665 $Y=1.41 $X2=0 $Y2=0
cc_88 B1_N N_A_209_21#_c_123_n 0.00262577f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_89 B1_N N_A_36_47#_M1003_s 0.00204566f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B1_N_c_85_n N_A_36_47#_c_259_n 0.00813204f $X=0.665 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B1_N_c_86_n N_A_36_47#_c_259_n 0.00311524f $X=0.69 $Y=0.995 $X2=0 $Y2=0
cc_92 B1_N N_A_36_47#_c_259_n 0.0496417f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B1_N_c_85_n N_A_36_47#_c_266_n 0.0118287f $X=0.665 $Y=1.41 $X2=0 $Y2=0
cc_94 B1_N N_A_36_47#_c_266_n 0.0103074f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B1_N_c_85_n N_A_36_47#_c_261_n 2.12172e-19 $X=0.665 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B1_N_c_86_n N_A_36_47#_c_261_n 0.016918f $X=0.69 $Y=0.995 $X2=0 $Y2=0
cc_97 B1_N N_A_36_47#_c_261_n 0.00346284f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_98 B1_N N_A_36_47#_c_270_n 0.00427105f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_99 B1_N N_VPWR_M1003_d 0.00183947f $X=0.575 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_100 N_B1_N_c_85_n N_VPWR_c_489_n 0.00485239f $X=0.665 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B1_N_c_85_n N_VPWR_c_498_n 0.0104595f $X=0.665 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B1_N_c_85_n N_VPWR_c_499_n 0.0032362f $X=0.665 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B1_N_c_86_n N_X_c_589_n 6.43894e-19 $X=0.69 $Y=0.995 $X2=0 $Y2=0
cc_104 N_B1_N_c_85_n X 8.8441e-19 $X=0.665 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B1_N_c_86_n X 0.00115679f $X=0.69 $Y=0.995 $X2=0 $Y2=0
cc_106 B1_N X 0.0390144f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_107 N_B1_N_c_86_n N_VGND_c_697_n 0.0149142f $X=0.69 $Y=0.995 $X2=0 $Y2=0
cc_108 B1_N N_VGND_c_697_n 0.00447855f $X=0.575 $Y=1.105 $X2=0 $Y2=0
cc_109 N_B1_N_c_86_n N_VGND_c_701_n 0.00582584f $X=0.69 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_209_21#_c_121_n N_A_36_47#_c_263_n 0.00270839f $X=3.83 $Y=1.62 $X2=0
+ $Y2=0
cc_111 N_A_209_21#_c_120_n N_A_36_47#_c_257_n 0.00497407f $X=2.945 $Y=0.995
+ $X2=0 $Y2=0
cc_112 N_A_209_21#_c_138_p N_A_36_47#_c_257_n 0.0162401f $X=3.745 $Y=0.7 $X2=0
+ $Y2=0
cc_113 N_A_209_21#_c_121_n N_A_36_47#_c_257_n 0.0026752f $X=3.83 $Y=1.62 $X2=0
+ $Y2=0
cc_114 N_A_209_21#_c_121_n N_A_36_47#_c_264_n 0.00222706f $X=3.83 $Y=1.62 $X2=0
+ $Y2=0
cc_115 N_A_209_21#_c_121_n N_A_36_47#_c_258_n 0.00335184f $X=3.83 $Y=1.62 $X2=0
+ $Y2=0
cc_116 N_A_209_21#_c_142_p N_A_36_47#_c_258_n 0.014874f $X=5.105 $Y=0.755 $X2=0
+ $Y2=0
cc_117 N_A_209_21#_c_124_n N_A_36_47#_c_266_n 0.0133781f $X=1.145 $Y=1.41 $X2=0
+ $Y2=0
cc_118 N_A_209_21#_c_125_n N_A_36_47#_c_266_n 0.0128321f $X=1.625 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_209_21#_c_126_n N_A_36_47#_c_266_n 0.0134306f $X=2.105 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_A_209_21#_c_127_n N_A_36_47#_c_266_n 0.0157717f $X=2.585 $Y=1.41 $X2=0
+ $Y2=0
cc_121 N_A_209_21#_c_122_n N_A_36_47#_c_266_n 0.00346564f $X=2.615 $Y=1.16 $X2=0
+ $Y2=0
cc_122 N_A_209_21#_c_123_n N_A_36_47#_c_266_n 0.00207988f $X=2.585 $Y=1.202
+ $X2=0 $Y2=0
cc_123 N_A_209_21#_c_127_n N_A_36_47#_c_267_n 0.0111131f $X=2.585 $Y=1.41 $X2=0
+ $Y2=0
cc_124 N_A_209_21#_c_121_n N_A_36_47#_c_267_n 0.00469861f $X=3.83 $Y=1.62 $X2=0
+ $Y2=0
cc_125 N_A_209_21#_c_127_n N_A_36_47#_c_268_n 0.00428396f $X=2.585 $Y=1.41 $X2=0
+ $Y2=0
cc_126 N_A_209_21#_c_138_p N_A_36_47#_c_268_n 0.00576396f $X=3.745 $Y=0.7 $X2=0
+ $Y2=0
cc_127 N_A_209_21#_c_121_n N_A_36_47#_c_268_n 0.0108546f $X=3.83 $Y=1.62 $X2=0
+ $Y2=0
cc_128 N_A_209_21#_c_122_n N_A_36_47#_c_268_n 0.00915628f $X=2.615 $Y=1.16 $X2=0
+ $Y2=0
cc_129 N_A_209_21#_c_123_n N_A_36_47#_c_268_n 0.00208042f $X=2.585 $Y=1.202
+ $X2=0 $Y2=0
cc_130 N_A_209_21#_c_138_p N_A_36_47#_c_260_n 0.0187942f $X=3.745 $Y=0.7 $X2=0
+ $Y2=0
cc_131 N_A_209_21#_c_121_n N_A_36_47#_c_260_n 0.0209295f $X=3.83 $Y=1.62 $X2=0
+ $Y2=0
cc_132 N_A_209_21#_c_122_n N_A_36_47#_c_260_n 0.0212365f $X=2.615 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_A_209_21#_c_123_n N_A_36_47#_c_260_n 0.00250931f $X=2.585 $Y=1.202
+ $X2=0 $Y2=0
cc_134 N_A_209_21#_c_138_p N_A_36_47#_c_262_n 0.00138581f $X=3.745 $Y=0.7 $X2=0
+ $Y2=0
cc_135 N_A_209_21#_c_121_n N_A_36_47#_c_262_n 0.0246205f $X=3.83 $Y=1.62 $X2=0
+ $Y2=0
cc_136 N_A_209_21#_c_142_p N_A_36_47#_c_262_n 3.64185e-19 $X=5.105 $Y=0.755
+ $X2=0 $Y2=0
cc_137 N_A_209_21#_c_122_n N_A_36_47#_c_262_n 8.52775e-19 $X=2.615 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_209_21#_c_123_n N_A_36_47#_c_262_n 0.00654167f $X=2.585 $Y=1.202
+ $X2=0 $Y2=0
cc_139 N_A_209_21#_c_121_n N_A2_c_361_n 4.32833e-19 $X=3.83 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_140 N_A_209_21#_c_142_p N_A2_c_361_n 0.00362527f $X=5.105 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A_209_21#_c_142_p N_A2_c_362_n 0.0120398f $X=5.105 $Y=0.755 $X2=0 $Y2=0
cc_142 N_A_209_21#_c_121_n N_A2_c_365_n 0.00424417f $X=3.83 $Y=1.62 $X2=0 $Y2=0
cc_143 N_A_209_21#_c_121_n N_A2_c_368_n 0.0102371f $X=3.83 $Y=1.62 $X2=0 $Y2=0
cc_144 N_A_209_21#_c_142_p N_A2_c_368_n 0.0283014f $X=5.105 $Y=0.755 $X2=0 $Y2=0
cc_145 N_A_209_21#_c_142_p N_A1_c_442_n 0.0117599f $X=5.105 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_146 N_A_209_21#_c_142_p A1 0.00870954f $X=5.105 $Y=0.755 $X2=0 $Y2=0
cc_147 N_A_209_21#_c_173_p A1 0.020986f $X=5.24 $Y=0.57 $X2=0 $Y2=0
cc_148 N_A_209_21#_c_173_p N_A1_c_444_n 0.00444199f $X=5.24 $Y=0.57 $X2=0 $Y2=0
cc_149 N_A_209_21#_c_124_n N_VPWR_c_490_n 0.00111962f $X=1.145 $Y=1.41 $X2=0
+ $Y2=0
cc_150 N_A_209_21#_c_125_n N_VPWR_c_490_n 0.0105269f $X=1.625 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_A_209_21#_c_126_n N_VPWR_c_490_n 0.00768958f $X=2.105 $Y=1.41 $X2=0
+ $Y2=0
cc_152 N_A_209_21#_c_127_n N_VPWR_c_490_n 0.00100315f $X=2.585 $Y=1.41 $X2=0
+ $Y2=0
cc_153 N_A_209_21#_c_124_n N_VPWR_c_491_n 0.00464324f $X=1.145 $Y=1.41 $X2=0
+ $Y2=0
cc_154 N_A_209_21#_c_125_n N_VPWR_c_491_n 0.0032362f $X=1.625 $Y=1.41 $X2=0
+ $Y2=0
cc_155 N_A_209_21#_c_126_n N_VPWR_c_492_n 0.00112904f $X=2.105 $Y=1.41 $X2=0
+ $Y2=0
cc_156 N_A_209_21#_c_127_n N_VPWR_c_492_n 0.011771f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_209_21#_c_126_n N_VPWR_c_493_n 0.00464324f $X=2.105 $Y=1.41 $X2=0
+ $Y2=0
cc_158 N_A_209_21#_c_127_n N_VPWR_c_493_n 0.00309549f $X=2.585 $Y=1.41 $X2=0
+ $Y2=0
cc_159 N_A_209_21#_M1005_s N_VPWR_c_489_n 0.00241663f $X=3.685 $Y=1.485 $X2=0
+ $Y2=0
cc_160 N_A_209_21#_c_124_n N_VPWR_c_489_n 0.00529844f $X=1.145 $Y=1.41 $X2=0
+ $Y2=0
cc_161 N_A_209_21#_c_125_n N_VPWR_c_489_n 0.00388795f $X=1.625 $Y=1.41 $X2=0
+ $Y2=0
cc_162 N_A_209_21#_c_126_n N_VPWR_c_489_n 0.00529844f $X=2.105 $Y=1.41 $X2=0
+ $Y2=0
cc_163 N_A_209_21#_c_127_n N_VPWR_c_489_n 0.0037469f $X=2.585 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_209_21#_c_124_n N_VPWR_c_498_n 0.00768031f $X=1.145 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_A_209_21#_c_125_n N_VPWR_c_498_n 0.00100586f $X=1.625 $Y=1.41 $X2=0
+ $Y2=0
cc_166 N_A_209_21#_c_117_n N_X_c_593_n 0.0130941f $X=1.6 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_209_21#_c_118_n N_X_c_593_n 0.0100176f $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_209_21#_c_119_n N_X_c_593_n 0.00347369f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_209_21#_c_195_p N_X_c_593_n 0.0437179f $X=2.585 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_209_21#_c_196_p N_X_c_593_n 0.00839667f $X=3.03 $Y=0.7 $X2=0 $Y2=0
cc_171 N_A_209_21#_c_123_n N_X_c_593_n 0.00655084f $X=2.585 $Y=1.202 $X2=0 $Y2=0
cc_172 N_A_209_21#_c_125_n N_X_c_599_n 0.0148235f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_209_21#_c_126_n N_X_c_599_n 0.0105501f $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_209_21#_c_127_n N_X_c_599_n 0.00597541f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_209_21#_c_195_p N_X_c_599_n 0.0384425f $X=2.585 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_209_21#_c_123_n N_X_c_599_n 0.0121227f $X=2.585 $Y=1.202 $X2=0 $Y2=0
cc_177 N_A_209_21#_c_116_n N_X_c_589_n 0.00736308f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_209_21#_c_117_n N_X_c_589_n 5.35717e-19 $X=1.6 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_209_21#_c_116_n X 0.00717333f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_209_21#_c_124_n X 0.00463973f $X=1.145 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_209_21#_c_117_n X 0.00545196f $X=1.6 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_209_21#_c_125_n X 0.00429671f $X=1.625 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_209_21#_c_118_n X 9.7202e-19 $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_209_21#_c_126_n X 8.22614e-19 $X=2.105 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_209_21#_c_195_p X 0.0269532f $X=2.585 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_209_21#_c_123_n X 0.037467f $X=2.585 $Y=1.202 $X2=0 $Y2=0
cc_187 N_A_209_21#_c_124_n N_X_c_614_n 0.00604641f $X=1.145 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_209_21#_c_127_n N_A_647_297#_c_638_n 0.00262841f $X=2.585 $Y=1.41
+ $X2=0 $Y2=0
cc_189 N_A_209_21#_c_121_n N_A_647_297#_c_638_n 0.00525856f $X=3.83 $Y=1.62
+ $X2=0 $Y2=0
cc_190 N_A_209_21#_M1005_s N_A_647_297#_c_640_n 0.00458721f $X=3.685 $Y=1.485
+ $X2=0 $Y2=0
cc_191 N_A_209_21#_c_121_n N_A_647_297#_c_640_n 0.00719556f $X=3.83 $Y=1.62
+ $X2=0 $Y2=0
cc_192 N_A_209_21#_c_121_n N_A_647_297#_c_635_n 0.00989862f $X=3.83 $Y=1.62
+ $X2=0 $Y2=0
cc_193 N_A_209_21#_c_142_p N_A_647_297#_c_635_n 0.00440519f $X=5.105 $Y=0.755
+ $X2=0 $Y2=0
cc_194 N_A_209_21#_c_120_n N_VGND_M1009_s 0.0031999f $X=2.945 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_209_21#_c_138_p N_VGND_M1009_s 0.014076f $X=3.745 $Y=0.7 $X2=0 $Y2=0
cc_196 N_A_209_21#_c_196_p N_VGND_M1009_s 0.0054155f $X=3.03 $Y=0.7 $X2=0 $Y2=0
cc_197 N_A_209_21#_c_142_p N_VGND_M1016_d 0.00639913f $X=5.105 $Y=0.755 $X2=0
+ $Y2=0
cc_198 N_A_209_21#_c_142_p N_VGND_c_690_n 0.0147553f $X=5.105 $Y=0.755 $X2=0
+ $Y2=0
cc_199 N_A_209_21#_c_116_n N_VGND_c_693_n 0.00106058f $X=1.12 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_209_21#_c_117_n N_VGND_c_693_n 0.00819243f $X=1.6 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_209_21#_c_118_n N_VGND_c_693_n 0.00939017f $X=2.08 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_209_21#_c_119_n N_VGND_c_693_n 0.00196005f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_209_21#_c_116_n N_VGND_c_694_n 0.00351635f $X=1.12 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_209_21#_c_117_n N_VGND_c_694_n 0.00351745f $X=1.6 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_209_21#_c_138_p N_VGND_c_695_n 0.00348385f $X=3.745 $Y=0.7 $X2=0
+ $Y2=0
cc_206 N_A_209_21#_c_232_p N_VGND_c_695_n 0.0116048f $X=3.83 $Y=0.42 $X2=0 $Y2=0
cc_207 N_A_209_21#_c_142_p N_VGND_c_695_n 0.00353953f $X=5.105 $Y=0.755 $X2=0
+ $Y2=0
cc_208 N_A_209_21#_c_142_p N_VGND_c_696_n 0.00804207f $X=5.105 $Y=0.755 $X2=0
+ $Y2=0
cc_209 N_A_209_21#_c_173_p N_VGND_c_696_n 0.00922285f $X=5.24 $Y=0.57 $X2=0
+ $Y2=0
cc_210 N_A_209_21#_c_116_n N_VGND_c_697_n 0.00787709f $X=1.12 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_209_21#_c_117_n N_VGND_c_697_n 0.00106105f $X=1.6 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_A_209_21#_c_118_n N_VGND_c_698_n 0.0035176f $X=2.08 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_209_21#_c_119_n N_VGND_c_698_n 0.00558173f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A_209_21#_c_119_n N_VGND_c_699_n 0.013604f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_209_21#_c_138_p N_VGND_c_699_n 0.0345011f $X=3.745 $Y=0.7 $X2=0 $Y2=0
cc_216 N_A_209_21#_c_196_p N_VGND_c_699_n 0.01398f $X=3.03 $Y=0.7 $X2=0 $Y2=0
cc_217 N_A_209_21#_c_122_n N_VGND_c_699_n 0.00414494f $X=2.615 $Y=1.16 $X2=0
+ $Y2=0
cc_218 N_A_209_21#_c_123_n N_VGND_c_699_n 4.02743e-19 $X=2.585 $Y=1.202 $X2=0
+ $Y2=0
cc_219 N_A_209_21#_M1010_s N_VGND_c_701_n 0.00311376f $X=3.695 $Y=0.235 $X2=0
+ $Y2=0
cc_220 N_A_209_21#_M1011_d N_VGND_c_701_n 0.00481352f $X=5.055 $Y=0.235 $X2=0
+ $Y2=0
cc_221 N_A_209_21#_c_116_n N_VGND_c_701_n 0.00424416f $X=1.12 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_209_21#_c_117_n N_VGND_c_701_n 0.00424592f $X=1.6 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_209_21#_c_118_n N_VGND_c_701_n 0.00424616f $X=2.08 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_209_21#_c_119_n N_VGND_c_701_n 0.011515f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_209_21#_c_138_p N_VGND_c_701_n 0.00826721f $X=3.745 $Y=0.7 $X2=0
+ $Y2=0
cc_226 N_A_209_21#_c_196_p N_VGND_c_701_n 8.76362e-19 $X=3.03 $Y=0.7 $X2=0 $Y2=0
cc_227 N_A_209_21#_c_232_p N_VGND_c_701_n 0.00646998f $X=3.83 $Y=0.42 $X2=0
+ $Y2=0
cc_228 N_A_209_21#_c_142_p N_VGND_c_701_n 0.0228608f $X=5.105 $Y=0.755 $X2=0
+ $Y2=0
cc_229 N_A_209_21#_c_173_p N_VGND_c_701_n 0.00967148f $X=5.24 $Y=0.57 $X2=0
+ $Y2=0
cc_230 N_A_209_21#_c_142_p A_1115_47# 0.00492452f $X=5.105 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_231 N_A_36_47#_c_264_n N_A2_c_361_n 0.0207407f $X=4.065 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_232 N_A_36_47#_c_262_n N_A2_c_361_n 0.0260722f $X=4.065 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_233 N_A_36_47#_c_258_n N_A2_c_362_n 0.0201748f $X=4.09 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_36_47#_c_262_n N_A2_c_365_n 4.38741e-19 $X=4.065 $Y=1.202 $X2=0 $Y2=0
cc_235 N_A_36_47#_c_262_n N_A2_c_368_n 0.00256018f $X=4.065 $Y=1.202 $X2=0 $Y2=0
cc_236 N_A_36_47#_c_266_n N_VPWR_M1003_d 0.00806509f $X=2.92 $Y=2.02 $X2=-0.19
+ $Y2=-0.24
cc_237 N_A_36_47#_c_266_n N_VPWR_M1006_s 0.00371167f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_238 N_A_36_47#_c_266_n N_VPWR_M1018_s 0.0090856f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_239 N_A_36_47#_c_267_n N_VPWR_M1018_s 0.00600737f $X=3.005 $Y=1.935 $X2=0
+ $Y2=0
cc_240 N_A_36_47#_c_268_n N_VPWR_M1018_s 7.73555e-19 $X=3.37 $Y=1.355 $X2=0
+ $Y2=0
cc_241 N_A_36_47#_c_266_n N_VPWR_c_490_n 0.019553f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_242 N_A_36_47#_c_266_n N_VPWR_c_491_n 0.00938267f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_243 N_A_36_47#_c_263_n N_VPWR_c_492_n 0.00450246f $X=3.595 $Y=1.41 $X2=0
+ $Y2=0
cc_244 N_A_36_47#_c_266_n N_VPWR_c_492_n 0.0248644f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_245 N_A_36_47#_c_266_n N_VPWR_c_493_n 0.00929692f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_246 N_A_36_47#_c_263_n N_VPWR_c_494_n 0.00450022f $X=3.595 $Y=1.41 $X2=0
+ $Y2=0
cc_247 N_A_36_47#_c_264_n N_VPWR_c_494_n 0.00450022f $X=4.065 $Y=1.41 $X2=0
+ $Y2=0
cc_248 N_A_36_47#_c_266_n N_VPWR_c_494_n 0.00209217f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_249 N_A_36_47#_M1003_s N_VPWR_c_489_n 0.00239749f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_250 N_A_36_47#_c_263_n N_VPWR_c_489_n 0.0074987f $X=3.595 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_36_47#_c_264_n N_VPWR_c_489_n 0.00619321f $X=4.065 $Y=1.41 $X2=0
+ $Y2=0
cc_252 N_A_36_47#_c_266_n N_VPWR_c_489_n 0.0427385f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_253 N_A_36_47#_c_270_n N_VPWR_c_489_n 0.0164007f $X=0.32 $Y=2.02 $X2=0 $Y2=0
cc_254 N_A_36_47#_c_266_n N_VPWR_c_498_n 0.019553f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_255 N_A_36_47#_c_266_n N_VPWR_c_499_n 0.00237813f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_256 N_A_36_47#_c_270_n N_VPWR_c_499_n 0.0292923f $X=0.32 $Y=2.02 $X2=0 $Y2=0
cc_257 N_A_36_47#_c_264_n N_VPWR_c_500_n 0.00158396f $X=4.065 $Y=1.41 $X2=0
+ $Y2=0
cc_258 N_A_36_47#_c_266_n N_X_M1000_d 0.00498114f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_259 N_A_36_47#_c_266_n N_X_M1012_d 0.00498533f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_260 N_A_36_47#_c_266_n N_X_c_599_n 0.0567413f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_261 N_A_36_47#_c_267_n N_X_c_599_n 0.00772309f $X=3.005 $Y=1.935 $X2=0 $Y2=0
cc_262 N_A_36_47#_c_261_n N_X_c_589_n 0.00573f $X=0.345 $Y=0.36 $X2=0 $Y2=0
cc_263 N_A_36_47#_c_261_n X 0.00179152f $X=0.345 $Y=0.36 $X2=0 $Y2=0
cc_264 N_A_36_47#_c_266_n N_X_c_614_n 0.0290987f $X=2.92 $Y=2.02 $X2=0 $Y2=0
cc_265 N_A_36_47#_c_268_n N_A_647_297#_M1005_d 0.00343438f $X=3.37 $Y=1.355
+ $X2=-0.19 $Y2=-0.24
cc_266 N_A_36_47#_c_266_n N_A_647_297#_c_638_n 0.0132908f $X=2.92 $Y=2.02 $X2=0
+ $Y2=0
cc_267 N_A_36_47#_c_267_n N_A_647_297#_c_638_n 0.0166633f $X=3.005 $Y=1.935
+ $X2=0 $Y2=0
cc_268 N_A_36_47#_c_268_n N_A_647_297#_c_638_n 0.0136764f $X=3.37 $Y=1.355 $X2=0
+ $Y2=0
cc_269 N_A_36_47#_c_263_n N_A_647_297#_c_640_n 0.0149823f $X=3.595 $Y=1.41 $X2=0
+ $Y2=0
cc_270 N_A_36_47#_c_264_n N_A_647_297#_c_640_n 0.0156264f $X=4.065 $Y=1.41 $X2=0
+ $Y2=0
cc_271 N_A_36_47#_c_264_n N_A_647_297#_c_635_n 6.1325e-19 $X=4.065 $Y=1.41 $X2=0
+ $Y2=0
cc_272 N_A_36_47#_c_258_n N_VGND_c_690_n 0.0018666f $X=4.09 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_36_47#_c_257_n N_VGND_c_695_n 0.00422112f $X=3.62 $Y=0.995 $X2=0
+ $Y2=0
cc_274 N_A_36_47#_c_258_n N_VGND_c_695_n 0.00430182f $X=4.09 $Y=0.995 $X2=0
+ $Y2=0
cc_275 N_A_36_47#_c_261_n N_VGND_c_697_n 0.0434499f $X=0.345 $Y=0.36 $X2=0 $Y2=0
cc_276 N_A_36_47#_c_257_n N_VGND_c_699_n 0.00749714f $X=3.62 $Y=0.995 $X2=0
+ $Y2=0
cc_277 N_A_36_47#_M1013_s N_VGND_c_701_n 0.00724027f $X=0.18 $Y=0.235 $X2=0
+ $Y2=0
cc_278 N_A_36_47#_c_257_n N_VGND_c_701_n 0.00713982f $X=3.62 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_A_36_47#_c_258_n N_VGND_c_701_n 0.00601154f $X=4.09 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_36_47#_c_261_n N_VGND_c_701_n 0.0154887f $X=0.345 $Y=0.36 $X2=0 $Y2=0
cc_281 N_A2_c_362_n N_A1_c_442_n 0.0516638f $X=4.6 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_282 N_A2_c_361_n N_A1_c_445_n 0.0380956f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_283 N_A2_c_365_n N_A1_c_445_n 0.00429595f $X=4.677 $Y=1.595 $X2=0 $Y2=0
cc_284 N_A2_c_387_p N_A1_c_445_n 0.0135879f $X=5.63 $Y=1.68 $X2=0 $Y2=0
cc_285 N_A2_c_364_n N_A1_c_446_n 0.0383045f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_286 N_A2_c_387_p N_A1_c_446_n 0.0173644f $X=5.63 $Y=1.68 $X2=0 $Y2=0
cc_287 A2 N_A1_c_446_n 0.00465095f $X=5.69 $Y=1.445 $X2=0 $Y2=0
cc_288 N_A2_c_363_n N_A1_c_443_n 0.0308723f $X=5.92 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A2_c_361_n A1 3.26318e-19 $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_290 N_A2_c_364_n A1 4.20876e-19 $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_291 N_A2_c_365_n A1 0.0065944f $X=4.677 $Y=1.595 $X2=0 $Y2=0
cc_292 N_A2_c_387_p A1 0.0218511f $X=5.63 $Y=1.68 $X2=0 $Y2=0
cc_293 N_A2_c_366_n A1 0.0147415f $X=5.86 $Y=1.172 $X2=0 $Y2=0
cc_294 N_A2_c_368_n A1 0.0218795f $X=4.677 $Y=1.142 $X2=0 $Y2=0
cc_295 A2 A1 0.00397009f $X=5.69 $Y=1.445 $X2=0 $Y2=0
cc_296 N_A2_c_361_n N_A1_c_444_n 0.0254638f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_297 N_A2_c_364_n N_A1_c_444_n 0.0308723f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_298 N_A2_c_365_n N_A1_c_444_n 0.00174922f $X=4.677 $Y=1.595 $X2=0 $Y2=0
cc_299 N_A2_c_387_p N_A1_c_444_n 0.00140717f $X=5.63 $Y=1.68 $X2=0 $Y2=0
cc_300 N_A2_c_366_n N_A1_c_444_n 0.0025976f $X=5.86 $Y=1.172 $X2=0 $Y2=0
cc_301 N_A2_c_368_n N_A1_c_444_n 0.00186335f $X=4.677 $Y=1.142 $X2=0 $Y2=0
cc_302 A2 N_A1_c_444_n 0.00193627f $X=5.69 $Y=1.445 $X2=0 $Y2=0
cc_303 N_A2_c_365_n N_VPWR_M1002_d 0.00127321f $X=4.677 $Y=1.595 $X2=0 $Y2=0
cc_304 N_A2_c_387_p N_VPWR_M1002_d 0.00327038f $X=5.63 $Y=1.68 $X2=0 $Y2=0
cc_305 N_A2_c_408_p N_VPWR_M1002_d 0.00117519f $X=4.79 $Y=1.68 $X2=0 $Y2=0
cc_306 N_A2_c_387_p N_VPWR_M1020_d 3.41682e-19 $X=5.63 $Y=1.68 $X2=0 $Y2=0
cc_307 A2 N_VPWR_M1020_d 0.0012454f $X=5.69 $Y=1.445 $X2=0 $Y2=0
cc_308 N_A2_c_411_p N_VPWR_M1020_d 0.00185505f $X=5.745 $Y=1.595 $X2=0 $Y2=0
cc_309 N_A2_c_361_n N_VPWR_c_494_n 0.00309549f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A2_c_364_n N_VPWR_c_496_n 0.00450253f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A2_c_361_n N_VPWR_c_489_n 0.00374672f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_312 N_A2_c_364_n N_VPWR_c_489_n 0.00607752f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_313 N_A2_c_361_n N_VPWR_c_500_n 0.0109362f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A2_c_364_n N_VPWR_c_501_n 0.0140442f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A2_c_387_p N_A_647_297#_M1014_s 0.00361554f $X=5.63 $Y=1.68 $X2=0 $Y2=0
cc_316 N_A2_c_361_n N_A_647_297#_c_635_n 0.00495235f $X=4.535 $Y=1.41 $X2=0
+ $Y2=0
cc_317 N_A2_c_365_n N_A_647_297#_c_635_n 0.0103551f $X=4.677 $Y=1.595 $X2=0
+ $Y2=0
cc_318 N_A2_c_408_p N_A_647_297#_c_635_n 0.0128305f $X=4.79 $Y=1.68 $X2=0 $Y2=0
cc_319 N_A2_c_368_n N_A_647_297#_c_635_n 0.00336061f $X=4.677 $Y=1.142 $X2=0
+ $Y2=0
cc_320 N_A2_c_361_n N_A_647_297#_c_636_n 0.0132067f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A2_c_364_n N_A_647_297#_c_636_n 0.013531f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A2_c_387_p N_A_647_297#_c_636_n 0.0425641f $X=5.63 $Y=1.68 $X2=0 $Y2=0
cc_323 N_A2_c_408_p N_A_647_297#_c_636_n 0.0129215f $X=4.79 $Y=1.68 $X2=0 $Y2=0
cc_324 A2 N_A_647_297#_c_636_n 0.00462982f $X=5.925 $Y=1.2 $X2=0 $Y2=0
cc_325 N_A2_c_368_n N_A_647_297#_c_636_n 0.00347175f $X=4.677 $Y=1.142 $X2=0
+ $Y2=0
cc_326 N_A2_c_411_p N_A_647_297#_c_636_n 0.0140114f $X=5.745 $Y=1.595 $X2=0
+ $Y2=0
cc_327 N_A2_c_364_n N_A_647_297#_c_637_n 0.00238772f $X=5.945 $Y=1.41 $X2=0
+ $Y2=0
cc_328 A2 N_A_647_297#_c_637_n 0.0108014f $X=5.925 $Y=1.2 $X2=0 $Y2=0
cc_329 A2 N_A_647_297#_c_637_n 0.00451327f $X=5.69 $Y=1.445 $X2=0 $Y2=0
cc_330 N_A2_c_361_n N_A_647_297#_c_666_n 0.00426194f $X=4.535 $Y=1.41 $X2=0
+ $Y2=0
cc_331 N_A2_c_362_n N_VGND_c_690_n 0.00319032f $X=4.6 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A2_c_363_n N_VGND_c_692_n 0.0184132f $X=5.92 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A2_c_364_n N_VGND_c_692_n 0.00248023f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_334 A2 N_VGND_c_692_n 0.0126389f $X=5.925 $Y=1.2 $X2=0 $Y2=0
cc_335 N_A2_c_362_n N_VGND_c_696_n 0.00430182f $X=4.6 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A2_c_363_n N_VGND_c_696_n 0.00585385f $X=5.92 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A2_c_362_n N_VGND_c_701_n 0.00587489f $X=4.6 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A2_c_363_n N_VGND_c_701_n 0.0116903f $X=5.92 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A1_c_445_n N_VPWR_c_495_n 0.00450253f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A1_c_446_n N_VPWR_c_495_n 0.00309549f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A1_c_445_n N_VPWR_c_489_n 0.00513103f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_342 N_A1_c_446_n N_VPWR_c_489_n 0.00372054f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A1_c_445_n N_VPWR_c_500_n 0.00780548f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A1_c_446_n N_VPWR_c_500_n 0.00100747f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_345 N_A1_c_445_n N_VPWR_c_501_n 0.00112257f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A1_c_446_n N_VPWR_c_501_n 0.0106109f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A1_c_445_n N_A_647_297#_c_636_n 0.0111059f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_348 N_A1_c_446_n N_A_647_297#_c_636_n 0.010665f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_349 N_A1_c_442_n N_VGND_c_696_n 0.00430182f $X=4.98 $Y=0.995 $X2=0 $Y2=0
cc_350 N_A1_c_443_n N_VGND_c_696_n 0.00585385f $X=5.5 $Y=0.995 $X2=0 $Y2=0
cc_351 N_A1_c_442_n N_VGND_c_701_n 0.00613555f $X=4.98 $Y=0.995 $X2=0 $Y2=0
cc_352 N_A1_c_443_n N_VGND_c_701_n 0.0110915f $X=5.5 $Y=0.995 $X2=0 $Y2=0
cc_353 N_VPWR_c_489_n N_X_M1000_d 0.00341753f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_354 N_VPWR_c_489_n N_X_M1012_d 0.00341753f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_355 N_VPWR_M1006_s N_X_c_599_n 0.00393239f $X=1.715 $Y=1.485 $X2=0 $Y2=0
cc_356 N_VPWR_c_489_n N_A_647_297#_M1005_d 0.00364058f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_357 N_VPWR_c_489_n N_A_647_297#_M1019_d 0.00258242f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_489_n N_A_647_297#_M1014_s 0.00330361f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_489_n N_A_647_297#_M1008_s 0.00308785f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_494_n N_A_647_297#_c_640_n 0.0267689f $X=4.555 $Y=2.72 $X2=0
+ $Y2=0
cc_361 N_VPWR_c_489_n N_A_647_297#_c_640_n 0.0250745f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_362 N_VPWR_c_492_n N_A_647_297#_c_675_n 0.0063501f $X=2.82 $Y=2.36 $X2=0
+ $Y2=0
cc_363 N_VPWR_c_494_n N_A_647_297#_c_675_n 0.00770731f $X=4.555 $Y=2.72 $X2=0
+ $Y2=0
cc_364 N_VPWR_c_489_n N_A_647_297#_c_675_n 0.00625935f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_365 N_VPWR_M1002_d N_A_647_297#_c_636_n 0.00364347f $X=4.625 $Y=1.485 $X2=0
+ $Y2=0
cc_366 N_VPWR_M1020_d N_A_647_297#_c_636_n 0.00365341f $X=5.565 $Y=1.485 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_494_n N_A_647_297#_c_636_n 0.00252264f $X=4.555 $Y=2.72 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_495_n N_A_647_297#_c_636_n 0.00901445f $X=5.495 $Y=2.72 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_496_n N_A_647_297#_c_636_n 0.00845292f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_489_n N_A_647_297#_c_636_n 0.0357556f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_500_n N_A_647_297#_c_636_n 0.0195044f $X=4.77 $Y=2.36 $X2=0
+ $Y2=0
cc_372 N_VPWR_c_501_n N_A_647_297#_c_636_n 0.0195044f $X=5.71 $Y=2.36 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_494_n N_A_647_297#_c_666_n 0.00793684f $X=4.555 $Y=2.72 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_489_n N_A_647_297#_c_666_n 0.00655231f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_500_n N_A_647_297#_c_666_n 0.00787162f $X=4.77 $Y=2.36 $X2=0
+ $Y2=0
cc_376 N_X_c_593_n N_VGND_M1004_s 0.00435335f $X=2.345 $Y=0.7 $X2=0 $Y2=0
cc_377 N_X_c_593_n N_VGND_c_693_n 0.0196989f $X=2.345 $Y=0.7 $X2=0 $Y2=0
cc_378 N_X_c_593_n N_VGND_c_694_n 0.00187977f $X=2.345 $Y=0.7 $X2=0 $Y2=0
cc_379 N_X_c_589_n N_VGND_c_694_n 0.00815715f $X=1.295 $Y=0.785 $X2=0 $Y2=0
cc_380 N_X_c_589_n N_VGND_c_697_n 0.00149282f $X=1.295 $Y=0.785 $X2=0 $Y2=0
cc_381 N_X_c_593_n N_VGND_c_698_n 0.00768849f $X=2.345 $Y=0.7 $X2=0 $Y2=0
cc_382 N_X_M1001_d N_VGND_c_701_n 0.00375459f $X=1.195 $Y=0.235 $X2=0 $Y2=0
cc_383 N_X_M1007_d N_VGND_c_701_n 0.00375928f $X=2.155 $Y=0.235 $X2=0 $Y2=0
cc_384 N_X_c_593_n N_VGND_c_701_n 0.0174455f $X=2.345 $Y=0.7 $X2=0 $Y2=0
cc_385 N_X_c_589_n N_VGND_c_701_n 0.0137373f $X=1.295 $Y=0.785 $X2=0 $Y2=0
cc_386 N_A_647_297#_c_637_n N_VGND_c_692_n 0.00477372f $X=6.18 $Y=1.63 $X2=0
+ $Y2=0
cc_387 N_VGND_c_701_n A_1115_47# 0.00280308f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_388 N_VGND_c_701_n A_935_47# 0.0115413f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
