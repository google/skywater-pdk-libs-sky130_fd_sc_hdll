* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xor3_2 A B C VGND VNB VPB VPWR X
X0 VPWR B a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_1050_365# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 a_1335_297# B a_465_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_465_325# C a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X4 a_1335_297# B a_483_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X5 a_483_49# C a_81_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_483_49# a_934_297# a_1335_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VGND C a_335_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_483_49# a_934_297# a_1050_365# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X10 a_81_21# a_335_93# a_483_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X11 VGND a_1050_365# a_1335_297# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_465_325# a_934_297# a_1050_365# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X13 a_465_325# a_934_297# a_1335_297# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X14 a_1050_365# B a_465_325# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X15 a_1050_365# B a_483_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VPWR a_1050_365# a_1335_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 a_81_21# a_335_93# a_465_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_1050_365# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 VGND B a_934_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR C a_335_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X22 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
