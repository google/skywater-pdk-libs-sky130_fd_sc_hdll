# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o32ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o32ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.090000 1.075000 10.925000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.520000 1.075000 8.010000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.170000 1.075000 5.980000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.075000 3.940000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.835000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 3.730000 0.905000 ;
        RECT 0.515000 1.495000 6.130000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.085000 ;
        RECT 1.455000 1.665000 1.850000 2.085000 ;
        RECT 2.055000 0.905000 2.235000 1.495000 ;
        RECT 4.860000 1.665000 5.190000 2.085000 ;
        RECT 5.750000 1.665000 6.130000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.040000 0.085000 ;
        RECT  4.420000  0.085000  4.590000 0.545000 ;
        RECT  5.360000  0.085000  5.690000 0.545000 ;
        RECT  6.820000  0.085000  6.990000 0.545000 ;
        RECT  7.760000  0.085000  7.930000 0.545000 ;
        RECT  9.220000  0.085000  9.390000 0.545000 ;
        RECT 10.160000  0.085000 10.375000 0.545000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 11.040000 2.805000 ;
        RECT  2.410000 2.175000  2.790000 2.635000 ;
        RECT  3.350000 2.175000  3.730000 2.635000 ;
        RECT  8.670000 1.835000  8.920000 2.635000 ;
        RECT  9.690000 1.835000  9.860000 2.635000 ;
        RECT 10.675000 1.495000 10.925000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.090000 0.255000  4.200000 0.465000 ;
      RECT  0.090000 0.465000  0.345000 0.905000 ;
      RECT  0.090000 1.495000  0.345000 2.255000 ;
      RECT  0.090000 2.255000  2.240000 2.465000 ;
      RECT  1.115000 1.835000  1.285000 2.255000 ;
      RECT  2.070000 1.835000  4.200000 2.005000 ;
      RECT  2.070000 2.005000  2.240000 2.255000 ;
      RECT  3.010000 2.005000  3.180000 2.425000 ;
      RECT  3.950000 0.465000  4.200000 0.735000 ;
      RECT  3.950000 0.735000 10.925000 0.905000 ;
      RECT  3.950000 2.005000  4.200000 2.465000 ;
      RECT  4.390000 1.835000  4.640000 2.255000 ;
      RECT  4.390000 2.255000  8.480000 2.465000 ;
      RECT  4.760000 0.255000  5.140000 0.735000 ;
      RECT  5.410000 1.835000  5.580000 2.255000 ;
      RECT  5.910000 0.255000  6.580000 0.735000 ;
      RECT  6.350000 1.835000  6.520000 2.255000 ;
      RECT  6.690000 1.495000 10.410000 1.665000 ;
      RECT  6.690000 1.665000  7.070000 2.085000 ;
      RECT  7.160000 0.255000  7.540000 0.735000 ;
      RECT  7.290000 1.835000  7.460000 2.255000 ;
      RECT  7.630000 1.665000  8.010000 2.085000 ;
      RECT  8.100000 0.255000  8.840000 0.735000 ;
      RECT  8.230000 1.835000  8.480000 2.255000 ;
      RECT  9.090000 1.665000  9.470000 2.465000 ;
      RECT  9.560000 0.255000  9.940000 0.735000 ;
      RECT 10.030000 1.665000 10.410000 2.465000 ;
      RECT 10.545000 0.255000 10.925000 0.735000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o32ai_4
