* File: sky130_fd_sc_hdll__bufbuf_16.spice
* Created: Wed Sep  2 08:24:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__bufbuf_16.pex.spice"
.subckt sky130_fd_sc_hdll__bufbuf_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1037 N_A_117_297#_M1037_d N_A_M1037_g N_VGND_M1037_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.2015 PD=1.82 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_A_117_297#_M1020_g N_A_225_47#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75011.5 A=0.0975 P=1.6 MULT=1
MM1038 N_VGND_M1020_d N_A_117_297#_M1038_g N_A_225_47#_M1038_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75011 A=0.0975 P=1.6 MULT=1
MM1050 N_VGND_M1050_d N_A_117_297#_M1050_g N_A_225_47#_M1038_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75010.5 A=0.0975 P=1.6 MULT=1
MM1012 N_A_589_47#_M1012_d N_A_225_47#_M1012_g N_VGND_M1050_d VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75010.1 A=0.0975 P=1.6 MULT=1
MM1014 N_A_589_47#_M1012_d N_A_225_47#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75009.6 A=0.0975 P=1.6 MULT=1
MM1023 N_A_589_47#_M1023_d N_A_225_47#_M1023_g N_VGND_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.5 SB=75009.2 A=0.0975 P=1.6 MULT=1
MM1033 N_A_589_47#_M1023_d N_A_225_47#_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003 SB=75008.7 A=0.0975 P=1.6 MULT=1
MM1045 N_A_589_47#_M1045_d N_A_225_47#_M1045_g N_VGND_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75008.2 A=0.0975 P=1.6 MULT=1
MM1047 N_A_589_47#_M1045_d N_A_225_47#_M1047_g N_VGND_M1047_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75004 SB=75007.7 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1047_s N_A_589_47#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.4
+ SB=75007.3 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A_589_47#_M1002_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1002_d N_A_589_47#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.4
+ SB=75006.3 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A_589_47#_M1006_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.8
+ SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1006_d N_A_589_47#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.3
+ SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_589_47#_M1015_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006.8
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1015_d N_A_589_47#_M1017_g N_X_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75007.2
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_A_589_47#_M1018_g N_X_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75007.7
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1018_d N_A_589_47#_M1021_g N_X_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75008.2
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1024_d N_A_589_47#_M1024_g N_X_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75008.6
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1026 N_VGND_M1024_d N_A_589_47#_M1026_g N_X_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75009.1
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1028 N_VGND_M1028_d N_A_589_47#_M1028_g N_X_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75009.6
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1034 N_VGND_M1028_d N_A_589_47#_M1034_g N_X_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75010.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1043 N_VGND_M1043_d N_A_589_47#_M1043_g N_X_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75010.5
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1048 N_VGND_M1043_d N_A_589_47#_M1048_g N_X_M1048_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75011
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1051 N_VGND_M1051_d N_A_589_47#_M1051_g N_X_M1048_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75011.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1022 N_A_117_297#_M1022_d N_A_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.27 PD=2.54 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1027 N_VPWR_M1027_d N_A_117_297#_M1027_g N_A_225_47#_M1027_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90011.5 A=0.18 P=2.36 MULT=1
MM1035 N_VPWR_M1027_d N_A_117_297#_M1035_g N_A_225_47#_M1035_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90011 A=0.18 P=2.36 MULT=1
MM1042 N_VPWR_M1042_d N_A_117_297#_M1042_g N_A_225_47#_M1035_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001.1 SB=90010.5 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1042_d N_A_225_47#_M1005_g N_A_589_47#_M1005_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90010 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_225_47#_M1008_g N_A_589_47#_M1005_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90009.6 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1008_d N_A_225_47#_M1010_g N_A_589_47#_M1010_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90009.1 A=0.18 P=2.36 MULT=1
MM1031 N_VPWR_M1031_d N_A_225_47#_M1031_g N_A_589_47#_M1010_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003 SB=90008.6 A=0.18 P=2.36 MULT=1
MM1039 N_VPWR_M1031_d N_A_225_47#_M1039_g N_A_589_47#_M1039_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90008.2 A=0.18 P=2.36 MULT=1
MM1049 N_VPWR_M1049_d N_A_225_47#_M1049_g N_A_589_47#_M1039_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.9 SB=90007.7 A=0.18 P=2.36 MULT=1
MM1000 N_X_M1000_d N_A_589_47#_M1000_g N_VPWR_M1049_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90007.2 A=0.18 P=2.36 MULT=1
MM1004 N_X_M1000_d N_A_589_47#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.9 SB=90006.8 A=0.18 P=2.36 MULT=1
MM1009 N_X_M1009_d N_A_589_47#_M1009_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.3 SB=90006.3 A=0.18 P=2.36 MULT=1
MM1011 N_X_M1009_d N_A_589_47#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.8 SB=90005.8 A=0.18 P=2.36 MULT=1
MM1013 N_X_M1013_d N_A_589_47#_M1013_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.3 SB=90005.3 A=0.18 P=2.36 MULT=1
MM1016 N_X_M1013_d N_A_589_47#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.8 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1019 N_X_M1019_d N_A_589_47#_M1019_g N_VPWR_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.2 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1025 N_X_M1019_d N_A_589_47#_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.7 SB=90003.9 A=0.18 P=2.36 MULT=1
MM1029 N_X_M1029_d N_A_589_47#_M1029_g N_VPWR_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90008.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1030 N_X_M1029_d N_A_589_47#_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90008.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1032 N_X_M1032_d N_A_589_47#_M1032_g N_VPWR_M1030_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90009.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1036 N_X_M1032_d N_A_589_47#_M1036_g N_VPWR_M1036_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90009.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1040 N_X_M1040_d N_A_589_47#_M1040_g N_VPWR_M1036_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90010
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1041 N_X_M1040_d N_A_589_47#_M1041_g N_VPWR_M1041_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90010.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1044 N_X_M1044_d N_A_589_47#_M1044_g N_VPWR_M1041_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90011
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1046 N_X_M1044_d N_A_589_47#_M1046_g N_VPWR_M1046_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90011.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX52_noxref VNB VPB NWDIODE A=22.0206 P=30.65
*
.include "sky130_fd_sc_hdll__bufbuf_16.pxi.spice"
*
.ends
*
*
