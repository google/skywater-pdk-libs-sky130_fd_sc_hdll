* File: sky130_fd_sc_hdll__dfrtp_4.spice
* Created: Wed Sep  2 08:28:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__dfrtp_4.pex.spice"
.subckt sky130_fd_sc_hdll__dfrtp_4  VNB VPB CLK D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_CLK_M1021_g N_A_27_47#_M1021_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_211_363#_M1002_d N_A_27_47#_M1002_g N_VGND_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_468_47#_M1012_d N_D_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0920769 AS=0.2205 PD=0.91 PS=1.89 NRD=12.852 NRS=68.568 M=1 R=2.8
+ SA=75000.4 SB=75005.5 A=0.063 P=1.14 MULT=1
MM1007 N_A_583_47#_M1007_d N_A_27_47#_M1007_g N_A_468_47#_M1012_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0684 AS=0.0789231 PD=0.74 PS=0.78 NRD=18.324 NRS=33.324 M=1
+ R=2.4 SA=75001 SB=75005.8 A=0.054 P=1.02 MULT=1
MM1014 A_689_47# N_A_211_363#_M1014_g N_A_583_47#_M1007_d VNB NSHORT L=0.15
+ W=0.36 AD=0.139015 AS=0.0684 PD=1.06154 PS=0.74 NRD=110.376 NRS=14.988 M=1
+ R=2.4 SA=75001.6 SB=75005.3 A=0.054 P=1.02 MULT=1
MM1001 A_865_47# N_A_811_289#_M1001_g A_689_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.162185 PD=0.63 PS=1.23846 NRD=14.28 NRS=94.608 M=1 R=2.8
+ SA=75002.2 SB=75004 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_RESET_B_M1003_g A_865_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.127664 AS=0.0441 PD=0.990566 PS=0.63 NRD=47.136 NRS=14.28 M=1 R=2.8
+ SA=75002.5 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1032 N_A_811_289#_M1032_d N_A_583_47#_M1032_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.64 AD=0.127872 AS=0.194536 PD=1.2608 PS=1.50943 NRD=2.808 NRS=30.936 M=1
+ R=4.26667 SA=75002.2 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1005 N_A_1188_47#_M1005_d N_A_211_363#_M1005_g N_A_811_289#_M1032_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0891 AS=0.071928 PD=0.855 PS=0.7092 NRD=39.996 NRS=16.656
+ M=1 R=2.4 SA=75004 SB=75002.8 A=0.054 P=1.02 MULT=1
MM1020 A_1317_47# N_A_27_47#_M1020_g N_A_1188_47#_M1005_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0797538 AS=0.0891 PD=0.784615 PS=0.855 NRD=55.512 NRS=31.656 M=1
+ R=2.4 SA=75004.7 SB=75002.2 A=0.054 P=1.02 MULT=1
MM1018 N_VGND_M1018_d N_A_1403_21#_M1018_g A_1317_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.15645 AS=0.0930462 PD=1.165 PS=0.915385 NRD=44.28 NRS=47.58 M=1 R=2.8
+ SA=75004.6 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1029 A_1612_47# N_RESET_B_M1029_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07455 AS=0.15645 PD=0.775 PS=1.165 NRD=34.992 NRS=88.56 M=1 R=2.8
+ SA=75005.4 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_A_1403_21#_M1013_d N_A_1188_47#_M1013_g A_1612_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.07455 PD=1.36 PS=0.775 NRD=0 NRS=34.992 M=1 R=2.8
+ SA=75006 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_1403_21#_M1008_g N_Q_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1023_d N_A_1403_21#_M1023_g N_Q_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1030 N_VGND_M1023_d N_A_1403_21#_M1030_g N_Q_M1030_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1031 N_VGND_M1031_d N_A_1403_21#_M1031_g N_Q_M1030_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.104 PD=1.86 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_CLK_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1027 N_A_211_363#_M1027_d N_A_27_47#_M1027_g N_VPWR_M1004_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1024 N_A_468_47#_M1024_d N_D_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0693 AS=0.1134 PD=0.75 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1025 N_A_583_47#_M1025_d N_A_211_363#_M1025_g N_A_468_47#_M1024_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.07665 AS=0.0693 PD=0.785 PS=0.75 NRD=4.6886 NRS=21.0987 M=1
+ R=2.33333 SA=90000.7 SB=90002 A=0.0756 P=1.2 MULT=1
MM1000 N_A_699_413#_M1000_d N_A_27_47#_M1000_g N_A_583_47#_M1025_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.1197 AS=0.07665 PD=0.99 PS=0.785 NRD=133.665 NRS=35.1645
+ M=1 R=2.33333 SA=90001.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1015 N_VPWR_M1015_d N_A_811_289#_M1015_g N_A_699_413#_M1000_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.07455 AS=0.1197 PD=0.775 PS=0.99 NRD=32.8202 NRS=2.3443 M=1
+ R=2.33333 SA=90002 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1033 N_A_699_413#_M1033_d N_RESET_B_M1033_g N_VPWR_M1015_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.07455 PD=1.38 PS=0.775 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90002.5 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1022 N_A_811_289#_M1022_d N_A_583_47#_M1022_g N_VPWR_M1022_s VPB PHIGHVT
+ L=0.18 W=0.84 AD=0.1806 AS=0.2688 PD=1.60667 PS=2.32 NRD=5.8509 NRS=1.1623 M=1
+ R=4.66667 SA=90000.2 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1028 N_A_1188_47#_M1028_d N_A_27_47#_M1028_g N_A_811_289#_M1022_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0735 AS=0.0903 PD=0.77 PS=0.803333 NRD=7.0329 NRS=28.1316
+ M=1 R=2.33333 SA=90000.8 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1009 A_1388_413# N_A_211_363#_M1009_g N_A_1188_47#_M1028_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0714 AS=0.0735 PD=0.76 PS=0.77 NRD=53.9386 NRS=25.7873 M=1
+ R=2.33333 SA=90001.3 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_1403_21#_M1006_g A_1388_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0861 AS=0.0714 PD=0.83 PS=0.76 NRD=58.6272 NRS=53.9386 M=1 R=2.33333
+ SA=90001.8 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1017 N_A_1403_21#_M1017_d N_RESET_B_M1017_g N_VPWR_M1006_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.0861 PD=0.71 PS=0.83 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90002.4 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1011 N_VPWR_M1011_d N_A_1188_47#_M1011_g N_A_1403_21#_M1017_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.1176 AS=0.0609 PD=1.4 PS=0.71 NRD=7.0329 NRS=2.3443 M=1
+ R=2.33333 SA=90002.9 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_1403_21#_M1010_g N_Q_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_A_1403_21#_M1016_g N_Q_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1016_d N_A_1403_21#_M1019_g N_Q_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1026 N_VPWR_M1026_d N_A_1403_21#_M1026_g N_Q_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.315 AS=0.145 PD=2.63 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX34_noxref VNB VPB NWDIODE A=19.0674 P=26.97
c_104 VNB 0 1.94832e-19 $X=0.145 $Y=-0.085
c_217 VPB 0 1.92806e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__dfrtp_4.pxi.spice"
*
.ends
*
*
