* File: sky130_fd_sc_hdll__o22ai_4.pxi.spice
* Created: Wed Sep  2 08:45:51 2020
* 
x_PM_SKY130_FD_SC_HDLL__O22AI_4%A1 N_A1_c_111_n N_A1_M1007_g N_A1_c_102_n
+ N_A1_M1005_g N_A1_c_112_n N_A1_M1011_g N_A1_c_103_n N_A1_M1006_g N_A1_c_113_n
+ N_A1_M1012_g N_A1_c_104_n N_A1_M1019_g N_A1_c_105_n N_A1_M1027_g N_A1_c_106_n
+ N_A1_M1031_g N_A1_c_115_n N_A1_c_116_n N_A1_c_117_n N_A1_c_107_n A1
+ N_A1_c_109_n N_A1_c_110_n A1 PM_SKY130_FD_SC_HDLL__O22AI_4%A1
x_PM_SKY130_FD_SC_HDLL__O22AI_4%A2 N_A2_c_223_n N_A2_M1002_g N_A2_c_229_n
+ N_A2_M1000_g N_A2_c_224_n N_A2_M1016_g N_A2_c_230_n N_A2_M1015_g N_A2_c_225_n
+ N_A2_M1024_g N_A2_c_231_n N_A2_M1022_g N_A2_c_232_n N_A2_M1025_g N_A2_c_226_n
+ N_A2_M1026_g A2 N_A2_c_227_n N_A2_c_228_n A2 PM_SKY130_FD_SC_HDLL__O22AI_4%A2
x_PM_SKY130_FD_SC_HDLL__O22AI_4%B1 N_B1_c_304_n N_B1_M1004_g N_B1_c_312_n
+ N_B1_M1003_g N_B1_c_305_n N_B1_M1014_g N_B1_c_313_n N_B1_M1018_g N_B1_c_314_n
+ N_B1_M1023_g N_B1_c_306_n N_B1_M1020_g N_B1_c_307_n N_B1_M1030_g N_B1_c_308_n
+ N_B1_M1029_g N_B1_c_316_n N_B1_c_309_n B1 N_B1_c_310_n B1 N_B1_c_311_n
+ PM_SKY130_FD_SC_HDLL__O22AI_4%B1
x_PM_SKY130_FD_SC_HDLL__O22AI_4%B2 N_B2_c_412_n N_B2_M1009_g N_B2_c_417_n
+ N_B2_M1001_g N_B2_c_413_n N_B2_M1010_g N_B2_c_418_n N_B2_M1008_g N_B2_c_414_n
+ N_B2_M1017_g N_B2_c_419_n N_B2_M1013_g N_B2_c_420_n N_B2_M1028_g N_B2_c_415_n
+ N_B2_M1021_g B2 N_B2_c_416_n B2 PM_SKY130_FD_SC_HDLL__O22AI_4%B2
x_PM_SKY130_FD_SC_HDLL__O22AI_4%VPWR N_VPWR_M1007_s N_VPWR_M1011_s
+ N_VPWR_M1027_s N_VPWR_M1018_s N_VPWR_M1030_s N_VPWR_c_476_n N_VPWR_c_477_n
+ N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_480_n N_VPWR_c_481_n N_VPWR_c_482_n
+ N_VPWR_c_483_n N_VPWR_c_484_n N_VPWR_c_485_n N_VPWR_c_486_n N_VPWR_c_487_n
+ VPWR N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_475_n
+ PM_SKY130_FD_SC_HDLL__O22AI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O22AI_4%A_123_297# N_A_123_297#_M1007_d
+ N_A_123_297#_M1012_d N_A_123_297#_M1015_s N_A_123_297#_M1025_s
+ N_A_123_297#_c_591_n N_A_123_297#_c_617_n N_A_123_297#_c_601_n
+ N_A_123_297#_c_640_p N_A_123_297#_c_608_n N_A_123_297#_c_624_n
+ N_A_123_297#_c_610_n N_A_123_297#_c_628_n N_A_123_297#_c_607_n
+ PM_SKY130_FD_SC_HDLL__O22AI_4%A_123_297#
x_PM_SKY130_FD_SC_HDLL__O22AI_4%Y N_Y_M1004_d N_Y_M1020_d N_Y_M1010_s
+ N_Y_M1021_s N_Y_M1000_d N_Y_M1022_d N_Y_M1001_d N_Y_M1013_d N_Y_c_654_n
+ N_Y_c_669_n N_Y_c_671_n N_Y_c_646_n N_Y_c_647_n N_Y_c_686_n N_Y_c_650_n
+ N_Y_c_648_n N_Y_c_658_n N_Y_c_659_n N_Y_c_694_n N_Y_c_695_n Y Y
+ PM_SKY130_FD_SC_HDLL__O22AI_4%Y
x_PM_SKY130_FD_SC_HDLL__O22AI_4%A_885_297# N_A_885_297#_M1003_d
+ N_A_885_297#_M1023_d N_A_885_297#_M1008_s N_A_885_297#_M1028_s
+ N_A_885_297#_c_770_n N_A_885_297#_c_774_n N_A_885_297#_c_778_n
+ N_A_885_297#_c_791_n N_A_885_297#_c_780_n N_A_885_297#_c_776_n
+ N_A_885_297#_c_777_n N_A_885_297#_c_798_n N_A_885_297#_c_800_n
+ PM_SKY130_FD_SC_HDLL__O22AI_4%A_885_297#
x_PM_SKY130_FD_SC_HDLL__O22AI_4%A_33_47# N_A_33_47#_M1005_d N_A_33_47#_M1006_d
+ N_A_33_47#_M1002_d N_A_33_47#_M1024_d N_A_33_47#_M1031_d N_A_33_47#_M1014_s
+ N_A_33_47#_M1009_d N_A_33_47#_M1017_d N_A_33_47#_M1029_s N_A_33_47#_c_818_n
+ N_A_33_47#_c_819_n N_A_33_47#_c_820_n N_A_33_47#_c_834_n N_A_33_47#_c_821_n
+ N_A_33_47#_c_839_n N_A_33_47#_c_822_n N_A_33_47#_c_859_n N_A_33_47#_c_823_n
+ N_A_33_47#_c_844_n N_A_33_47#_c_845_n N_A_33_47#_c_824_n N_A_33_47#_c_825_n
+ N_A_33_47#_c_826_n N_A_33_47#_c_827_n PM_SKY130_FD_SC_HDLL__O22AI_4%A_33_47#
x_PM_SKY130_FD_SC_HDLL__O22AI_4%VGND N_VGND_M1005_s N_VGND_M1019_s
+ N_VGND_M1016_s N_VGND_M1026_s N_VGND_c_937_n N_VGND_c_938_n N_VGND_c_939_n
+ N_VGND_c_940_n N_VGND_c_941_n N_VGND_c_942_n N_VGND_c_943_n N_VGND_c_944_n
+ N_VGND_c_945_n N_VGND_c_946_n VGND N_VGND_c_947_n N_VGND_c_948_n
+ N_VGND_c_949_n PM_SKY130_FD_SC_HDLL__O22AI_4%VGND
cc_1 VNB N_A1_c_102_n 0.0219752f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_2 VNB N_A1_c_103_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=0.995
cc_3 VNB N_A1_c_104_n 0.0164985f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=0.995
cc_4 VNB N_A1_c_105_n 0.0226064f $X=-0.19 $Y=-0.24 $X2=3.815 $Y2=1.41
cc_5 VNB N_A1_c_106_n 0.017129f $X=-0.19 $Y=-0.24 $X2=3.84 $Y2=0.995
cc_6 VNB N_A1_c_107_n 0.00412135f $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.16
cc_7 VNB A1 0.00149193f $X=-0.19 $Y=-0.24 $X2=1.165 $Y2=1.105
cc_8 VNB N_A1_c_109_n 0.0643539f $X=-0.19 $Y=-0.24 $X2=1.465 $Y2=1.202
cc_9 VNB N_A1_c_110_n 0.0174592f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.175
cc_10 VNB N_A2_c_223_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.41
cc_11 VNB N_A2_c_224_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=1.41
cc_12 VNB N_A2_c_225_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.465 $Y2=1.41
cc_13 VNB N_A2_c_226_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=3.84 $Y2=0.995
cc_14 VNB N_A2_c_227_n 0.00275279f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.202
cc_15 VNB N_A2_c_228_n 0.0725593f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.202
cc_16 VNB N_B1_c_304_n 0.0167043f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.41
cc_17 VNB N_B1_c_305_n 0.0173774f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=1.41
cc_18 VNB N_B1_c_306_n 0.0171738f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=0.995
cc_19 VNB N_B1_c_307_n 0.0292917f $X=-0.19 $Y=-0.24 $X2=3.815 $Y2=1.41
cc_20 VNB N_B1_c_308_n 0.019994f $X=-0.19 $Y=-0.24 $X2=3.84 $Y2=0.995
cc_21 VNB N_B1_c_309_n 0.00111724f $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.16
cc_22 VNB N_B1_c_310_n 0.0583907f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.16
cc_23 VNB N_B1_c_311_n 0.00297731f $X=-0.19 $Y=-0.24 $X2=3.815 $Y2=1.16
cc_24 VNB N_B2_c_412_n 0.0167331f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.41
cc_25 VNB N_B2_c_413_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=1.41
cc_26 VNB N_B2_c_414_n 0.0174167f $X=-0.19 $Y=-0.24 $X2=1.465 $Y2=1.41
cc_27 VNB N_B2_c_415_n 0.0176314f $X=-0.19 $Y=-0.24 $X2=3.84 $Y2=0.995
cc_28 VNB N_B2_c_416_n 0.0748537f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.202
cc_29 VNB N_VPWR_c_475_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_646_n 0.00106329f $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.16
cc_31 VNB N_Y_c_647_n 0.0105127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_648_n 0.0249014f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.202
cc_33 VNB N_A_33_47#_c_818_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.16
cc_34 VNB N_A_33_47#_c_819_n 0.00258371f $X=-0.19 $Y=-0.24 $X2=3.827 $Y2=1.53
cc_35 VNB N_A_33_47#_c_820_n 0.0104861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_33_47#_c_821_n 0.00424033f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.202
cc_37 VNB N_A_33_47#_c_822_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.202
cc_38 VNB N_A_33_47#_c_823_n 0.0111224f $X=-0.19 $Y=-0.24 $X2=3.815 $Y2=1.16
cc_39 VNB N_A_33_47#_c_824_n 0.0103442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_33_47#_c_825_n 0.00232405f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_33_47#_c_826_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_33_47#_c_827_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_937_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=0.56
cc_44 VNB N_VGND_c_938_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=3.815 $Y2=1.985
cc_45 VNB N_VGND_c_939_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=3.625 $Y2=1.53
cc_46 VNB N_VGND_c_940_n 0.00467885f $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.16
cc_47 VNB N_VGND_c_941_n 0.0192906f $X=-0.19 $Y=-0.24 $X2=3.827 $Y2=1.53
cc_48 VNB N_VGND_c_942_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_943_n 0.019187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_944_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_945_n 0.0193072f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.202
cc_52 VNB N_VGND_c_946_n 0.00323927f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.202
cc_53 VNB N_VGND_c_947_n 0.107043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_948_n 0.394167f $X=-0.19 $Y=-0.24 $X2=1.207 $Y2=1.175
cc_55 VNB N_VGND_c_949_n 0.0229511f $X=-0.19 $Y=-0.24 $X2=1.407 $Y2=1.175
cc_56 VPB N_A1_c_111_n 0.0200169f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.41
cc_57 VPB N_A1_c_112_n 0.01623f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=1.41
cc_58 VPB N_A1_c_113_n 0.0156258f $X=-0.19 $Y=1.305 $X2=1.465 $Y2=1.41
cc_59 VPB N_A1_c_105_n 0.0253766f $X=-0.19 $Y=1.305 $X2=3.815 $Y2=1.41
cc_60 VPB N_A1_c_115_n 0.012067f $X=-0.19 $Y=1.305 $X2=3.625 $Y2=1.53
cc_61 VPB N_A1_c_116_n 3.20327e-19 $X=-0.19 $Y=1.305 $X2=1.565 $Y2=1.53
cc_62 VPB N_A1_c_117_n 0.00160641f $X=-0.19 $Y=1.305 $X2=1.407 $Y2=1.445
cc_63 VPB N_A1_c_107_n 0.00292279f $X=-0.19 $Y=1.305 $X2=3.79 $Y2=1.16
cc_64 VPB N_A1_c_109_n 0.0392633f $X=-0.19 $Y=1.305 $X2=1.465 $Y2=1.202
cc_65 VPB N_A2_c_229_n 0.01598f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_66 VPB N_A2_c_230_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=0.995
cc_67 VPB N_A2_c_231_n 0.0158907f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=0.995
cc_68 VPB N_A2_c_232_n 0.0159964f $X=-0.19 $Y=1.305 $X2=3.815 $Y2=1.41
cc_69 VPB N_A2_c_228_n 0.0449077f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.202
cc_70 VPB N_B1_c_312_n 0.016212f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_71 VPB N_B1_c_313_n 0.0158859f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=0.995
cc_72 VPB N_B1_c_314_n 0.0156395f $X=-0.19 $Y=1.305 $X2=1.465 $Y2=1.41
cc_73 VPB N_B1_c_307_n 0.0311051f $X=-0.19 $Y=1.305 $X2=3.815 $Y2=1.41
cc_74 VPB N_B1_c_316_n 0.011552f $X=-0.19 $Y=1.305 $X2=3.625 $Y2=1.53
cc_75 VPB N_B1_c_309_n 0.00234935f $X=-0.19 $Y=1.305 $X2=3.79 $Y2=1.16
cc_76 VPB N_B1_c_310_n 0.0353049f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.16
cc_77 VPB N_B1_c_311_n 0.001579f $X=-0.19 $Y=1.305 $X2=3.815 $Y2=1.16
cc_78 VPB N_B2_c_417_n 0.0159762f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_79 VPB N_B2_c_418_n 0.0158727f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=0.995
cc_80 VPB N_B2_c_419_n 0.0158729f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=0.995
cc_81 VPB N_B2_c_420_n 0.015978f $X=-0.19 $Y=1.305 $X2=3.815 $Y2=1.41
cc_82 VPB N_B2_c_416_n 0.04485f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.202
cc_83 VPB N_VPWR_c_476_n 0.012247f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=0.995
cc_84 VPB N_VPWR_c_477_n 0.00937472f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=0.56
cc_85 VPB N_VPWR_c_478_n 0.0195604f $X=-0.19 $Y=1.305 $X2=3.84 $Y2=0.995
cc_86 VPB N_VPWR_c_479_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.565 $Y2=1.53
cc_87 VPB N_VPWR_c_480_n 0.00498084f $X=-0.19 $Y=1.305 $X2=3.79 $Y2=1.16
cc_88 VPB N_VPWR_c_481_n 0.00510984f $X=-0.19 $Y=1.305 $X2=1.165 $Y2=1.105
cc_89 VPB N_VPWR_c_482_n 0.0154711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_483_n 0.0190376f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.202
cc_91 VPB N_VPWR_c_484_n 0.0619203f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.16
cc_92 VPB N_VPWR_c_485_n 0.00420242f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.16
cc_93 VPB N_VPWR_c_486_n 0.0200246f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.202
cc_94 VPB N_VPWR_c_487_n 0.00459045f $X=-0.19 $Y=1.305 $X2=1.35 $Y2=1.202
cc_95 VPB N_VPWR_c_488_n 0.0611287f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_489_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_475_n 0.0480802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_123_297#_c_591_n 0.00231366f $X=-0.19 $Y=1.305 $X2=1.465 $Y2=1.985
cc_99 VPB N_Y_c_646_n 0.00319318f $X=-0.19 $Y=1.305 $X2=3.79 $Y2=1.16
cc_100 VPB N_Y_c_650_n 0.010711f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.16
cc_101 VPB N_Y_c_648_n 0.0221969f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.202
cc_102 N_A1_c_104_n N_A2_c_223_n 0.0239161f $X=1.49 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_103 N_A1_c_113_n N_A2_c_229_n 0.0226278f $X=1.465 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A1_c_115_n N_A2_c_229_n 0.0152542f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_105 N_A1_c_117_n N_A2_c_229_n 7.03078e-19 $X=1.407 $Y=1.445 $X2=0 $Y2=0
cc_106 N_A1_c_115_n N_A2_c_230_n 0.01191f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_107 N_A1_c_115_n N_A2_c_231_n 0.011867f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_108 N_A1_c_105_n N_A2_c_232_n 0.0378352f $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A1_c_115_n N_A2_c_232_n 0.0112841f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_110 N_A1_c_107_n N_A2_c_232_n 0.00102531f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A1_c_106_n N_A2_c_226_n 0.0212656f $X=3.84 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A1_c_105_n N_A2_c_227_n 2.32333e-19 $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A1_c_115_n N_A2_c_227_n 0.113835f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_114 N_A1_c_107_n N_A2_c_227_n 0.0161602f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_115 A1 N_A2_c_227_n 0.0115402f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_116 N_A1_c_109_n N_A2_c_227_n 2.49913e-19 $X=1.465 $Y=1.202 $X2=0 $Y2=0
cc_117 N_A1_c_105_n N_A2_c_228_n 0.0263635f $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A1_c_115_n N_A2_c_228_n 0.0231495f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_119 N_A1_c_117_n N_A2_c_228_n 9.22604e-19 $X=1.407 $Y=1.445 $X2=0 $Y2=0
cc_120 N_A1_c_107_n N_A2_c_228_n 0.00400307f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_121 A1 N_A2_c_228_n 2.49913e-19 $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A1_c_109_n N_A2_c_228_n 0.0239161f $X=1.465 $Y=1.202 $X2=0 $Y2=0
cc_123 N_A1_c_106_n N_B1_c_304_n 0.00984352f $X=3.84 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_124 N_A1_c_105_n N_B1_c_312_n 0.0297781f $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A1_c_107_n N_B1_c_312_n 8.79448e-19 $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A1_c_105_n N_B1_c_310_n 0.0203555f $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A1_c_107_n N_B1_c_310_n 0.00286642f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A1_c_116_n N_VPWR_M1011_s 0.00230525f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_129 N_A1_c_107_n N_VPWR_M1027_s 0.00181837f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A1_c_111_n N_VPWR_c_477_n 0.00578236f $X=0.525 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A1_c_109_n N_VPWR_c_477_n 8.41451e-19 $X=1.465 $Y=1.202 $X2=0 $Y2=0
cc_132 N_A1_c_110_n N_VPWR_c_477_n 0.0210492f $X=1.25 $Y=1.175 $X2=0 $Y2=0
cc_133 N_A1_c_111_n N_VPWR_c_478_n 0.00702461f $X=0.525 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A1_c_112_n N_VPWR_c_478_n 0.00702461f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A1_c_112_n N_VPWR_c_479_n 0.00300743f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A1_c_113_n N_VPWR_c_479_n 0.00300743f $X=1.465 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A1_c_105_n N_VPWR_c_480_n 0.00443541f $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A1_c_113_n N_VPWR_c_484_n 0.00702461f $X=1.465 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A1_c_105_n N_VPWR_c_484_n 0.00673617f $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A1_c_111_n N_VPWR_c_475_n 0.0133474f $X=0.525 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A1_c_112_n N_VPWR_c_475_n 0.00693457f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A1_c_113_n N_VPWR_c_475_n 0.00695979f $X=1.465 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A1_c_105_n N_VPWR_c_475_n 0.00708752f $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A1_c_115_n N_A_123_297#_M1012_d 0.00183902f $X=3.625 $Y=1.53 $X2=0
+ $Y2=0
cc_145 N_A1_c_115_n N_A_123_297#_M1015_s 0.00187547f $X=3.625 $Y=1.53 $X2=0
+ $Y2=0
cc_146 N_A1_c_115_n N_A_123_297#_M1025_s 0.00172342f $X=3.625 $Y=1.53 $X2=0
+ $Y2=0
cc_147 N_A1_c_107_n N_A_123_297#_M1025_s 7.76441e-19 $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A1_c_111_n N_A_123_297#_c_591_n 3.55815e-19 $X=0.525 $Y=1.41 $X2=0
+ $Y2=0
cc_149 N_A1_c_112_n N_A_123_297#_c_591_n 4.44016e-19 $X=0.995 $Y=1.41 $X2=0
+ $Y2=0
cc_150 N_A1_c_116_n N_A_123_297#_c_591_n 0.00532569f $X=1.565 $Y=1.53 $X2=0
+ $Y2=0
cc_151 N_A1_c_109_n N_A_123_297#_c_591_n 0.00658737f $X=1.465 $Y=1.202 $X2=0
+ $Y2=0
cc_152 N_A1_c_110_n N_A_123_297#_c_591_n 0.0202219f $X=1.25 $Y=1.175 $X2=0 $Y2=0
cc_153 N_A1_c_112_n N_A_123_297#_c_601_n 0.0132594f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A1_c_113_n N_A_123_297#_c_601_n 0.0112647f $X=1.465 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A1_c_115_n N_A_123_297#_c_601_n 0.014075f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_156 N_A1_c_116_n N_A_123_297#_c_601_n 0.0188459f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_157 N_A1_c_109_n N_A_123_297#_c_601_n 0.00332181f $X=1.465 $Y=1.202 $X2=0
+ $Y2=0
cc_158 N_A1_c_110_n N_A_123_297#_c_601_n 0.00936841f $X=1.25 $Y=1.175 $X2=0
+ $Y2=0
cc_159 N_A1_c_105_n N_A_123_297#_c_607_n 0.00441302f $X=3.815 $Y=1.41 $X2=0
+ $Y2=0
cc_160 N_A1_c_115_n N_Y_M1000_d 0.00187091f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_161 N_A1_c_115_n N_Y_M1022_d 0.00187091f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_162 N_A1_c_115_n N_Y_c_654_n 0.0371166f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_163 N_A1_c_105_n N_Y_c_646_n 9.95759e-19 $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A1_c_106_n N_Y_c_646_n 4.63754e-19 $X=3.84 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_107_n N_Y_c_646_n 0.0265298f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A1_c_115_n N_Y_c_658_n 0.0184746f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_167 N_A1_c_105_n N_Y_c_659_n 0.0137372f $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A1_c_115_n N_Y_c_659_n 0.0218268f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_169 N_A1_c_107_n N_Y_c_659_n 0.0221538f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A1_c_115_n Y 0.0135474f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_171 N_A1_c_102_n N_A_33_47#_c_819_n 0.0110832f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A1_c_103_n N_A_33_47#_c_819_n 0.00622594f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A1_c_109_n N_A_33_47#_c_819_n 0.00403238f $X=1.465 $Y=1.202 $X2=0 $Y2=0
cc_174 N_A1_c_110_n N_A_33_47#_c_819_n 0.0398177f $X=1.25 $Y=1.175 $X2=0 $Y2=0
cc_175 N_A1_c_109_n N_A_33_47#_c_820_n 0.00201748f $X=1.465 $Y=1.202 $X2=0 $Y2=0
cc_176 N_A1_c_110_n N_A_33_47#_c_820_n 0.0277903f $X=1.25 $Y=1.175 $X2=0 $Y2=0
cc_177 N_A1_c_102_n N_A_33_47#_c_834_n 5.82315e-19 $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A1_c_103_n N_A_33_47#_c_834_n 0.00850899f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A1_c_104_n N_A_33_47#_c_821_n 0.0103603f $X=1.49 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A1_c_115_n N_A_33_47#_c_821_n 0.00911016f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_181 A1 N_A_33_47#_c_821_n 0.0127403f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A1_c_104_n N_A_33_47#_c_839_n 5.32212e-19 $X=1.49 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A1_c_105_n N_A_33_47#_c_823_n 0.00442788f $X=3.815 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A1_c_106_n N_A_33_47#_c_823_n 0.00861051f $X=3.84 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A1_c_115_n N_A_33_47#_c_823_n 0.00608471f $X=3.625 $Y=1.53 $X2=0 $Y2=0
cc_186 N_A1_c_107_n N_A_33_47#_c_823_n 0.0330607f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A1_c_106_n N_A_33_47#_c_844_n 0.00373464f $X=3.84 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_106_n N_A_33_47#_c_845_n 0.00499625f $X=3.84 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_103_n N_A_33_47#_c_825_n 0.00273722f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_190 A1 N_A_33_47#_c_825_n 0.0126709f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_191 N_A1_c_109_n N_A_33_47#_c_825_n 0.00358162f $X=1.465 $Y=1.202 $X2=0 $Y2=0
cc_192 N_A1_c_110_n N_A_33_47#_c_825_n 0.0186972f $X=1.25 $Y=1.175 $X2=0 $Y2=0
cc_193 N_A1_c_102_n N_VGND_c_937_n 0.00276126f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A1_c_103_n N_VGND_c_937_n 0.00359159f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A1_c_104_n N_VGND_c_938_n 0.00268723f $X=1.49 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_106_n N_VGND_c_940_n 0.00358858f $X=3.84 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A1_c_103_n N_VGND_c_941_n 0.00396605f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A1_c_104_n N_VGND_c_941_n 0.00439206f $X=1.49 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_106_n N_VGND_c_947_n 0.00395719f $X=3.84 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A1_c_102_n N_VGND_c_948_n 0.00703627f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A1_c_103_n N_VGND_c_948_n 0.00581484f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A1_c_104_n N_VGND_c_948_n 0.00606547f $X=1.49 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A1_c_106_n N_VGND_c_948_n 0.00587228f $X=3.84 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A1_c_102_n N_VGND_c_949_n 0.00437852f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A2_c_229_n N_VPWR_c_484_n 0.00429453f $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A2_c_230_n N_VPWR_c_484_n 0.00429453f $X=2.405 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A2_c_231_n N_VPWR_c_484_n 0.00429453f $X=2.875 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A2_c_232_n N_VPWR_c_484_n 0.00429453f $X=3.345 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A2_c_229_n N_VPWR_c_475_n 0.00609021f $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A2_c_230_n N_VPWR_c_475_n 0.00606499f $X=2.405 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A2_c_231_n N_VPWR_c_475_n 0.00606499f $X=2.875 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A2_c_232_n N_VPWR_c_475_n 0.00609021f $X=3.345 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A2_c_229_n N_A_123_297#_c_608_n 0.0122046f $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A2_c_230_n N_A_123_297#_c_608_n 0.0100164f $X=2.405 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A2_c_231_n N_A_123_297#_c_610_n 0.0099733f $X=2.875 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A2_c_232_n N_A_123_297#_c_610_n 0.0099733f $X=3.345 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A2_c_230_n N_Y_c_654_n 0.0108425f $X=2.405 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A2_c_231_n N_Y_c_654_n 0.0108425f $X=2.875 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A2_c_229_n N_Y_c_658_n 0.00662959f $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A2_c_232_n N_Y_c_659_n 0.0108425f $X=3.345 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A2_c_223_n N_A_33_47#_c_821_n 0.00845772f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_c_227_n N_A_33_47#_c_821_n 0.00820272f $X=3.23 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A2_c_223_n N_A_33_47#_c_839_n 0.00644736f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A2_c_224_n N_A_33_47#_c_839_n 0.00686626f $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A2_c_225_n N_A_33_47#_c_839_n 5.45498e-19 $X=2.85 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A2_c_224_n N_A_33_47#_c_822_n 0.00901745f $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A2_c_225_n N_A_33_47#_c_822_n 0.00901745f $X=2.85 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A2_c_227_n N_A_33_47#_c_822_n 0.0397461f $X=3.23 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A2_c_228_n N_A_33_47#_c_822_n 0.00345541f $X=3.345 $Y=1.202 $X2=0 $Y2=0
cc_230 N_A2_c_224_n N_A_33_47#_c_859_n 5.24597e-19 $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A2_c_225_n N_A_33_47#_c_859_n 0.00651696f $X=2.85 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A2_c_226_n N_A_33_47#_c_823_n 0.0106793f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A2_c_227_n N_A_33_47#_c_823_n 0.0117061f $X=3.23 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A2_c_226_n N_A_33_47#_c_845_n 5.51303e-19 $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A2_c_223_n N_A_33_47#_c_826_n 0.00132158f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A2_c_224_n N_A_33_47#_c_826_n 0.00116636f $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A2_c_227_n N_A_33_47#_c_826_n 0.0306016f $X=3.23 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A2_c_228_n N_A_33_47#_c_826_n 0.00358305f $X=3.345 $Y=1.202 $X2=0 $Y2=0
cc_239 N_A2_c_225_n N_A_33_47#_c_827_n 0.00119564f $X=2.85 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A2_c_227_n N_A_33_47#_c_827_n 0.0307352f $X=3.23 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A2_c_228_n N_A_33_47#_c_827_n 0.00486271f $X=3.345 $Y=1.202 $X2=0 $Y2=0
cc_242 N_A2_c_223_n N_VGND_c_938_n 0.00268723f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A2_c_224_n N_VGND_c_939_n 0.00379224f $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A2_c_225_n N_VGND_c_939_n 0.00276126f $X=2.85 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A2_c_226_n N_VGND_c_940_n 0.00276126f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A2_c_223_n N_VGND_c_943_n 0.00424416f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A2_c_224_n N_VGND_c_943_n 0.00423334f $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A2_c_225_n N_VGND_c_945_n 0.00423334f $X=2.85 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A2_c_226_n N_VGND_c_945_n 0.00439206f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A2_c_223_n N_VGND_c_948_n 0.00589024f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A2_c_224_n N_VGND_c_948_n 0.006093f $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A2_c_225_n N_VGND_c_948_n 0.00608558f $X=2.85 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A2_c_226_n N_VGND_c_948_n 0.00629903f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_254 N_B1_c_306_n N_B2_c_412_n 0.0271098f $X=5.3 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_255 N_B1_c_314_n N_B2_c_417_n 0.0225943f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B1_c_316_n N_B2_c_417_n 0.0174354f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_257 N_B1_c_311_n N_B2_c_417_n 9.74913e-19 $X=5.49 $Y=1.305 $X2=0 $Y2=0
cc_258 N_B1_c_316_n N_B2_c_418_n 0.01191f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_259 N_B1_c_316_n N_B2_c_419_n 0.01191f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_260 N_B1_c_307_n N_B2_c_420_n 0.0372921f $X=7.625 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B1_c_316_n N_B2_c_420_n 0.0130729f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_262 N_B1_c_309_n N_B2_c_420_n 7.32389e-19 $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B1_c_308_n N_B2_c_415_n 0.0220973f $X=7.65 $Y=0.995 $X2=0 $Y2=0
cc_264 N_B1_c_307_n B2 6.03085e-19 $X=7.625 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B1_c_316_n B2 0.10621f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_266 N_B1_c_309_n B2 0.00974021f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B1_c_310_n B2 2.11472e-19 $X=5.275 $Y=1.202 $X2=0 $Y2=0
cc_268 N_B1_c_311_n B2 0.0176522f $X=5.49 $Y=1.305 $X2=0 $Y2=0
cc_269 N_B1_c_307_n N_B2_c_416_n 0.0262867f $X=7.625 $Y=1.41 $X2=0 $Y2=0
cc_270 N_B1_c_316_n N_B2_c_416_n 0.0232657f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_271 N_B1_c_309_n N_B2_c_416_n 0.0037099f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B1_c_310_n N_B2_c_416_n 0.0256085f $X=5.275 $Y=1.202 $X2=0 $Y2=0
cc_273 N_B1_c_311_n N_B2_c_416_n 0.00748181f $X=5.49 $Y=1.305 $X2=0 $Y2=0
cc_274 N_B1_c_311_n N_VPWR_M1018_s 0.00195154f $X=5.49 $Y=1.305 $X2=0 $Y2=0
cc_275 N_B1_c_312_n N_VPWR_c_480_n 0.00417414f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B1_c_313_n N_VPWR_c_481_n 0.00293739f $X=4.805 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B1_c_314_n N_VPWR_c_481_n 0.00299501f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_278 N_B1_c_307_n N_VPWR_c_483_n 0.00482583f $X=7.625 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B1_c_312_n N_VPWR_c_486_n 0.00597712f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_280 N_B1_c_313_n N_VPWR_c_486_n 0.00702461f $X=4.805 $Y=1.41 $X2=0 $Y2=0
cc_281 N_B1_c_314_n N_VPWR_c_488_n 0.00702461f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_282 N_B1_c_307_n N_VPWR_c_488_n 0.00702461f $X=7.625 $Y=1.41 $X2=0 $Y2=0
cc_283 N_B1_c_312_n N_VPWR_c_475_n 0.00674904f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_284 N_B1_c_313_n N_VPWR_c_475_n 0.00695966f $X=4.805 $Y=1.41 $X2=0 $Y2=0
cc_285 N_B1_c_314_n N_VPWR_c_475_n 0.00695979f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_286 N_B1_c_307_n N_VPWR_c_475_n 0.00798959f $X=7.625 $Y=1.41 $X2=0 $Y2=0
cc_287 N_B1_c_316_n N_Y_M1001_d 0.00187091f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_288 N_B1_c_316_n N_Y_M1013_d 0.00187091f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_289 N_B1_c_312_n N_Y_c_669_n 0.00565588f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_290 N_B1_c_313_n N_Y_c_669_n 9.67426e-19 $X=4.805 $Y=1.41 $X2=0 $Y2=0
cc_291 N_B1_c_304_n N_Y_c_671_n 0.00226162f $X=4.31 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B1_c_304_n N_Y_c_646_n 0.00353043f $X=4.31 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B1_c_312_n N_Y_c_646_n 0.0130916f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_294 N_B1_c_305_n N_Y_c_646_n 0.00378693f $X=4.78 $Y=0.995 $X2=0 $Y2=0
cc_295 N_B1_c_313_n N_Y_c_646_n 0.00132304f $X=4.805 $Y=1.41 $X2=0 $Y2=0
cc_296 N_B1_c_310_n N_Y_c_646_n 0.023979f $X=5.275 $Y=1.202 $X2=0 $Y2=0
cc_297 N_B1_c_311_n N_Y_c_646_n 0.0493476f $X=5.49 $Y=1.305 $X2=0 $Y2=0
cc_298 N_B1_c_305_n N_Y_c_647_n 0.0102655f $X=4.78 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B1_c_306_n N_Y_c_647_n 0.00909383f $X=5.3 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B1_c_307_n N_Y_c_647_n 0.00283632f $X=7.625 $Y=1.41 $X2=0 $Y2=0
cc_301 N_B1_c_308_n N_Y_c_647_n 0.0103189f $X=7.65 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B1_c_316_n N_Y_c_647_n 0.0115516f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_303 N_B1_c_309_n N_Y_c_647_n 0.0177167f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_304 N_B1_c_310_n N_Y_c_647_n 0.00694474f $X=5.275 $Y=1.202 $X2=0 $Y2=0
cc_305 N_B1_c_311_n N_Y_c_647_n 0.0501453f $X=5.49 $Y=1.305 $X2=0 $Y2=0
cc_306 N_B1_c_316_n N_Y_c_686_n 0.0371166f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_307 N_B1_c_307_n N_Y_c_650_n 0.0169016f $X=7.625 $Y=1.41 $X2=0 $Y2=0
cc_308 N_B1_c_316_n N_Y_c_650_n 0.0386255f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_309 N_B1_c_307_n N_Y_c_648_n 0.0164716f $X=7.625 $Y=1.41 $X2=0 $Y2=0
cc_310 N_B1_c_308_n N_Y_c_648_n 0.00621452f $X=7.65 $Y=0.995 $X2=0 $Y2=0
cc_311 N_B1_c_316_n N_Y_c_648_n 0.0085043f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_312 N_B1_c_309_n N_Y_c_648_n 0.0349273f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_313 N_B1_c_312_n N_Y_c_659_n 0.00813042f $X=4.335 $Y=1.41 $X2=0 $Y2=0
cc_314 N_B1_c_316_n N_Y_c_694_n 0.0135474f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_315 N_B1_c_316_n N_Y_c_695_n 0.0135474f $X=7.465 $Y=1.53 $X2=0 $Y2=0
cc_316 N_B1_c_316_n N_A_885_297#_M1023_d 0.00113743f $X=7.465 $Y=1.53 $X2=0
+ $Y2=0
cc_317 N_B1_c_311_n N_A_885_297#_M1023_d 7.52159e-19 $X=5.49 $Y=1.305 $X2=0
+ $Y2=0
cc_318 N_B1_c_316_n N_A_885_297#_M1008_s 0.00187547f $X=7.465 $Y=1.53 $X2=0
+ $Y2=0
cc_319 N_B1_c_316_n N_A_885_297#_M1028_s 0.00185904f $X=7.465 $Y=1.53 $X2=0
+ $Y2=0
cc_320 N_B1_c_313_n N_A_885_297#_c_770_n 0.0136249f $X=4.805 $Y=1.41 $X2=0 $Y2=0
cc_321 N_B1_c_314_n N_A_885_297#_c_770_n 0.011229f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_322 N_B1_c_310_n N_A_885_297#_c_770_n 0.00102745f $X=5.275 $Y=1.202 $X2=0
+ $Y2=0
cc_323 N_B1_c_311_n N_A_885_297#_c_770_n 0.0537421f $X=5.49 $Y=1.305 $X2=0 $Y2=0
cc_324 N_B1_c_312_n N_A_885_297#_c_774_n 0.00125802f $X=4.335 $Y=1.41 $X2=0
+ $Y2=0
cc_325 N_B1_c_310_n N_A_885_297#_c_774_n 0.00367845f $X=5.275 $Y=1.202 $X2=0
+ $Y2=0
cc_326 N_B1_c_312_n N_A_885_297#_c_776_n 0.00694965f $X=4.335 $Y=1.41 $X2=0
+ $Y2=0
cc_327 N_B1_c_312_n N_A_885_297#_c_777_n 0.00369299f $X=4.335 $Y=1.41 $X2=0
+ $Y2=0
cc_328 N_B1_c_304_n N_A_33_47#_c_824_n 0.0130858f $X=4.31 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B1_c_305_n N_A_33_47#_c_824_n 0.00931157f $X=4.78 $Y=0.995 $X2=0 $Y2=0
cc_330 N_B1_c_306_n N_A_33_47#_c_824_n 0.00886996f $X=5.3 $Y=0.995 $X2=0 $Y2=0
cc_331 N_B1_c_308_n N_A_33_47#_c_824_n 0.00923997f $X=7.65 $Y=0.995 $X2=0 $Y2=0
cc_332 N_B1_c_310_n N_A_33_47#_c_824_n 4.02536e-19 $X=5.275 $Y=1.202 $X2=0 $Y2=0
cc_333 N_B1_c_304_n N_VGND_c_947_n 0.00357877f $X=4.31 $Y=0.995 $X2=0 $Y2=0
cc_334 N_B1_c_305_n N_VGND_c_947_n 0.00357877f $X=4.78 $Y=0.995 $X2=0 $Y2=0
cc_335 N_B1_c_306_n N_VGND_c_947_n 0.00357877f $X=5.3 $Y=0.995 $X2=0 $Y2=0
cc_336 N_B1_c_308_n N_VGND_c_947_n 0.00357877f $X=7.65 $Y=0.995 $X2=0 $Y2=0
cc_337 N_B1_c_304_n N_VGND_c_948_n 0.00550244f $X=4.31 $Y=0.995 $X2=0 $Y2=0
cc_338 N_B1_c_305_n N_VGND_c_948_n 0.00559933f $X=4.78 $Y=0.995 $X2=0 $Y2=0
cc_339 N_B1_c_306_n N_VGND_c_948_n 0.00549573f $X=5.3 $Y=0.995 $X2=0 $Y2=0
cc_340 N_B1_c_308_n N_VGND_c_948_n 0.00645241f $X=7.65 $Y=0.995 $X2=0 $Y2=0
cc_341 N_B2_c_417_n N_VPWR_c_488_n 0.00429453f $X=5.745 $Y=1.41 $X2=0 $Y2=0
cc_342 N_B2_c_418_n N_VPWR_c_488_n 0.00429453f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_343 N_B2_c_419_n N_VPWR_c_488_n 0.00429453f $X=6.685 $Y=1.41 $X2=0 $Y2=0
cc_344 N_B2_c_420_n N_VPWR_c_488_n 0.00429453f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_345 N_B2_c_417_n N_VPWR_c_475_n 0.00609021f $X=5.745 $Y=1.41 $X2=0 $Y2=0
cc_346 N_B2_c_418_n N_VPWR_c_475_n 0.00606499f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_347 N_B2_c_419_n N_VPWR_c_475_n 0.00606499f $X=6.685 $Y=1.41 $X2=0 $Y2=0
cc_348 N_B2_c_420_n N_VPWR_c_475_n 0.00609021f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_349 N_B2_c_412_n N_Y_c_647_n 0.00942464f $X=5.72 $Y=0.995 $X2=0 $Y2=0
cc_350 N_B2_c_413_n N_Y_c_647_n 0.00929111f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_351 N_B2_c_414_n N_Y_c_647_n 0.00955778f $X=6.66 $Y=0.995 $X2=0 $Y2=0
cc_352 N_B2_c_415_n N_Y_c_647_n 0.0105624f $X=7.18 $Y=0.995 $X2=0 $Y2=0
cc_353 B2 N_Y_c_647_n 0.0677865f $X=6.825 $Y=1.105 $X2=0 $Y2=0
cc_354 N_B2_c_416_n N_Y_c_647_n 0.0109421f $X=7.155 $Y=1.202 $X2=0 $Y2=0
cc_355 N_B2_c_418_n N_Y_c_686_n 0.0108425f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_356 N_B2_c_419_n N_Y_c_686_n 0.0108425f $X=6.685 $Y=1.41 $X2=0 $Y2=0
cc_357 N_B2_c_420_n N_Y_c_650_n 0.0108425f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_358 N_B2_c_417_n N_A_885_297#_c_778_n 0.0143148f $X=5.745 $Y=1.41 $X2=0 $Y2=0
cc_359 N_B2_c_418_n N_A_885_297#_c_778_n 0.0100164f $X=6.215 $Y=1.41 $X2=0 $Y2=0
cc_360 N_B2_c_419_n N_A_885_297#_c_780_n 0.0099733f $X=6.685 $Y=1.41 $X2=0 $Y2=0
cc_361 N_B2_c_420_n N_A_885_297#_c_780_n 0.0099733f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_362 N_B2_c_412_n N_A_33_47#_c_824_n 0.00886996f $X=5.72 $Y=0.995 $X2=0 $Y2=0
cc_363 N_B2_c_413_n N_A_33_47#_c_824_n 0.00931157f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_364 N_B2_c_414_n N_A_33_47#_c_824_n 0.00931157f $X=6.66 $Y=0.995 $X2=0 $Y2=0
cc_365 N_B2_c_415_n N_A_33_47#_c_824_n 0.00923997f $X=7.18 $Y=0.995 $X2=0 $Y2=0
cc_366 N_B2_c_412_n N_VGND_c_947_n 0.00357877f $X=5.72 $Y=0.995 $X2=0 $Y2=0
cc_367 N_B2_c_413_n N_VGND_c_947_n 0.00357877f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_368 N_B2_c_414_n N_VGND_c_947_n 0.00357877f $X=6.66 $Y=0.995 $X2=0 $Y2=0
cc_369 N_B2_c_415_n N_VGND_c_947_n 0.00357877f $X=7.18 $Y=0.995 $X2=0 $Y2=0
cc_370 N_B2_c_412_n N_VGND_c_948_n 0.00538038f $X=5.72 $Y=0.995 $X2=0 $Y2=0
cc_371 N_B2_c_413_n N_VGND_c_948_n 0.00548399f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_372 N_B2_c_414_n N_VGND_c_948_n 0.00559933f $X=6.66 $Y=0.995 $X2=0 $Y2=0
cc_373 N_B2_c_415_n N_VGND_c_948_n 0.00561849f $X=7.18 $Y=0.995 $X2=0 $Y2=0
cc_374 N_VPWR_c_475_n N_A_123_297#_M1007_d 0.0031047f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_375 N_VPWR_c_475_n N_A_123_297#_M1012_d 0.00241848f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_475_n N_A_123_297#_M1015_s 0.00229658f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_475_n N_A_123_297#_M1025_s 0.0023046f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_477_n N_A_123_297#_c_591_n 0.00259649f $X=0.29 $Y=1.62 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_478_n N_A_123_297#_c_617_n 0.0149311f $X=1.105 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_475_n N_A_123_297#_c_617_n 0.00955092f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_M1011_s N_A_123_297#_c_601_n 0.00409206f $X=1.085 $Y=1.485 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_479_n N_A_123_297#_c_601_n 0.0139109f $X=1.23 $Y=2.3 $X2=0 $Y2=0
cc_383 N_VPWR_c_475_n N_A_123_297#_c_601_n 0.0141598f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_484_n N_A_123_297#_c_608_n 0.0400924f $X=3.965 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_475_n N_A_123_297#_c_608_n 0.0253962f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_484_n N_A_123_297#_c_624_n 0.0134783f $X=3.965 $Y=2.72 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_475_n N_A_123_297#_c_624_n 0.00808747f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_484_n N_A_123_297#_c_610_n 0.0386815f $X=3.965 $Y=2.72 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_475_n N_A_123_297#_c_610_n 0.0239224f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_484_n N_A_123_297#_c_628_n 0.014332f $X=3.965 $Y=2.72 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_475_n N_A_123_297#_c_628_n 0.00938745f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_480_n N_A_123_297#_c_607_n 0.0207828f $X=4.09 $Y=2.3 $X2=0 $Y2=0
cc_393 N_VPWR_c_484_n N_A_123_297#_c_607_n 0.0162495f $X=3.965 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_475_n N_A_123_297#_c_607_n 0.0107392f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_475_n N_Y_M1000_d 0.00232092f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_396 N_VPWR_c_475_n N_Y_M1022_d 0.00231289f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_c_475_n N_Y_M1001_d 0.00232092f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_c_475_n N_Y_M1013_d 0.00231289f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_c_475_n N_Y_c_654_n 0.00153883f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_400 N_VPWR_c_475_n N_Y_c_686_n 0.00153883f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_M1030_s N_Y_c_650_n 0.00710404f $X=7.715 $Y=1.485 $X2=0 $Y2=0
cc_402 N_VPWR_c_482_n N_Y_c_650_n 0.00245087f $X=7.875 $Y=2.635 $X2=0 $Y2=0
cc_403 N_VPWR_c_483_n N_Y_c_650_n 0.0200542f $X=7.86 $Y=2.3 $X2=0 $Y2=0
cc_404 N_VPWR_c_475_n N_Y_c_650_n 0.0130164f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_M1030_s N_Y_c_648_n 0.00449515f $X=7.715 $Y=1.485 $X2=0 $Y2=0
cc_406 N_VPWR_M1027_s N_Y_c_659_n 0.00903367f $X=3.905 $Y=1.485 $X2=0 $Y2=0
cc_407 N_VPWR_c_480_n N_Y_c_659_n 0.0172305f $X=4.09 $Y=2.3 $X2=0 $Y2=0
cc_408 N_VPWR_c_475_n N_Y_c_659_n 0.0145575f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_c_475_n N_A_885_297#_M1003_d 0.00227246f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_410 N_VPWR_c_475_n N_A_885_297#_M1023_d 0.00241844f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_475_n N_A_885_297#_M1008_s 0.00229658f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_475_n N_A_885_297#_M1028_s 0.00241598f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_M1018_s N_A_885_297#_c_770_n 0.00347905f $X=4.895 $Y=1.485 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_481_n N_A_885_297#_c_770_n 0.0139109f $X=5.04 $Y=2.3 $X2=0 $Y2=0
cc_415 N_VPWR_c_475_n N_A_885_297#_c_770_n 0.0139702f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_488_n N_A_885_297#_c_778_n 0.0386815f $X=7.735 $Y=2.72 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_475_n N_A_885_297#_c_778_n 0.0239144f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_488_n N_A_885_297#_c_791_n 0.015002f $X=7.735 $Y=2.72 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_475_n N_A_885_297#_c_791_n 0.00962794f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_488_n N_A_885_297#_c_780_n 0.0386815f $X=7.735 $Y=2.72 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_475_n N_A_885_297#_c_780_n 0.0239224f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_480_n N_A_885_297#_c_776_n 0.0257341f $X=4.09 $Y=2.3 $X2=0 $Y2=0
cc_423 N_VPWR_c_486_n N_A_885_297#_c_776_n 0.0204601f $X=4.925 $Y=2.72 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_475_n N_A_885_297#_c_776_n 0.0130874f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_488_n N_A_885_297#_c_798_n 0.014332f $X=7.735 $Y=2.72 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_475_n N_A_885_297#_c_798_n 0.00938745f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_488_n N_A_885_297#_c_800_n 0.0143076f $X=7.735 $Y=2.72 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_475_n N_A_885_297#_c_800_n 0.00938089f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_429 N_A_123_297#_c_608_n N_Y_M1000_d 0.00352392f $X=2.515 $Y=2.38 $X2=0 $Y2=0
cc_430 N_A_123_297#_c_610_n N_Y_M1022_d 0.00352392f $X=3.455 $Y=2.38 $X2=0 $Y2=0
cc_431 N_A_123_297#_M1015_s N_Y_c_654_n 0.00347905f $X=2.495 $Y=1.485 $X2=0
+ $Y2=0
cc_432 N_A_123_297#_c_608_n N_Y_c_654_n 0.00608347f $X=2.515 $Y=2.38 $X2=0 $Y2=0
cc_433 N_A_123_297#_c_610_n N_Y_c_654_n 0.00608347f $X=3.455 $Y=2.38 $X2=0 $Y2=0
cc_434 N_A_123_297#_c_628_n N_Y_c_654_n 0.0131392f $X=2.64 $Y=2.3 $X2=0 $Y2=0
cc_435 N_A_123_297#_c_601_n N_Y_c_658_n 0.0140678f $X=1.575 $Y=1.87 $X2=0 $Y2=0
cc_436 N_A_123_297#_c_640_p N_Y_c_658_n 0.0127426f $X=1.7 $Y=1.96 $X2=0 $Y2=0
cc_437 N_A_123_297#_c_608_n N_Y_c_658_n 0.0173581f $X=2.515 $Y=2.38 $X2=0 $Y2=0
cc_438 N_A_123_297#_M1025_s N_Y_c_659_n 0.00367036f $X=3.435 $Y=1.485 $X2=0
+ $Y2=0
cc_439 N_A_123_297#_c_610_n N_Y_c_659_n 0.00608347f $X=3.455 $Y=2.38 $X2=0 $Y2=0
cc_440 N_A_123_297#_c_607_n N_Y_c_659_n 0.0143527f $X=3.58 $Y=2.3 $X2=0 $Y2=0
cc_441 N_A_123_297#_c_610_n Y 0.0127274f $X=3.455 $Y=2.38 $X2=0 $Y2=0
cc_442 N_Y_c_646_n N_A_885_297#_M1003_d 0.00252049f $X=4.465 $Y=1.445 $X2=-0.19
+ $Y2=-0.24
cc_443 N_Y_c_686_n N_A_885_297#_M1008_s 0.00347905f $X=6.795 $Y=1.87 $X2=0 $Y2=0
cc_444 N_Y_c_650_n N_A_885_297#_M1028_s 0.00372618f $X=7.905 $Y=1.87 $X2=0 $Y2=0
cc_445 N_Y_c_646_n N_A_885_297#_c_774_n 0.00284755f $X=4.465 $Y=1.445 $X2=0
+ $Y2=0
cc_446 N_Y_c_659_n N_A_885_297#_c_774_n 0.0148586f $X=4.2 $Y=1.87 $X2=0 $Y2=0
cc_447 N_Y_M1001_d N_A_885_297#_c_778_n 0.00352392f $X=5.835 $Y=1.485 $X2=0
+ $Y2=0
cc_448 N_Y_c_686_n N_A_885_297#_c_778_n 0.00608347f $X=6.795 $Y=1.87 $X2=0 $Y2=0
cc_449 N_Y_c_694_n N_A_885_297#_c_778_n 0.0127274f $X=5.98 $Y=1.87 $X2=0 $Y2=0
cc_450 N_Y_M1013_d N_A_885_297#_c_780_n 0.00352392f $X=6.775 $Y=1.485 $X2=0
+ $Y2=0
cc_451 N_Y_c_686_n N_A_885_297#_c_780_n 0.00608347f $X=6.795 $Y=1.87 $X2=0 $Y2=0
cc_452 N_Y_c_650_n N_A_885_297#_c_780_n 0.00608347f $X=7.905 $Y=1.87 $X2=0 $Y2=0
cc_453 N_Y_c_695_n N_A_885_297#_c_780_n 0.0127274f $X=6.92 $Y=1.87 $X2=0 $Y2=0
cc_454 N_Y_c_646_n N_A_885_297#_c_776_n 0.0035794f $X=4.465 $Y=1.445 $X2=0 $Y2=0
cc_455 N_Y_c_659_n N_A_885_297#_c_776_n 0.00103696f $X=4.2 $Y=1.87 $X2=0 $Y2=0
cc_456 N_Y_c_686_n N_A_885_297#_c_798_n 0.0131392f $X=6.795 $Y=1.87 $X2=0 $Y2=0
cc_457 N_Y_c_650_n N_A_885_297#_c_800_n 0.0124948f $X=7.905 $Y=1.87 $X2=0 $Y2=0
cc_458 N_Y_c_647_n N_A_33_47#_M1014_s 0.00504965f $X=7.905 $Y=0.732 $X2=0 $Y2=0
cc_459 N_Y_c_647_n N_A_33_47#_M1009_d 0.00434237f $X=7.905 $Y=0.732 $X2=0 $Y2=0
cc_460 N_Y_c_647_n N_A_33_47#_M1017_d 0.00544525f $X=7.905 $Y=0.732 $X2=0 $Y2=0
cc_461 N_Y_c_647_n N_A_33_47#_M1029_s 0.00667482f $X=7.905 $Y=0.732 $X2=0 $Y2=0
cc_462 N_Y_c_648_n N_A_33_47#_M1029_s 0.00104005f $X=8.037 $Y=1.785 $X2=0 $Y2=0
cc_463 N_Y_c_646_n N_A_33_47#_c_823_n 0.00386175f $X=4.465 $Y=1.445 $X2=0 $Y2=0
cc_464 N_Y_M1004_d N_A_33_47#_c_824_n 0.00399124f $X=4.385 $Y=0.235 $X2=0 $Y2=0
cc_465 N_Y_M1020_d N_A_33_47#_c_824_n 0.00312026f $X=5.375 $Y=0.235 $X2=0 $Y2=0
cc_466 N_Y_M1010_s N_A_33_47#_c_824_n 0.00400389f $X=6.265 $Y=0.235 $X2=0 $Y2=0
cc_467 N_Y_M1021_s N_A_33_47#_c_824_n 0.00410384f $X=7.255 $Y=0.235 $X2=0 $Y2=0
cc_468 N_Y_c_671_n N_A_33_47#_c_824_n 0.012594f $X=4.465 $Y=0.82 $X2=0 $Y2=0
cc_469 N_Y_c_647_n N_A_33_47#_c_824_n 0.184537f $X=7.905 $Y=0.732 $X2=0 $Y2=0
cc_470 N_Y_c_647_n N_VGND_c_947_n 0.00248637f $X=7.905 $Y=0.732 $X2=0 $Y2=0
cc_471 N_Y_M1004_d N_VGND_c_948_n 0.00256987f $X=4.385 $Y=0.235 $X2=0 $Y2=0
cc_472 N_Y_M1020_d N_VGND_c_948_n 0.00216833f $X=5.375 $Y=0.235 $X2=0 $Y2=0
cc_473 N_Y_M1010_s N_VGND_c_948_n 0.00256987f $X=6.265 $Y=0.235 $X2=0 $Y2=0
cc_474 N_Y_M1021_s N_VGND_c_948_n 0.00256987f $X=7.255 $Y=0.235 $X2=0 $Y2=0
cc_475 N_Y_c_647_n N_VGND_c_948_n 0.0040842f $X=7.905 $Y=0.732 $X2=0 $Y2=0
cc_476 N_A_33_47#_c_819_n N_VGND_M1005_s 0.00251047f $X=1.015 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_477 N_A_33_47#_c_821_n N_VGND_M1019_s 0.00165819f $X=1.955 $Y=0.82 $X2=0
+ $Y2=0
cc_478 N_A_33_47#_c_822_n N_VGND_M1016_s 0.00251047f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_479 N_A_33_47#_c_823_n N_VGND_M1026_s 0.00255557f $X=3.835 $Y=0.82 $X2=0
+ $Y2=0
cc_480 N_A_33_47#_c_819_n N_VGND_c_937_n 0.0127273f $X=1.015 $Y=0.815 $X2=0
+ $Y2=0
cc_481 N_A_33_47#_c_834_n N_VGND_c_937_n 0.0223967f $X=1.23 $Y=0.39 $X2=0 $Y2=0
cc_482 N_A_33_47#_c_821_n N_VGND_c_938_n 0.0116529f $X=1.955 $Y=0.82 $X2=0 $Y2=0
cc_483 N_A_33_47#_c_839_n N_VGND_c_939_n 0.0183628f $X=2.17 $Y=0.39 $X2=0 $Y2=0
cc_484 N_A_33_47#_c_822_n N_VGND_c_939_n 0.0127273f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_485 N_A_33_47#_c_823_n N_VGND_c_940_n 0.012101f $X=3.835 $Y=0.82 $X2=0 $Y2=0
cc_486 N_A_33_47#_c_844_n N_VGND_c_940_n 0.0172916f $X=4.01 $Y=0.475 $X2=0 $Y2=0
cc_487 N_A_33_47#_c_845_n N_VGND_c_940_n 0.00589622f $X=4.05 $Y=0.73 $X2=0 $Y2=0
cc_488 N_A_33_47#_c_819_n N_VGND_c_941_n 0.00199443f $X=1.015 $Y=0.815 $X2=0
+ $Y2=0
cc_489 N_A_33_47#_c_834_n N_VGND_c_941_n 0.023074f $X=1.23 $Y=0.39 $X2=0 $Y2=0
cc_490 N_A_33_47#_c_821_n N_VGND_c_941_n 0.00248202f $X=1.955 $Y=0.82 $X2=0
+ $Y2=0
cc_491 N_A_33_47#_c_821_n N_VGND_c_943_n 0.00193763f $X=1.955 $Y=0.82 $X2=0
+ $Y2=0
cc_492 N_A_33_47#_c_839_n N_VGND_c_943_n 0.0223596f $X=2.17 $Y=0.39 $X2=0 $Y2=0
cc_493 N_A_33_47#_c_822_n N_VGND_c_943_n 0.00266636f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_494 N_A_33_47#_c_822_n N_VGND_c_945_n 0.00198695f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_495 N_A_33_47#_c_859_n N_VGND_c_945_n 0.0231806f $X=3.11 $Y=0.39 $X2=0 $Y2=0
cc_496 N_A_33_47#_c_823_n N_VGND_c_945_n 0.00248202f $X=3.835 $Y=0.82 $X2=0
+ $Y2=0
cc_497 N_A_33_47#_c_823_n N_VGND_c_947_n 0.00194552f $X=3.835 $Y=0.82 $X2=0
+ $Y2=0
cc_498 N_A_33_47#_c_844_n N_VGND_c_947_n 0.022113f $X=4.01 $Y=0.475 $X2=0 $Y2=0
cc_499 N_A_33_47#_c_824_n N_VGND_c_947_n 0.220057f $X=7.86 $Y=0.39 $X2=0 $Y2=0
cc_500 N_A_33_47#_M1005_d N_VGND_c_948_n 0.00258952f $X=0.165 $Y=0.235 $X2=0
+ $Y2=0
cc_501 N_A_33_47#_M1006_d N_VGND_c_948_n 0.00264276f $X=1.095 $Y=0.235 $X2=0
+ $Y2=0
cc_502 N_A_33_47#_M1002_d N_VGND_c_948_n 0.0025535f $X=1.985 $Y=0.235 $X2=0
+ $Y2=0
cc_503 N_A_33_47#_M1024_d N_VGND_c_948_n 0.00304426f $X=2.925 $Y=0.235 $X2=0
+ $Y2=0
cc_504 N_A_33_47#_M1031_d N_VGND_c_948_n 0.00255355f $X=3.915 $Y=0.235 $X2=0
+ $Y2=0
cc_505 N_A_33_47#_M1014_s N_VGND_c_948_n 0.00295535f $X=4.855 $Y=0.235 $X2=0
+ $Y2=0
cc_506 N_A_33_47#_M1009_d N_VGND_c_948_n 0.00255381f $X=5.795 $Y=0.235 $X2=0
+ $Y2=0
cc_507 N_A_33_47#_M1017_d N_VGND_c_948_n 0.00295535f $X=6.735 $Y=0.235 $X2=0
+ $Y2=0
cc_508 N_A_33_47#_M1029_s N_VGND_c_948_n 0.00209344f $X=7.725 $Y=0.235 $X2=0
+ $Y2=0
cc_509 N_A_33_47#_c_818_n N_VGND_c_948_n 0.0126169f $X=0.29 $Y=0.39 $X2=0 $Y2=0
cc_510 N_A_33_47#_c_819_n N_VGND_c_948_n 0.00977515f $X=1.015 $Y=0.815 $X2=0
+ $Y2=0
cc_511 N_A_33_47#_c_834_n N_VGND_c_948_n 0.0141066f $X=1.23 $Y=0.39 $X2=0 $Y2=0
cc_512 N_A_33_47#_c_821_n N_VGND_c_948_n 0.00938601f $X=1.955 $Y=0.82 $X2=0
+ $Y2=0
cc_513 N_A_33_47#_c_839_n N_VGND_c_948_n 0.0141302f $X=2.17 $Y=0.39 $X2=0 $Y2=0
cc_514 N_A_33_47#_c_822_n N_VGND_c_948_n 0.00972452f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_515 N_A_33_47#_c_859_n N_VGND_c_948_n 0.0143352f $X=3.11 $Y=0.39 $X2=0 $Y2=0
cc_516 N_A_33_47#_c_823_n N_VGND_c_948_n 0.0096764f $X=3.835 $Y=0.82 $X2=0 $Y2=0
cc_517 N_A_33_47#_c_844_n N_VGND_c_948_n 0.013025f $X=4.01 $Y=0.475 $X2=0 $Y2=0
cc_518 N_A_33_47#_c_824_n N_VGND_c_948_n 0.138536f $X=7.86 $Y=0.39 $X2=0 $Y2=0
cc_519 N_A_33_47#_c_818_n N_VGND_c_949_n 0.0217962f $X=0.29 $Y=0.39 $X2=0 $Y2=0
cc_520 N_A_33_47#_c_819_n N_VGND_c_949_n 0.00254521f $X=1.015 $Y=0.815 $X2=0
+ $Y2=0
