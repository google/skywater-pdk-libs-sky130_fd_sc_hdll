* File: sky130_fd_sc_hdll__einvp_2.spice
* Created: Wed Sep  2 08:31:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__einvp_2.pex.spice"
.subckt sky130_fd_sc_hdll__einvp_2  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_TE_M1008_g N_A_27_47#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0843925 AS=0.1092 PD=0.804673 PS=1.36 NRD=21.42 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1008_d N_TE_M1004_g N_A_214_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.130607 AS=0.104 PD=1.24533 PS=0.97 NRD=3.684 NRS=8.304 M=1 R=4.33333
+ SA=75000.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_TE_M1005_g N_A_214_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.195 AS=0.104 PD=1.9 PS=0.97 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_Z_M1000_d N_A_M1000_g N_A_214_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.23075 PD=1.02 PS=2.01 NRD=8.304 NRS=16.608 M=1 R=4.33333
+ SA=75000.3 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_Z_M1000_d N_A_M1006_g N_A_214_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_TE_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1728 AS=0.1728 PD=1.82 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1001 N_VPWR_M1001_d N_A_27_47#_M1001_g N_A_235_309#_M1001_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.2538 PD=1.23 PS=2.42 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90000.2 SB=90001.7 A=0.1692 P=2.24 MULT=1
MM1009 N_VPWR_M1001_d N_A_27_47#_M1009_g N_A_235_309#_M1009_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.210725 PD=1.23 PS=1.39546 NRD=1.0441 NRS=7.3284 M=1
+ R=5.22222 SA=90000.6 SB=90001.3 A=0.1692 P=2.24 MULT=1
MM1003 N_A_235_309#_M1009_s N_A_M1003_g N_Z_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.224175 AS=0.145 PD=1.48454 PS=1.29 NRD=24.6053 NRS=0.9653 M=1 R=5.55556
+ SA=90001.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1007 N_A_235_309#_M1007_d N_A_M1007_g N_Z_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.7 SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_58 VPB 0 1.1096e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__einvp_2.pxi.spice"
*
.ends
*
*
