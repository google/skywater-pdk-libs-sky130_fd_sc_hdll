# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a21bo_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21bo_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.960000 1.010000 5.375000 1.360000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.010000 4.790000 1.275000 ;
        RECT 4.565000 1.275000 4.790000 1.595000 ;
        RECT 4.565000 1.595000 5.860000 1.765000 ;
        RECT 5.630000 1.055000 6.220000 1.290000 ;
        RECT 5.630000 1.290000 5.860000 1.595000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.470000 1.010000 0.850000 1.625000 ;
    END
  END B1_N
  PIN VGND
    ANTENNADIFFAREA  1.423500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.470000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  1.029000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.615000 2.510000 0.785000 ;
        RECT 1.050000 0.785000 1.540000 1.595000 ;
        RECT 1.050000 1.595000 2.580000 1.765000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.105000  0.255000 0.510000 0.840000 ;
      RECT 0.105000  0.840000 0.300000 1.795000 ;
      RECT 0.105000  1.795000 0.535000 1.935000 ;
      RECT 0.105000  1.935000 3.090000 2.105000 ;
      RECT 0.105000  2.105000 0.520000 2.465000 ;
      RECT 0.680000  0.085000 1.070000 0.445000 ;
      RECT 0.690000  2.275000 1.070000 2.635000 ;
      RECT 1.650000  0.085000 2.030000 0.445000 ;
      RECT 1.650000  2.275000 2.030000 2.635000 ;
      RECT 1.710000  0.995000 3.030000 1.185000 ;
      RECT 1.710000  1.185000 2.750000 1.325000 ;
      RECT 2.605000  2.275000 2.990000 2.635000 ;
      RECT 2.735000  0.085000 3.505000 0.445000 ;
      RECT 2.860000  0.615000 3.915000 0.670000 ;
      RECT 2.860000  0.670000 5.385000 0.785000 ;
      RECT 2.860000  0.785000 3.030000 0.995000 ;
      RECT 2.920000  1.355000 3.525000 1.525000 ;
      RECT 2.920000  1.525000 3.090000 1.935000 ;
      RECT 3.215000  0.995000 3.525000 1.355000 ;
      RECT 3.275000  1.695000 3.445000 2.210000 ;
      RECT 3.275000  2.210000 4.385000 2.380000 ;
      RECT 3.745000  0.255000 3.915000 0.615000 ;
      RECT 3.745000  0.785000 5.385000 0.840000 ;
      RECT 3.745000  0.840000 3.915000 1.805000 ;
      RECT 4.175000  0.085000 4.505000 0.445000 ;
      RECT 4.205000  1.445000 4.385000 1.935000 ;
      RECT 4.205000  1.935000 6.345000 2.105000 ;
      RECT 4.205000  2.105000 4.385000 2.210000 ;
      RECT 4.555000  2.275000 4.935000 2.635000 ;
      RECT 5.105000  0.405000 5.385000 0.670000 ;
      RECT 5.495000  2.275000 5.875000 2.635000 ;
      RECT 6.065000  0.085000 6.345000 0.885000 ;
      RECT 6.090000  1.460000 6.345000 1.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21bo_4
