* File: sky130_fd_sc_hdll__a221oi_4.spice
* Created: Thu Aug 27 18:53:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a221oi_4.pex.spice"
.subckt sky130_fd_sc_hdll__a221oi_4  VNB VPB C1 B2 B1 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_C1_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.2145 PD=0.97 PS=1.96 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.3 SB=75009.7
+ A=0.0975 P=1.6 MULT=1
MM1020 N_Y_M1007_d N_C1_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7 SB=75009.2
+ A=0.0975 P=1.6 MULT=1
MM1024 N_Y_M1024_d N_C1_M1024_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2 SB=75008.8
+ A=0.0975 P=1.6 MULT=1
MM1033 N_Y_M1024_d N_C1_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.1105 PD=0.97 PS=0.99 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7 SB=75008.3
+ A=0.0975 P=1.6 MULT=1
MM1001 N_A_503_47#_M1001_d N_B2_M1001_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.1105 PD=0.97 PS=0.99 NRD=0 NRS=11.988 M=1 R=4.33333 SA=75002.2
+ SB=75007.8 A=0.0975 P=1.6 MULT=1
MM1015 N_A_503_47#_M1001_d N_B2_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75007.3 A=0.0975 P=1.6 MULT=1
MM1027 N_A_503_47#_M1027_d N_B2_M1027_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2665 AS=0.104 PD=1.47 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.1
+ SB=75006.9 A=0.0975 P=1.6 MULT=1
MM1021 N_A_503_47#_M1027_d N_B1_M1021_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2665 AS=0.104 PD=1.47 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.1
+ SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1022 N_A_503_47#_M1022_d N_B1_M1022_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1029 N_A_503_47#_M1022_d N_B1_M1029_g N_Y_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1038 N_A_503_47#_M1038_d N_B1_M1038_g N_Y_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.5
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1036 N_A_503_47#_M1038_d N_B2_M1036_g N_VGND_M1036_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333 SA=75006
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1006 N_A_1375_47#_M1006_d N_A2_M1006_g N_VGND_M1036_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.5
+ SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1002 N_A_1375_47#_M1006_d N_A1_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.9
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1011 N_A_1375_47#_M1011_d N_A1_M1011_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75007.4
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1017 N_A_1375_47#_M1011_d N_A1_M1017_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75007.9
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1039 N_A_1375_47#_M1039_d N_A1_M1039_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75008.4
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1009 N_A_1375_47#_M1039_d N_A2_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75008.8
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1025 N_A_1375_47#_M1025_d N_A2_M1025_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75009.3
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1037 N_A_1375_47#_M1025_d N_A2_M1037_g N_VGND_M1037_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.18525 PD=0.97 PS=1.87 NRD=0 NRS=0 M=1 R=4.33333 SA=75009.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1010 N_Y_M1003_d N_C1_M1010_g N_A_27_297#_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1016 N_Y_M1016_d N_C1_M1016_g N_A_27_297#_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1028 N_Y_M1016_d N_C1_M1028_g N_A_27_297#_M1028_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1014 N_A_511_297#_M1014_d N_B2_M1014_g N_A_27_297#_M1014_s VPB PHIGHVT L=0.18
+ W=1 AD=0.32 AS=0.145 PD=2.64 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90007.3 A=0.18 P=2.36 MULT=1
MM1018 N_A_511_297#_M1018_d N_B2_M1018_g N_A_27_297#_M1014_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90006.8 A=0.18 P=2.36 MULT=1
MM1030 N_A_511_297#_M1018_d N_B2_M1030_g N_A_27_297#_M1030_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.2 SB=90006.4 A=0.18 P=2.36 MULT=1
MM1004 N_A_27_297#_M1030_s N_B1_M1004_g N_A_511_297#_M1004_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90005.9 A=0.18 P=2.36 MULT=1
MM1012 N_A_27_297#_M1012_d N_B1_M1012_g N_A_511_297#_M1004_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90005.4 A=0.18 P=2.36 MULT=1
MM1026 N_A_27_297#_M1012_d N_B1_M1026_g N_A_511_297#_M1026_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1032 N_A_27_297#_M1032_d N_B1_M1032_g N_A_511_297#_M1026_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003 SB=90004.5 A=0.18 P=2.36 MULT=1
MM1034 N_A_511_297#_M1034_d N_B2_M1034_g N_A_27_297#_M1032_d VPB PHIGHVT L=0.18
+ W=1 AD=0.17 AS=0.145 PD=1.34 PS=1.29 NRD=8.8453 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90004 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_511_297#_M1034_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.17 PD=1.29 PS=1.34 NRD=0.9653 NRS=2.9353 M=1 R=5.55556 SA=90004
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1000 N_A_511_297#_M1000_d N_A1_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.5 SB=90003 A=0.18 P=2.36 MULT=1
MM1019 N_A_511_297#_M1000_d N_A1_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1031 N_A_511_297#_M1031_d N_A1_M1031_g N_VPWR_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.4 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1035 N_A_511_297#_M1031_d N_A1_M1035_g N_VPWR_M1035_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.9 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1035_s N_A2_M1008_g N_A_511_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.4 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A2_M1013_g N_A_511_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.9 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1013_d N_A2_M1023_g N_A_511_297#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX40_noxref VNB VPB NWDIODE A=17.5908 P=25.13
pX41_noxref noxref_15 A2 A2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a221oi_4.pxi.spice"
*
.ends
*
*
