# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xnor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xnor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.495000 1.075000 8.215000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.625000 0.995000 6.845000 1.445000 ;
        RECT 6.625000 1.445000 7.255000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715000 1.075000 2.330000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.472000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.345000 1.440000 ;
        RECT 0.085000 1.440000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.200000 0.085000 ;
        RECT 0.515000  0.085000 0.815000 0.525000 ;
        RECT 3.675000  0.085000 3.845000 0.865000 ;
        RECT 8.050000  0.085000 8.510000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.200000 2.805000 ;
        RECT 0.535000 2.215000 0.920000 2.635000 ;
        RECT 3.425000 2.235000 3.755000 2.635000 ;
        RECT 7.915000 2.275000 8.595000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515000 0.695000 1.205000 0.865000 ;
      RECT 0.515000 0.865000 0.755000 1.330000 ;
      RECT 0.535000 1.330000 0.755000 1.875000 ;
      RECT 0.535000 1.875000 1.320000 2.045000 ;
      RECT 0.985000 0.255000 2.655000 0.425000 ;
      RECT 0.985000 0.425000 1.205000 0.695000 ;
      RECT 0.985000 1.535000 2.670000 1.705000 ;
      RECT 1.100000 2.045000 1.320000 2.235000 ;
      RECT 1.100000 2.235000 2.670000 2.405000 ;
      RECT 1.375000 0.595000 1.545000 1.535000 ;
      RECT 1.660000 1.895000 4.360000 2.065000 ;
      RECT 1.845000 0.625000 3.165000 0.795000 ;
      RECT 1.845000 0.795000 2.225000 0.905000 ;
      RECT 2.170000 0.425000 2.655000 0.455000 ;
      RECT 2.500000 0.995000 2.825000 1.325000 ;
      RECT 2.500000 1.325000 2.670000 1.535000 ;
      RECT 2.875000 0.285000 3.505000 0.455000 ;
      RECT 2.890000 1.525000 3.275000 1.695000 ;
      RECT 2.995000 0.795000 3.165000 1.375000 ;
      RECT 2.995000 1.375000 3.275000 1.525000 ;
      RECT 3.335000 0.455000 3.505000 1.035000 ;
      RECT 3.335000 1.035000 3.615000 1.205000 ;
      RECT 3.445000 1.205000 3.615000 1.895000 ;
      RECT 3.845000 1.445000 4.365000 1.715000 ;
      RECT 4.075000 0.415000 4.365000 1.445000 ;
      RECT 4.190000 2.065000 4.360000 2.275000 ;
      RECT 4.190000 2.275000 7.485000 2.445000 ;
      RECT 4.545000 0.265000 4.955000 0.485000 ;
      RECT 4.545000 0.485000 4.755000 0.595000 ;
      RECT 4.545000 0.595000 4.715000 2.105000 ;
      RECT 4.885000 0.720000 5.345000 0.825000 ;
      RECT 4.885000 0.825000 5.145000 0.890000 ;
      RECT 4.885000 0.890000 5.055000 2.275000 ;
      RECT 4.925000 0.655000 5.345000 0.720000 ;
      RECT 5.175000 0.320000 5.345000 0.655000 ;
      RECT 5.285000 1.445000 6.115000 1.615000 ;
      RECT 5.285000 1.615000 5.700000 2.045000 ;
      RECT 5.300000 0.995000 5.725000 1.270000 ;
      RECT 5.515000 0.630000 5.725000 0.995000 ;
      RECT 5.945000 0.255000 7.140000 0.425000 ;
      RECT 5.945000 0.425000 6.115000 1.445000 ;
      RECT 6.285000 0.595000 6.455000 1.935000 ;
      RECT 6.285000 1.935000 9.110000 2.105000 ;
      RECT 6.625000 0.425000 7.140000 0.465000 ;
      RECT 7.015000 0.730000 7.220000 0.945000 ;
      RECT 7.015000 0.945000 7.325000 1.275000 ;
      RECT 7.475000 1.495000 8.660000 1.705000 ;
      RECT 7.515000 0.295000 7.805000 0.735000 ;
      RECT 7.515000 0.735000 8.660000 0.750000 ;
      RECT 7.555000 0.750000 8.660000 0.905000 ;
      RECT 8.490000 0.905000 8.660000 0.995000 ;
      RECT 8.490000 0.995000 8.770000 1.325000 ;
      RECT 8.490000 1.325000 8.660000 1.495000 ;
      RECT 8.575000 1.875000 9.110000 1.935000 ;
      RECT 8.810000 0.255000 9.110000 0.585000 ;
      RECT 8.815000 2.105000 9.110000 2.465000 ;
      RECT 8.940000 0.585000 9.110000 1.875000 ;
    LAYER mcon ;
      RECT 3.105000 1.445000 3.275000 1.615000 ;
      RECT 4.075000 0.765000 4.245000 0.935000 ;
      RECT 4.585000 0.425000 4.755000 0.595000 ;
      RECT 5.555000 0.765000 5.725000 0.935000 ;
      RECT 5.555000 1.445000 5.725000 1.615000 ;
      RECT 7.035000 0.765000 7.205000 0.935000 ;
      RECT 7.545000 0.425000 7.715000 0.595000 ;
    LAYER met1 ;
      RECT 3.045000 1.415000 3.335000 1.460000 ;
      RECT 3.045000 1.460000 5.785000 1.600000 ;
      RECT 3.045000 1.600000 3.335000 1.645000 ;
      RECT 4.015000 0.735000 4.305000 0.780000 ;
      RECT 4.015000 0.780000 7.265000 0.920000 ;
      RECT 4.015000 0.920000 4.305000 0.965000 ;
      RECT 4.525000 0.395000 4.815000 0.440000 ;
      RECT 4.525000 0.440000 7.775000 0.580000 ;
      RECT 4.525000 0.580000 4.815000 0.625000 ;
      RECT 5.495000 0.735000 5.785000 0.780000 ;
      RECT 5.495000 0.920000 5.785000 0.965000 ;
      RECT 5.495000 1.415000 5.785000 1.460000 ;
      RECT 5.495000 1.600000 5.785000 1.645000 ;
      RECT 6.975000 0.735000 7.265000 0.780000 ;
      RECT 6.975000 0.920000 7.265000 0.965000 ;
      RECT 7.485000 0.395000 7.775000 0.440000 ;
      RECT 7.485000 0.580000 7.775000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor3_1
