# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xor2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.04000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 3.100000 1.275000 ;
        RECT 2.880000 1.275000 3.100000 1.445000 ;
        RECT 2.880000 1.445000 6.815000 1.615000 ;
        RECT 6.595000 1.075000 8.120000 1.275000 ;
        RECT 6.595000 1.275000 6.815000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 1.075000 5.500000 1.105000 ;
        RECT 3.270000 1.105000 6.340000 1.275000 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  1.318500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.650000 0.725000  9.480000 0.735000 ;
        RECT  8.650000 0.735000 10.955000 0.905000 ;
        RECT  8.680000 1.445000 10.955000 1.625000 ;
        RECT  8.680000 1.625000  9.910000 1.665000 ;
        RECT  8.680000 1.665000  8.970000 2.125000 ;
        RECT  9.100000 0.255000  9.480000 0.725000 ;
        RECT  9.660000 1.665000  9.910000 2.125000 ;
        RECT 10.040000 0.255000 10.420000 0.735000 ;
        RECT 10.550000 1.625000 10.955000 2.465000 ;
        RECT 10.635000 0.905000 10.955000 1.445000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.085000  0.085000  0.360000 0.565000 ;
      RECT  0.085000  0.735000  3.730000 0.905000 ;
      RECT  0.085000  0.905000  0.255000 1.445000 ;
      RECT  0.085000  1.445000  2.670000 1.615000 ;
      RECT  0.085000  1.785000  2.280000 2.005000 ;
      RECT  0.085000  2.005000  0.400000 2.465000 ;
      RECT  0.530000  0.255000  0.910000 0.725000 ;
      RECT  0.530000  0.725000  3.730000 0.735000 ;
      RECT  0.620000  2.175000  0.870000 2.635000 ;
      RECT  1.090000  2.005000  1.340000 2.465000 ;
      RECT  1.130000  0.085000  1.300000 0.555000 ;
      RECT  1.470000  0.255000  1.850000 0.725000 ;
      RECT  1.560000  2.175000  1.810000 2.635000 ;
      RECT  2.030000  2.005000  2.280000 2.295000 ;
      RECT  2.030000  2.295000  4.160000 2.465000 ;
      RECT  2.070000  0.085000  2.240000 0.555000 ;
      RECT  2.410000  0.255000  2.790000 0.725000 ;
      RECT  2.500000  1.615000  2.670000 1.785000 ;
      RECT  2.500000  1.785000  3.690000 1.955000 ;
      RECT  2.500000  1.955000  2.750000 2.125000 ;
      RECT  2.970000  2.125000  3.220000 2.295000 ;
      RECT  3.010000  0.085000  3.180000 0.555000 ;
      RECT  3.350000  0.255000  3.730000 0.725000 ;
      RECT  3.440000  1.955000  3.690000 2.125000 ;
      RECT  3.910000  1.795000  4.160000 2.295000 ;
      RECT  3.950000  0.085000  4.220000 0.895000 ;
      RECT  4.390000  0.255000  6.600000 0.475000 ;
      RECT  4.430000  1.785000  8.440000 2.005000 ;
      RECT  4.430000  2.005000  4.680000 2.465000 ;
      RECT  4.565000  0.645000  6.130000 0.905000 ;
      RECT  4.900000  2.175000  5.150000 2.635000 ;
      RECT  5.370000  2.005000  5.620000 2.465000 ;
      RECT  5.650000  0.905000  6.130000 0.935000 ;
      RECT  5.840000  2.175000  6.090000 2.635000 ;
      RECT  6.310000  2.005000  6.560000 2.465000 ;
      RECT  6.350000  0.475000  6.600000 0.725000 ;
      RECT  6.350000  0.725000  8.480000 0.905000 ;
      RECT  6.780000  2.175000  7.030000 2.635000 ;
      RECT  6.820000  0.085000  6.990000 0.555000 ;
      RECT  7.160000  0.255000  7.540000 0.725000 ;
      RECT  7.250000  1.455000  7.500000 1.785000 ;
      RECT  7.250000  2.005000  7.500000 2.465000 ;
      RECT  7.720000  2.175000  7.970000 2.635000 ;
      RECT  7.760000  0.085000  7.930000 0.555000 ;
      RECT  8.010000  1.445000  8.510000 1.615000 ;
      RECT  8.100000  0.255000  8.480000 0.725000 ;
      RECT  8.190000  2.005000  8.440000 2.295000 ;
      RECT  8.190000  2.295000 10.380000 2.465000 ;
      RECT  8.340000  1.075000 10.130000 1.275000 ;
      RECT  8.340000  1.275000  8.510000 1.445000 ;
      RECT  8.760000  0.085000  8.930000 0.555000 ;
      RECT  9.190000  1.835000  9.440000 2.295000 ;
      RECT  9.700000  0.085000  9.870000 0.555000 ;
      RECT 10.130000  1.795000 10.380000 2.295000 ;
      RECT 10.640000  0.085000 10.810000 0.555000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.185000  1.445000  2.355000 1.615000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.705000  0.725000  5.875000 0.895000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.305000  1.445000  8.475000 1.615000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.765000  0.725000  8.935000 0.895000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 2.125000 1.415000 2.415000 1.460000 ;
      RECT 2.125000 1.460000 8.535000 1.600000 ;
      RECT 2.125000 1.600000 2.415000 1.645000 ;
      RECT 5.645000 0.695000 5.935000 0.780000 ;
      RECT 5.645000 0.780000 8.995000 0.925000 ;
      RECT 8.245000 1.415000 8.535000 1.460000 ;
      RECT 8.245000 1.600000 8.535000 1.645000 ;
      RECT 8.705000 0.695000 8.995000 0.780000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor2_4
END LIBRARY
