# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.005000 1.075000 8.695000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.085000 0.995000 7.305000 1.445000 ;
        RECT 7.085000 1.445000 7.715000 1.725000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 0.995000 2.645000 1.325000 ;
    END
  END C
  PIN VGND
    ANTENNADIFFAREA  0.970950 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.309400 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.472000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.590000 0.925000 ;
        RECT 0.085000 0.925000 0.400000 1.440000 ;
        RECT 0.085000 1.440000 0.610000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.800000  0.695000 1.450000 0.865000 ;
      RECT 0.800000  0.865000 1.000000 1.875000 ;
      RECT 0.800000  1.875000 1.570000 2.045000 ;
      RECT 0.810000  0.085000 1.060000 0.525000 ;
      RECT 0.830000  2.215000 1.165000 2.635000 ;
      RECT 1.230000  0.255000 2.890000 0.425000 ;
      RECT 1.230000  0.425000 1.450000 0.695000 ;
      RECT 1.235000  1.535000 2.985000 1.705000 ;
      RECT 1.350000  2.045000 1.570000 2.235000 ;
      RECT 1.350000  2.235000 3.045000 2.405000 ;
      RECT 1.620000  0.595000 1.790000 1.535000 ;
      RECT 1.970000  1.895000 3.375000 2.065000 ;
      RECT 2.070000  0.655000 3.280000 0.825000 ;
      RECT 2.490000  0.425000 2.890000 0.455000 ;
      RECT 2.815000  0.995000 3.140000 1.325000 ;
      RECT 2.815000  1.325000 2.985000 1.535000 ;
      RECT 3.060000  0.255000 3.960000 0.425000 ;
      RECT 3.060000  0.425000 3.280000 0.655000 ;
      RECT 3.205000  1.525000 3.735000 1.695000 ;
      RECT 3.205000  1.695000 3.375000 1.895000 ;
      RECT 3.310000  2.235000 3.715000 2.405000 ;
      RECT 3.450000  0.595000 3.620000 1.375000 ;
      RECT 3.450000  1.375000 3.735000 1.525000 ;
      RECT 3.545000  1.895000 4.820000 2.065000 ;
      RECT 3.545000  2.065000 3.715000 2.235000 ;
      RECT 3.790000  0.425000 3.960000 1.035000 ;
      RECT 3.790000  1.035000 4.075000 1.205000 ;
      RECT 3.885000  2.235000 4.215000 2.635000 ;
      RECT 3.905000  1.205000 4.075000 1.895000 ;
      RECT 4.130000  0.085000 4.300000 0.865000 ;
      RECT 4.305000  1.445000 4.820000 1.715000 ;
      RECT 4.530000  0.415000 4.820000 1.445000 ;
      RECT 4.650000  2.065000 4.820000 2.275000 ;
      RECT 4.650000  2.275000 7.945000 2.445000 ;
      RECT 4.995000  0.265000 5.410000 0.485000 ;
      RECT 4.995000  0.485000 5.215000 0.595000 ;
      RECT 4.995000  0.595000 5.165000 2.105000 ;
      RECT 5.335000  0.720000 5.800000 0.825000 ;
      RECT 5.335000  0.825000 5.605000 0.890000 ;
      RECT 5.335000  0.890000 5.505000 2.275000 ;
      RECT 5.385000  0.655000 5.800000 0.720000 ;
      RECT 5.630000  0.320000 5.800000 0.655000 ;
      RECT 5.745000  1.445000 6.575000 1.615000 ;
      RECT 5.745000  1.615000 6.160000 2.045000 ;
      RECT 5.760000  0.995000 6.185000 1.270000 ;
      RECT 5.970000  0.630000 6.185000 0.995000 ;
      RECT 6.405000  0.255000 7.600000 0.425000 ;
      RECT 6.405000  0.425000 6.575000 1.445000 ;
      RECT 6.745000  0.595000 6.915000 1.935000 ;
      RECT 6.745000  1.935000 9.565000 2.105000 ;
      RECT 7.085000  0.425000 7.600000 0.465000 ;
      RECT 7.475000  0.730000 7.680000 0.945000 ;
      RECT 7.475000  0.945000 7.785000 1.275000 ;
      RECT 7.935000  1.495000 9.115000 1.705000 ;
      RECT 7.975000  0.295000 8.265000 0.735000 ;
      RECT 7.975000  0.735000 9.115000 0.750000 ;
      RECT 8.015000  0.750000 9.115000 0.905000 ;
      RECT 8.355000  2.275000 9.050000 2.635000 ;
      RECT 8.485000  0.085000 8.935000 0.565000 ;
      RECT 8.945000  0.905000 9.115000 0.995000 ;
      RECT 8.945000  0.995000 9.225000 1.325000 ;
      RECT 8.945000  1.325000 9.115000 1.495000 ;
      RECT 9.030000  1.875000 9.565000 1.935000 ;
      RECT 9.265000  0.255000 9.565000 0.585000 ;
      RECT 9.270000  2.105000 9.565000 2.465000 ;
      RECT 9.395000  0.585000 9.565000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.565000  1.445000 3.735000 1.615000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.535000  0.765000 4.705000 0.935000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.045000  0.425000 5.215000 0.595000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.015000  0.765000 6.185000 0.935000 ;
      RECT 6.015000  1.445000 6.185000 1.615000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.495000  0.765000 7.665000 0.935000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.005000  0.425000 8.175000 0.595000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 3.505000 1.415000 3.795000 1.460000 ;
      RECT 3.505000 1.460000 6.245000 1.600000 ;
      RECT 3.505000 1.600000 3.795000 1.645000 ;
      RECT 4.475000 0.735000 4.765000 0.780000 ;
      RECT 4.475000 0.780000 7.725000 0.920000 ;
      RECT 4.475000 0.920000 4.765000 0.965000 ;
      RECT 4.985000 0.395000 5.275000 0.440000 ;
      RECT 4.985000 0.440000 8.235000 0.580000 ;
      RECT 4.985000 0.580000 5.275000 0.625000 ;
      RECT 5.955000 0.735000 6.245000 0.780000 ;
      RECT 5.955000 0.920000 6.245000 0.965000 ;
      RECT 5.955000 1.415000 6.245000 1.460000 ;
      RECT 5.955000 1.600000 6.245000 1.645000 ;
      RECT 7.435000 0.735000 7.725000 0.780000 ;
      RECT 7.435000 0.920000 7.725000 0.965000 ;
      RECT 7.945000 0.395000 8.235000 0.440000 ;
      RECT 7.945000 0.580000 8.235000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor3_1
