* File: sky130_fd_sc_hdll__and4b_4.pxi.spice
* Created: Wed Sep  2 08:23:27 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND4B_4%A_N N_A_N_c_79_n N_A_N_c_80_n N_A_N_M1003_g
+ N_A_N_M1013_g A_N A_N A_N N_A_N_c_78_n PM_SKY130_FD_SC_HDLL__AND4B_4%A_N
x_PM_SKY130_FD_SC_HDLL__AND4B_4%A_184_21# N_A_184_21#_M1000_d
+ N_A_184_21#_M1016_d N_A_184_21#_M1004_d N_A_184_21#_c_116_n
+ N_A_184_21#_M1006_g N_A_184_21#_c_124_n N_A_184_21#_M1008_g
+ N_A_184_21#_c_117_n N_A_184_21#_M1007_g N_A_184_21#_c_125_n
+ N_A_184_21#_M1010_g N_A_184_21#_c_118_n N_A_184_21#_M1014_g
+ N_A_184_21#_c_126_n N_A_184_21#_M1011_g N_A_184_21#_c_119_n
+ N_A_184_21#_M1015_g N_A_184_21#_c_127_n N_A_184_21#_M1017_g
+ N_A_184_21#_c_120_n N_A_184_21#_c_129_n N_A_184_21#_c_142_p
+ N_A_184_21#_c_170_p N_A_184_21#_c_121_n N_A_184_21#_c_151_p
+ N_A_184_21#_c_122_n N_A_184_21#_c_123_n
+ PM_SKY130_FD_SC_HDLL__AND4B_4%A_184_21#
x_PM_SKY130_FD_SC_HDLL__AND4B_4%D N_D_c_239_n N_D_M1016_g N_D_c_240_n
+ N_D_M1002_g D D PM_SKY130_FD_SC_HDLL__AND4B_4%D
x_PM_SKY130_FD_SC_HDLL__AND4B_4%C N_C_c_267_n N_C_M1009_g N_C_c_268_n
+ N_C_M1001_g C C PM_SKY130_FD_SC_HDLL__AND4B_4%C
x_PM_SKY130_FD_SC_HDLL__AND4B_4%B N_B_c_296_n N_B_M1005_g N_B_c_297_n
+ N_B_M1004_g B B PM_SKY130_FD_SC_HDLL__AND4B_4%B
x_PM_SKY130_FD_SC_HDLL__AND4B_4%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1003_s
+ N_A_27_47#_c_331_n N_A_27_47#_M1000_g N_A_27_47#_c_336_n N_A_27_47#_M1012_g
+ N_A_27_47#_c_332_n N_A_27_47#_c_338_n N_A_27_47#_c_339_n N_A_27_47#_c_333_n
+ N_A_27_47#_c_334_n N_A_27_47#_c_341_n N_A_27_47#_c_335_n
+ PM_SKY130_FD_SC_HDLL__AND4B_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND4B_4%VPWR N_VPWR_M1003_d N_VPWR_M1010_d
+ N_VPWR_M1017_d N_VPWR_M1009_d N_VPWR_M1012_d N_VPWR_c_414_n N_VPWR_c_415_n
+ N_VPWR_c_416_n VPWR N_VPWR_c_417_n N_VPWR_c_418_n N_VPWR_c_419_n
+ N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_413_n
+ PM_SKY130_FD_SC_HDLL__AND4B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__AND4B_4%X N_X_M1006_s N_X_M1014_s N_X_M1008_s
+ N_X_M1011_s N_X_c_490_n N_X_c_498_n N_X_c_502_n N_X_c_507_n X X X N_X_c_493_n
+ X X PM_SKY130_FD_SC_HDLL__AND4B_4%X
x_PM_SKY130_FD_SC_HDLL__AND4B_4%VGND N_VGND_M1013_d N_VGND_M1007_d
+ N_VGND_M1015_d N_VGND_c_537_n N_VGND_c_538_n N_VGND_c_539_n N_VGND_c_540_n
+ N_VGND_c_541_n VGND N_VGND_c_542_n N_VGND_c_543_n N_VGND_c_544_n
+ N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n
+ PM_SKY130_FD_SC_HDLL__AND4B_4%VGND
cc_1 VNB N_A_N_M1013_g 0.0334873f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A_N 0.00546996f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.765
cc_3 VNB N_A_N_c_78_n 0.0270822f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.16
cc_4 VNB N_A_184_21#_c_116_n 0.0167071f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.765
cc_5 VNB N_A_184_21#_c_117_n 0.0166965f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.16
cc_6 VNB N_A_184_21#_c_118_n 0.0167366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_184_21#_c_119_n 0.0184873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_184_21#_c_120_n 0.00536809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_184_21#_c_121_n 0.0025288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_184_21#_c_122_n 0.00772384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_184_21#_c_123_n 0.0742298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_D_c_239_n 0.0273737f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_13 VNB N_D_c_240_n 0.0186714f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_14 VNB D 0.00203113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_C_c_267_n 0.0265992f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_16 VNB N_C_c_268_n 0.0161967f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_17 VNB C 0.00187039f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_18 VNB N_B_c_296_n 0.0166902f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_19 VNB N_B_c_297_n 0.0256606f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_20 VNB B 0.00326204f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_21 VNB N_A_27_47#_c_331_n 0.0225264f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_22 VNB N_A_27_47#_c_332_n 0.0334241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_333_n 0.00162417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_334_n 0.0128993f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.53
cc_25 VNB N_A_27_47#_c_335_n 0.0454575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_413_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB X 0.00106859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_537_n 0.00237268f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.445
cc_29 VNB N_VGND_c_538_n 4.17955e-19 $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.16
cc_30 VNB N_VGND_c_539_n 0.00507395f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.325
cc_31 VNB N_VGND_c_540_n 0.0168771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_541_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.16
cc_33 VNB N_VGND_c_542_n 0.0166487f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.53
cc_34 VNB N_VGND_c_543_n 0.017234f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_544_n 0.067158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_545_n 0.259805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_546_n 0.0035381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_547_n 0.00502664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VPB N_A_N_c_79_n 0.0348074f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_40 VPB N_A_N_c_80_n 0.0263351f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_41 VPB A_N 0.00195298f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=0.765
cc_42 VPB N_A_N_c_78_n 0.0048049f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.16
cc_43 VPB N_A_184_21#_c_124_n 0.016467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_184_21#_c_125_n 0.0157874f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_45 VPB N_A_184_21#_c_126_n 0.0160856f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.19
cc_46 VPB N_A_184_21#_c_127_n 0.0167386f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_184_21#_c_120_n 3.4877e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_184_21#_c_129_n 0.00301444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_184_21#_c_121_n 0.00174356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_184_21#_c_123_n 0.0468861f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_D_c_239_n 0.0275854f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_52 VPB N_C_c_267_n 0.0270315f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_53 VPB C 0.00110938f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_54 VPB N_B_c_297_n 0.0278996f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_55 VPB B 0.00194477f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_56 VPB N_A_27_47#_c_336_n 0.0182304f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=0.765
cc_57 VPB N_A_27_47#_c_332_n 0.029221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_338_n 0.0147617f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.16
cc_59 VPB N_A_27_47#_c_339_n 0.00224522f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_60 VPB N_A_27_47#_c_333_n 0.00644926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_47#_c_341_n 0.0110158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_47#_c_335_n 0.0173824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_414_n 0.0132269f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.16
cc_64 VPB N_VPWR_c_415_n 0.0087077f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_65 VPB N_VPWR_c_416_n 0.0175651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_417_n 0.0143107f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.53
cc_67 VPB N_VPWR_c_418_n 0.0157854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_419_n 0.0175377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_420_n 0.00810608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_421_n 0.00538861f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_422_n 0.00862719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_423_n 0.0249726f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_413_n 0.0440984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB X 0.00155996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 N_A_N_M1013_g N_A_184_21#_c_116_n 0.0193948f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_76 A_N N_A_184_21#_c_116_n 0.00520387f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_77 N_A_N_c_79_n N_A_184_21#_c_124_n 0.0208412f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_78 N_A_N_c_80_n N_A_184_21#_c_124_n 0.015366f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_79 A_N N_A_184_21#_c_124_n 0.00185147f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_80 N_A_N_c_79_n N_A_184_21#_c_123_n 0.00281774f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_81 N_A_N_c_78_n N_A_184_21#_c_123_n 0.0216201f $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_N_c_79_n N_A_27_47#_c_332_n 0.0168522f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_83 N_A_N_M1013_g N_A_27_47#_c_332_n 0.00716967f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_84 A_N N_A_27_47#_c_332_n 0.0646399f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_85 N_A_N_c_78_n N_A_27_47#_c_332_n 0.00775443f $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_N_c_80_n N_A_27_47#_c_338_n 0.00467732f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_87 N_A_N_c_80_n N_A_27_47#_c_339_n 0.0172144f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_88 A_N N_A_27_47#_c_339_n 0.021838f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_89 N_A_N_c_78_n N_A_27_47#_c_339_n 5.33633e-19 $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_90 A_N N_VPWR_M1003_d 0.00412295f $X=0.66 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_91 N_A_N_c_80_n N_VPWR_c_417_n 0.00315013f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_92 N_A_N_c_80_n N_VPWR_c_420_n 0.0109875f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_93 N_A_N_c_80_n N_VPWR_c_413_n 0.0046225f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_94 N_A_N_M1013_g N_X_c_490_n 4.43136e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_N_M1013_g X 6.02166e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_96 A_N X 0.0042163f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_97 N_A_N_c_79_n N_X_c_493_n 4.77684e-19 $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_98 A_N N_X_c_493_n 0.00689942f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_99 A_N X 0.0532601f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A_N_c_78_n X 2.75633e-19 $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_101 A_N N_VGND_M1013_d 0.00351948f $X=0.66 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_102 N_A_N_M1013_g N_VGND_c_537_n 0.0094371f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_103 A_N N_VGND_c_537_n 0.0150919f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_104 N_A_N_c_78_n N_VGND_c_537_n 4.16036e-19 $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_N_M1013_g N_VGND_c_542_n 0.0046653f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_N_M1013_g N_VGND_c_545_n 0.00519791f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_107 A_N N_VGND_c_545_n 0.00643138f $X=0.66 $Y=0.765 $X2=0 $Y2=0
cc_108 N_A_184_21#_c_127_n N_D_c_239_n 0.0292626f $X=2.43 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_184_21#_c_120_n N_D_c_239_n 0.00272373f $X=2.53 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_110 N_A_184_21#_c_129_n N_D_c_239_n 0.00451629f $X=2.615 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_184_21#_c_142_p N_D_c_239_n 0.0141956f $X=4.36 $Y=1.63 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_184_21#_c_123_n N_D_c_239_n 0.0153196f $X=2.405 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_113 N_A_184_21#_c_119_n N_D_c_240_n 0.0216649f $X=2.405 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_184_21#_c_120_n D 0.0272791f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_184_21#_c_142_p D 0.0126596f $X=4.36 $Y=1.63 $X2=0 $Y2=0
cc_116 N_A_184_21#_c_123_n D 2.72861e-19 $X=2.405 $Y=1.202 $X2=0 $Y2=0
cc_117 N_A_184_21#_c_142_p N_C_c_267_n 0.0115213f $X=4.36 $Y=1.63 $X2=-0.19
+ $Y2=-0.24
cc_118 N_A_184_21#_c_142_p C 0.0156423f $X=4.36 $Y=1.63 $X2=0 $Y2=0
cc_119 N_A_184_21#_c_121_n N_B_c_296_n 4.7301e-19 $X=4.445 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A_184_21#_c_151_p N_B_c_296_n 0.00245876f $X=4.53 $Y=0.725 $X2=-0.19
+ $Y2=-0.24
cc_121 N_A_184_21#_c_142_p N_B_c_297_n 0.0128028f $X=4.36 $Y=1.63 $X2=0 $Y2=0
cc_122 N_A_184_21#_c_121_n N_B_c_297_n 0.00599214f $X=4.445 $Y=1.545 $X2=0 $Y2=0
cc_123 N_A_184_21#_c_142_p B 0.0206496f $X=4.36 $Y=1.63 $X2=0 $Y2=0
cc_124 N_A_184_21#_c_121_n B 0.0396479f $X=4.445 $Y=1.545 $X2=0 $Y2=0
cc_125 N_A_184_21#_c_151_p B 0.00633981f $X=4.53 $Y=0.725 $X2=0 $Y2=0
cc_126 N_A_184_21#_c_121_n N_A_27_47#_c_331_n 0.00965007f $X=4.445 $Y=1.545
+ $X2=0 $Y2=0
cc_127 N_A_184_21#_c_151_p N_A_27_47#_c_331_n 0.00446778f $X=4.53 $Y=0.725 $X2=0
+ $Y2=0
cc_128 N_A_184_21#_c_122_n N_A_27_47#_c_331_n 0.0056493f $X=4.735 $Y=0.725 $X2=0
+ $Y2=0
cc_129 N_A_184_21#_c_142_p N_A_27_47#_c_336_n 0.00361166f $X=4.36 $Y=1.63 $X2=0
+ $Y2=0
cc_130 N_A_184_21#_c_121_n N_A_27_47#_c_336_n 0.00254145f $X=4.445 $Y=1.545
+ $X2=0 $Y2=0
cc_131 N_A_184_21#_M1016_d N_A_27_47#_c_339_n 0.00506751f $X=3.11 $Y=1.485 $X2=0
+ $Y2=0
cc_132 N_A_184_21#_M1004_d N_A_27_47#_c_339_n 0.00672307f $X=4.11 $Y=1.485 $X2=0
+ $Y2=0
cc_133 N_A_184_21#_c_124_n N_A_27_47#_c_339_n 0.0169293f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_134 N_A_184_21#_c_125_n N_A_27_47#_c_339_n 0.0131122f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_135 N_A_184_21#_c_126_n N_A_27_47#_c_339_n 0.0135818f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_136 N_A_184_21#_c_127_n N_A_27_47#_c_339_n 0.0155916f $X=2.43 $Y=1.41 $X2=0
+ $Y2=0
cc_137 N_A_184_21#_c_120_n N_A_27_47#_c_339_n 0.0042851f $X=2.53 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_184_21#_c_142_p N_A_27_47#_c_339_n 0.0897443f $X=4.36 $Y=1.63 $X2=0
+ $Y2=0
cc_139 N_A_184_21#_c_170_p N_A_27_47#_c_339_n 0.00886703f $X=2.7 $Y=1.63 $X2=0
+ $Y2=0
cc_140 N_A_184_21#_c_123_n N_A_27_47#_c_339_n 6.73635e-19 $X=2.405 $Y=1.202
+ $X2=0 $Y2=0
cc_141 N_A_184_21#_c_142_p N_A_27_47#_c_333_n 0.0125099f $X=4.36 $Y=1.63 $X2=0
+ $Y2=0
cc_142 N_A_184_21#_c_121_n N_A_27_47#_c_333_n 0.0355232f $X=4.445 $Y=1.545 $X2=0
+ $Y2=0
cc_143 N_A_184_21#_c_122_n N_A_27_47#_c_333_n 0.0123955f $X=4.735 $Y=0.725 $X2=0
+ $Y2=0
cc_144 N_A_184_21#_c_121_n N_A_27_47#_c_335_n 0.0106671f $X=4.445 $Y=1.545 $X2=0
+ $Y2=0
cc_145 N_A_184_21#_c_122_n N_A_27_47#_c_335_n 0.00523519f $X=4.735 $Y=0.725
+ $X2=0 $Y2=0
cc_146 N_A_184_21#_c_129_n N_VPWR_M1017_d 9.8524e-19 $X=2.615 $Y=1.545 $X2=0
+ $Y2=0
cc_147 N_A_184_21#_c_142_p N_VPWR_M1017_d 0.00703959f $X=4.36 $Y=1.63 $X2=0
+ $Y2=0
cc_148 N_A_184_21#_c_170_p N_VPWR_M1017_d 0.00261169f $X=2.7 $Y=1.63 $X2=0 $Y2=0
cc_149 N_A_184_21#_c_142_p N_VPWR_M1009_d 0.00970882f $X=4.36 $Y=1.63 $X2=0
+ $Y2=0
cc_150 N_A_184_21#_c_126_n N_VPWR_c_414_n 0.00453434f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_A_184_21#_c_127_n N_VPWR_c_414_n 0.00311736f $X=2.43 $Y=1.41 $X2=0
+ $Y2=0
cc_152 N_A_184_21#_c_124_n N_VPWR_c_418_n 0.00510113f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_153 N_A_184_21#_c_125_n N_VPWR_c_418_n 0.00311736f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_154 N_A_184_21#_c_124_n N_VPWR_c_420_n 0.00294646f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_155 N_A_184_21#_c_124_n N_VPWR_c_421_n 0.00122179f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_156 N_A_184_21#_c_125_n N_VPWR_c_421_n 0.0113834f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_184_21#_c_126_n N_VPWR_c_421_n 0.00820729f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_158 N_A_184_21#_c_127_n N_VPWR_c_421_n 0.00106505f $X=2.43 $Y=1.41 $X2=0
+ $Y2=0
cc_159 N_A_184_21#_c_126_n N_VPWR_c_422_n 0.00118604f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_160 N_A_184_21#_c_127_n N_VPWR_c_422_n 0.0112002f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_184_21#_M1016_d N_VPWR_c_413_n 0.00338665f $X=3.11 $Y=1.485 $X2=0
+ $Y2=0
cc_162 N_A_184_21#_M1004_d N_VPWR_c_413_n 0.00408734f $X=4.11 $Y=1.485 $X2=0
+ $Y2=0
cc_163 N_A_184_21#_c_124_n N_VPWR_c_413_n 0.00683693f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_184_21#_c_125_n N_VPWR_c_413_n 0.00375605f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_A_184_21#_c_126_n N_VPWR_c_413_n 0.00518254f $X=1.96 $Y=1.41 $X2=0
+ $Y2=0
cc_166 N_A_184_21#_c_127_n N_VPWR_c_413_n 0.00375605f $X=2.43 $Y=1.41 $X2=0
+ $Y2=0
cc_167 N_A_184_21#_c_116_n N_X_c_490_n 0.00631952f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_184_21#_c_117_n N_X_c_498_n 0.0163676f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_184_21#_c_118_n N_X_c_498_n 0.0117148f $X=1.935 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_184_21#_c_120_n N_X_c_498_n 0.048601f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_184_21#_c_123_n N_X_c_498_n 0.0063496f $X=2.405 $Y=1.202 $X2=0 $Y2=0
cc_172 N_A_184_21#_c_125_n N_X_c_502_n 0.0140558f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_184_21#_c_126_n N_X_c_502_n 0.0103731f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_184_21#_c_127_n N_X_c_502_n 0.0023821f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_184_21#_c_120_n N_X_c_502_n 0.042746f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_184_21#_c_123_n N_X_c_502_n 0.012208f $X=2.405 $Y=1.202 $X2=0 $Y2=0
cc_177 N_A_184_21#_c_118_n N_X_c_507_n 0.00418768f $X=1.935 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_184_21#_c_116_n X 0.00540833f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_184_21#_c_124_n N_X_c_493_n 0.0046246f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_184_21#_c_116_n X 0.00396032f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_184_21#_c_124_n X 0.0027388f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_184_21#_c_117_n X 0.0034321f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_184_21#_c_125_n X 0.00206809f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_184_21#_c_120_n X 0.0261825f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_184_21#_c_123_n X 0.0307164f $X=2.405 $Y=1.202 $X2=0 $Y2=0
cc_186 N_A_184_21#_c_116_n N_VGND_c_537_n 0.00392299f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_184_21#_c_116_n N_VGND_c_538_n 0.00103743f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_184_21#_c_117_n N_VGND_c_538_n 0.00817542f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_184_21#_c_118_n N_VGND_c_538_n 0.00751263f $X=1.935 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A_184_21#_c_119_n N_VGND_c_538_n 5.45278e-19 $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_184_21#_c_119_n N_VGND_c_539_n 0.00321134f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_184_21#_c_120_n N_VGND_c_539_n 0.00635328f $X=2.53 $Y=1.16 $X2=0
+ $Y2=0
cc_193 N_A_184_21#_c_118_n N_VGND_c_540_n 0.00341112f $X=1.935 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_184_21#_c_119_n N_VGND_c_540_n 0.00585385f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_184_21#_c_116_n N_VGND_c_543_n 0.00526178f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_184_21#_c_117_n N_VGND_c_543_n 0.00341112f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_184_21#_c_151_p N_VGND_c_544_n 0.0026036f $X=4.53 $Y=0.725 $X2=0
+ $Y2=0
cc_198 N_A_184_21#_c_122_n N_VGND_c_544_n 0.00590729f $X=4.735 $Y=0.725 $X2=0
+ $Y2=0
cc_199 N_A_184_21#_M1000_d N_VGND_c_545_n 0.00306852f $X=4.6 $Y=0.235 $X2=0
+ $Y2=0
cc_200 N_A_184_21#_c_116_n N_VGND_c_545_n 0.00953809f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_184_21#_c_117_n N_VGND_c_545_n 0.00410013f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_184_21#_c_118_n N_VGND_c_545_n 0.00410013f $X=1.935 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_184_21#_c_119_n N_VGND_c_545_n 0.0112463f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_184_21#_c_151_p N_VGND_c_545_n 0.00468565f $X=4.53 $Y=0.725 $X2=0
+ $Y2=0
cc_205 N_A_184_21#_c_122_n N_VGND_c_545_n 0.0100774f $X=4.735 $Y=0.725 $X2=0
+ $Y2=0
cc_206 N_A_184_21#_c_121_n A_814_47# 6.48296e-19 $X=4.445 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_207 N_A_184_21#_c_151_p A_814_47# 0.00265374f $X=4.53 $Y=0.725 $X2=-0.19
+ $Y2=-0.24
cc_208 N_D_c_239_n N_C_c_267_n 0.0652141f $X=3.02 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_209 D N_C_c_267_n 0.00113897f $X=2.995 $Y=1.19 $X2=-0.19 $Y2=-0.24
cc_210 N_D_c_240_n N_C_c_268_n 0.0362902f $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_211 N_D_c_239_n C 4.1478e-19 $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_212 N_D_c_240_n C 0.00540919f $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_213 D C 0.0203441f $X=2.995 $Y=1.19 $X2=0 $Y2=0
cc_214 N_D_c_239_n N_A_27_47#_c_339_n 0.0142936f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_215 N_D_c_239_n N_VPWR_c_415_n 0.00221617f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_216 N_D_c_239_n N_VPWR_c_416_n 0.00510113f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_217 N_D_c_239_n N_VPWR_c_422_n 0.00923358f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_218 N_D_c_239_n N_VPWR_c_413_n 0.00716145f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_219 N_D_c_239_n N_VGND_c_539_n 0.00184285f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_220 N_D_c_240_n N_VGND_c_539_n 0.00862748f $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_221 N_D_c_240_n N_VGND_c_544_n 0.00585385f $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_222 N_D_c_240_n N_VGND_c_545_n 0.0114566f $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_223 N_C_c_268_n N_B_c_296_n 0.0366786f $X=3.515 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_224 C N_B_c_296_n 4.03026e-19 $X=3.405 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_225 N_C_c_267_n N_B_c_297_n 0.0571094f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_226 C N_B_c_297_n 3.40276e-19 $X=3.405 $Y=0.765 $X2=0 $Y2=0
cc_227 N_C_c_267_n B 0.00218188f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_228 N_C_c_268_n B 0.00126232f $X=3.515 $Y=0.995 $X2=0 $Y2=0
cc_229 C B 0.04079f $X=3.405 $Y=0.765 $X2=0 $Y2=0
cc_230 N_C_c_267_n N_A_27_47#_c_339_n 0.0133477f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_231 N_C_c_267_n N_VPWR_c_415_n 0.0123252f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_232 N_C_c_267_n N_VPWR_c_416_n 0.00311736f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_233 N_C_c_267_n N_VPWR_c_413_n 0.00378223f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_234 N_C_c_268_n N_VGND_c_544_n 0.00441743f $X=3.515 $Y=0.995 $X2=0 $Y2=0
cc_235 C N_VGND_c_544_n 0.00359489f $X=3.405 $Y=0.765 $X2=0 $Y2=0
cc_236 N_C_c_268_n N_VGND_c_545_n 0.00649598f $X=3.515 $Y=0.995 $X2=0 $Y2=0
cc_237 C N_VGND_c_545_n 0.00763934f $X=3.405 $Y=0.765 $X2=0 $Y2=0
cc_238 C A_624_47# 0.00274039f $X=3.405 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_239 N_B_c_296_n N_A_27_47#_c_331_n 0.0305402f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_240 B N_A_27_47#_c_331_n 8.15039e-19 $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_241 N_B_c_297_n N_A_27_47#_c_336_n 0.0313704f $X=4.02 $Y=1.41 $X2=0 $Y2=0
cc_242 N_B_c_297_n N_A_27_47#_c_339_n 0.0143402f $X=4.02 $Y=1.41 $X2=0 $Y2=0
cc_243 N_B_c_297_n N_A_27_47#_c_335_n 0.0233493f $X=4.02 $Y=1.41 $X2=0 $Y2=0
cc_244 B N_A_27_47#_c_335_n 3.15965e-19 $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_245 N_B_c_297_n N_VPWR_c_415_n 0.00436918f $X=4.02 $Y=1.41 $X2=0 $Y2=0
cc_246 N_B_c_297_n N_VPWR_c_419_n 0.00510113f $X=4.02 $Y=1.41 $X2=0 $Y2=0
cc_247 N_B_c_297_n N_VPWR_c_423_n 0.00210708f $X=4.02 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B_c_297_n N_VPWR_c_413_n 0.00702798f $X=4.02 $Y=1.41 $X2=0 $Y2=0
cc_249 N_B_c_296_n N_VGND_c_544_n 0.00439071f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_250 B N_VGND_c_544_n 0.00478585f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_251 N_B_c_296_n N_VGND_c_545_n 0.00657939f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_252 B N_VGND_c_545_n 0.00972142f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_253 B A_718_47# 0.00245366f $X=3.825 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_254 B A_814_47# 0.00258501f $X=3.825 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_255 N_A_27_47#_c_339_n N_VPWR_M1003_d 0.00586137f $X=4.715 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_256 N_A_27_47#_c_339_n N_VPWR_M1010_d 0.00362631f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_339_n N_VPWR_M1017_d 0.00705129f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_339_n N_VPWR_M1009_d 0.005075f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_339_n N_VPWR_M1012_d 0.0105254f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_333_n N_VPWR_M1012_d 0.0232645f $X=4.8 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_339_n N_VPWR_c_414_n 0.00861424f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_339_n N_VPWR_c_415_n 0.0228926f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_339_n N_VPWR_c_416_n 0.0102519f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_338_n N_VPWR_c_417_n 0.0181194f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_339_n N_VPWR_c_417_n 0.00238709f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_339_n N_VPWR_c_418_n 0.00928399f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_336_n N_VPWR_c_419_n 0.00311027f $X=4.55 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_339_n N_VPWR_c_419_n 0.0103733f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_338_n N_VPWR_c_420_n 0.0161786f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_339_n N_VPWR_c_420_n 0.0225111f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_339_n N_VPWR_c_421_n 0.0196308f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_339_n N_VPWR_c_422_n 0.0241133f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_336_n N_VPWR_c_423_n 0.0136446f $X=4.55 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_339_n N_VPWR_c_423_n 0.0205438f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_275 N_A_27_47#_M1003_s N_VPWR_c_413_n 0.00238238f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_336_n N_VPWR_c_413_n 0.00390769f $X=4.55 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_338_n N_VPWR_c_413_n 0.00991829f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_339_n N_VPWR_c_413_n 0.0786087f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_339_n N_X_M1008_s 0.00489221f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_339_n N_X_M1011_s 0.004896f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_339_n N_X_c_502_n 0.0451915f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_339_n N_X_c_493_n 0.0179584f $X=4.715 $Y=2 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_334_n N_VGND_c_537_n 0.0177603f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_334_n N_VGND_c_542_n 0.0179125f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_331_n N_VGND_c_544_n 0.00425753f $X=4.525 $Y=0.995 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1013_s N_VGND_c_545_n 0.00584642f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_331_n N_VGND_c_545_n 0.00722198f $X=4.525 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_334_n N_VGND_c_545_n 0.00987844f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_289 N_VPWR_c_413_n N_X_M1008_s 0.00338665f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_290 N_VPWR_c_413_n N_X_M1011_s 0.00338665f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_291 N_VPWR_M1010_d N_X_c_502_n 0.00366978f $X=1.58 $Y=1.485 $X2=0 $Y2=0
cc_292 N_X_c_498_n N_VGND_M1007_d 0.00405996f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_293 N_X_c_490_n N_VGND_c_537_n 0.0183101f $X=1.255 $Y=0.42 $X2=0 $Y2=0
cc_294 N_X_c_498_n N_VGND_c_538_n 0.0188758f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_295 N_X_c_507_n N_VGND_c_538_n 0.01316f $X=2.195 $Y=0.42 $X2=0 $Y2=0
cc_296 N_X_c_498_n N_VGND_c_540_n 0.00314446f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_297 N_X_c_507_n N_VGND_c_540_n 0.0114519f $X=2.195 $Y=0.42 $X2=0 $Y2=0
cc_298 N_X_c_490_n N_VGND_c_543_n 0.0193477f $X=1.255 $Y=0.42 $X2=0 $Y2=0
cc_299 N_X_c_498_n N_VGND_c_543_n 0.00216966f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_300 N_X_M1006_s N_VGND_c_545_n 0.00273459f $X=1.07 $Y=0.235 $X2=0 $Y2=0
cc_301 N_X_M1014_s N_VGND_c_545_n 0.00466393f $X=2.01 $Y=0.235 $X2=0 $Y2=0
cc_302 N_X_c_490_n N_VGND_c_545_n 0.0116108f $X=1.255 $Y=0.42 $X2=0 $Y2=0
cc_303 N_X_c_498_n N_VGND_c_545_n 0.0107874f $X=2.11 $Y=0.735 $X2=0 $Y2=0
cc_304 N_X_c_507_n N_VGND_c_545_n 0.0064389f $X=2.195 $Y=0.42 $X2=0 $Y2=0
cc_305 X N_VGND_c_545_n 5.95167e-19 $X=1.17 $Y=0.765 $X2=0 $Y2=0
cc_306 N_VGND_c_545_n A_624_47# 0.0104837f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
cc_307 N_VGND_c_545_n A_718_47# 0.00944229f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
cc_308 N_VGND_c_545_n A_814_47# 0.00992884f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
