* File: sky130_fd_sc_hdll__nand3b_1.spice
* Created: Thu Aug 27 19:13:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand3b_1.pex.spice"
.subckt sky130_fd_sc_hdll__nand3b_1  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_N_M1003_g N_A_53_93#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0914579 AS=0.1302 PD=0.812523 PS=1.46 NRD=46.5 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1006 A_252_47# N_C_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.141542 PD=0.98 PS=1.25748 NRD=20.304 NRS=8.304 M=1 R=4.33333 SA=75000.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1002 A_348_47# N_B_M1002_g A_252_47# VNB NSHORT L=0.15 W=0.65 AD=0.105625
+ AS=0.10725 PD=0.975 PS=0.98 NRD=19.836 NRS=20.304 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_A_53_93#_M1004_g A_348_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.105625 PD=1.87 PS=0.975 NRD=0 NRS=19.836 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_53_93#_M1000_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0904183 AS=0.1134 PD=0.801549 PS=1.38 NRD=32.8202 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1005 N_Y_M1005_d N_C_M1005_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.215282 PD=1.3 PS=1.90845 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.4
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_Y_M1005_d VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=0.9653 NRS=2.9353 M=1 R=5.55556 SA=90000.9
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1007 N_Y_M1007_d N_A_53_93#_M1007_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.15 PD=2.58 PS=1.3 NRD=0.9653 NRS=2.9353 M=1 R=5.55556 SA=90001.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
pX9_noxref noxref_12 B B PROBETYPE=1
c_43 VPB 0 1.78374e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__nand3b_1.pxi.spice"
*
.ends
*
*
