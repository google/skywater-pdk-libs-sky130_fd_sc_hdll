* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
X0 a_514_297# C a_305_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_754_21# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 Y a_754_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_305_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_297# B a_305_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y a_754_21# a_514_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_754_21# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_514_297# a_754_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VGND a_754_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_305_297# C a_514_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
