* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or4_1 A B C D VGND VNB VPB VPWR X
M1000 a_27_297# D VGND VNB nshort w=420000u l=150000u
+  ad=3.15e+11p pd=3.18e+06u as=4.7985e+11p ps=4.92e+06u
M1001 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.73e+11p pd=2.14e+06u as=0p ps=0u
M1002 VGND A a_27_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_117_297# D a_27_297# VPB phighvt w=420000u l=180000u
+  ad=1.47e+11p pd=1.54e+06u as=1.134e+11p ps=1.38e+06u
M1004 VPWR A a_307_297# VPB phighvt w=420000u l=180000u
+  ad=3.107e+11p pd=2.72e+06u as=1.428e+11p ps=1.52e+06u
M1005 VGND C a_27_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_307_297# B a_223_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_27_297# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.3e+11p pd=2.86e+06u as=0p ps=0u
M1009 a_223_297# C a_117_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
