* File: sky130_fd_sc_hdll__clkinv_1.spice
* Created: Wed Sep  2 08:26:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkinv_1.pex.spice"
.subckt sky130_fd_sc_hdll__clkinv_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.1323 PD=1.41 PS=1.47 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.2 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=0.84
+ AD=0.1218 AS=0.2268 PD=1.13 PS=2.22 NRD=1.1623 NRS=1.1623 M=1 R=4.66667
+ SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1002 N_Y_M1001_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=0.84
+ AD=0.1218 AS=0.2436 PD=1.13 PS=2.26 NRD=1.1623 NRS=1.1623 M=1 R=4.66667
+ SA=90000.6 SB=90000.2 A=0.1512 P=2.04 MULT=1
DX3_noxref VNB VPB NWDIODE A=3.5631 P=7.65
pX4_noxref noxref_7 Y Y PROBETYPE=1
pX5_noxref noxref_8 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__clkinv_1.pxi.spice"
*
.ends
*
*
