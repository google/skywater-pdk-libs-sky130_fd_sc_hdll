* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__einvp_1 A TE VGND VNB VPB VPWR Z
M1000 a_332_297# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=4.55e+11p pd=2.91e+06u as=8.457e+11p ps=3.79e+06u
M1001 VPWR TE a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1002 Z A a_204_47# VNB nshort w=650000u l=150000u
+  ad=2.08e+11p pd=1.94e+06u as=7.0525e+11p ps=3.47e+06u
M1003 VGND TE a_27_47# VNB nshort w=420000u l=150000u
+  ad=1.94e+11p pd=1.95e+06u as=1.092e+11p ps=1.36e+06u
M1004 Z A a_332_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1005 a_204_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
