* File: sky130_fd_sc_hdll__sdfrtp_4.pxi.spice
* Created: Wed Sep  2 08:51:20 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%CLK N_CLK_c_269_n N_CLK_M1016_g N_CLK_c_266_n
+ N_CLK_M1031_g CLK CLK N_CLK_c_268_n PM_SKY130_FD_SC_HDLL__SDFRTP_4%CLK
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_27_47# N_A_27_47#_M1031_s N_A_27_47#_M1016_s
+ N_A_27_47#_c_297_n N_A_27_47#_M1033_g N_A_27_47#_c_298_n N_A_27_47#_M1002_g
+ N_A_27_47#_c_299_n N_A_27_47#_c_300_n N_A_27_47#_c_301_n N_A_27_47#_c_302_n
+ N_A_27_47#_M1010_g N_A_27_47#_c_320_n N_A_27_47#_c_321_n N_A_27_47#_M1026_g
+ N_A_27_47#_c_322_n N_A_27_47#_c_323_n N_A_27_47#_M1035_g N_A_27_47#_M1027_g
+ N_A_27_47#_c_304_n N_A_27_47#_c_305_n N_A_27_47#_c_306_n N_A_27_47#_c_334_n
+ N_A_27_47#_c_307_n N_A_27_47#_c_339_n N_A_27_47#_c_325_n N_A_27_47#_c_326_n
+ N_A_27_47#_c_308_n N_A_27_47#_c_344_n N_A_27_47#_c_309_n N_A_27_47#_c_416_p
+ N_A_27_47#_c_310_n N_A_27_47#_c_311_n N_A_27_47#_c_312_n N_A_27_47#_c_313_n
+ N_A_27_47#_c_314_n N_A_27_47#_c_315_n N_A_27_47#_c_316_n N_A_27_47#_c_317_n
+ PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_331_66# N_A_331_66#_M1040_s
+ N_A_331_66#_M1030_s N_A_331_66#_c_565_n N_A_331_66#_c_566_n
+ N_A_331_66#_M1021_g N_A_331_66#_c_567_n N_A_331_66#_M1039_g
+ N_A_331_66#_c_648_p N_A_331_66#_c_568_n N_A_331_66#_c_569_n
+ N_A_331_66#_c_652_p N_A_331_66#_c_578_n N_A_331_66#_c_579_n
+ N_A_331_66#_c_570_n N_A_331_66#_c_571_n N_A_331_66#_c_572_n
+ N_A_331_66#_c_573_n N_A_331_66#_c_574_n N_A_331_66#_c_575_n
+ N_A_331_66#_c_576_n PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_331_66#
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%D N_D_c_709_n N_D_M1020_g N_D_M1008_g D D
+ PM_SKY130_FD_SC_HDLL__SDFRTP_4%D
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%SCE N_SCE_M1040_g N_SCE_c_759_n N_SCE_c_753_n
+ N_SCE_c_754_n N_SCE_c_760_n N_SCE_c_761_n N_SCE_c_762_n N_SCE_M1030_g
+ N_SCE_c_763_n N_SCE_c_764_n N_SCE_M1017_g N_SCE_c_755_n N_SCE_M1034_g
+ N_SCE_c_756_n N_SCE_c_757_n N_SCE_c_767_n SCE SCE
+ PM_SKY130_FD_SC_HDLL__SDFRTP_4%SCE
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%SCD N_SCD_c_857_n N_SCD_M1007_g N_SCD_M1038_g
+ SCD SCD PM_SKY130_FD_SC_HDLL__SDFRTP_4%SCD
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_213_47# N_A_213_47#_M1002_d
+ N_A_213_47#_M1033_d N_A_213_47#_c_904_n N_A_213_47#_M1025_g
+ N_A_213_47#_c_894_n N_A_213_47#_M1036_g N_A_213_47#_c_895_n
+ N_A_213_47#_M1028_g N_A_213_47#_c_905_n N_A_213_47#_M1018_g
+ N_A_213_47#_c_896_n N_A_213_47#_c_897_n N_A_213_47#_c_898_n
+ N_A_213_47#_c_899_n N_A_213_47#_c_907_n N_A_213_47#_c_1027_p
+ N_A_213_47#_c_900_n N_A_213_47#_c_908_n N_A_213_47#_c_901_n
+ N_A_213_47#_c_910_n N_A_213_47#_c_911_n N_A_213_47#_c_912_n
+ N_A_213_47#_c_913_n N_A_213_47#_c_914_n N_A_213_47#_c_915_n
+ N_A_213_47#_c_916_n N_A_213_47#_c_917_n N_A_213_47#_c_902_n
+ N_A_213_47#_c_918_n N_A_213_47#_c_903_n
+ PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_213_47#
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1380_303# N_A_1380_303#_M1041_d
+ N_A_1380_303#_M1009_d N_A_1380_303#_c_1149_n N_A_1380_303#_M1015_g
+ N_A_1380_303#_M1000_g N_A_1380_303#_c_1151_n N_A_1380_303#_c_1175_n
+ N_A_1380_303#_c_1160_n N_A_1380_303#_c_1163_n N_A_1380_303#_c_1196_p
+ N_A_1380_303#_c_1164_n N_A_1380_303#_c_1152_n N_A_1380_303#_c_1148_n
+ PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1380_303#
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%RESET_B N_RESET_B_M1022_g N_RESET_B_c_1255_n
+ N_RESET_B_c_1269_n N_RESET_B_M1023_g N_RESET_B_M1006_g N_RESET_B_c_1270_n
+ N_RESET_B_c_1271_n N_RESET_B_M1004_g N_RESET_B_c_1257_n N_RESET_B_c_1258_n
+ N_RESET_B_c_1259_n N_RESET_B_c_1260_n N_RESET_B_c_1261_n N_RESET_B_c_1262_n
+ RESET_B N_RESET_B_c_1264_n N_RESET_B_c_1265_n N_RESET_B_c_1266_n
+ N_RESET_B_c_1267_n PM_SKY130_FD_SC_HDLL__SDFRTP_4%RESET_B
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1202_413# N_A_1202_413#_M1010_d
+ N_A_1202_413#_M1025_d N_A_1202_413#_M1041_g N_A_1202_413#_c_1429_n
+ N_A_1202_413#_c_1430_n N_A_1202_413#_M1009_g N_A_1202_413#_c_1462_n
+ N_A_1202_413#_c_1423_n N_A_1202_413#_c_1424_n N_A_1202_413#_c_1425_n
+ N_A_1202_413#_c_1426_n N_A_1202_413#_c_1447_n N_A_1202_413#_c_1433_n
+ N_A_1202_413#_c_1434_n N_A_1202_413#_c_1427_n N_A_1202_413#_c_1428_n
+ PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1202_413#
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1972_21# N_A_1972_21#_M1012_d
+ N_A_1972_21#_M1004_d N_A_1972_21#_M1032_g N_A_1972_21#_c_1562_n
+ N_A_1972_21#_c_1580_n N_A_1972_21#_M1003_g N_A_1972_21#_c_1563_n
+ N_A_1972_21#_M1013_g N_A_1972_21#_c_1581_n N_A_1972_21#_M1001_g
+ N_A_1972_21#_c_1564_n N_A_1972_21#_c_1565_n N_A_1972_21#_c_1584_n
+ N_A_1972_21#_M1005_g N_A_1972_21#_c_1566_n N_A_1972_21#_M1014_g
+ N_A_1972_21#_c_1585_n N_A_1972_21#_M1024_g N_A_1972_21#_c_1567_n
+ N_A_1972_21#_M1019_g N_A_1972_21#_c_1586_n N_A_1972_21#_M1037_g
+ N_A_1972_21#_c_1568_n N_A_1972_21#_M1029_g N_A_1972_21#_c_1569_n
+ N_A_1972_21#_c_1570_n N_A_1972_21#_c_1571_n N_A_1972_21#_c_1572_n
+ N_A_1972_21#_c_1573_n N_A_1972_21#_c_1574_n N_A_1972_21#_c_1626_n
+ N_A_1972_21#_c_1669_p N_A_1972_21#_c_1588_n N_A_1972_21#_c_1589_n
+ N_A_1972_21#_c_1575_n N_A_1972_21#_c_1590_n N_A_1972_21#_c_1576_n
+ N_A_1972_21#_c_1577_n N_A_1972_21#_c_1578_n
+ PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1972_21#
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1757_47# N_A_1757_47#_M1028_d
+ N_A_1757_47#_M1035_d N_A_1757_47#_M1012_g N_A_1757_47#_c_1758_n
+ N_A_1757_47#_M1011_g N_A_1757_47#_c_1754_n N_A_1757_47#_c_1755_n
+ N_A_1757_47#_c_1756_n N_A_1757_47#_c_1764_n N_A_1757_47#_c_1767_n
+ N_A_1757_47#_c_1757_n N_A_1757_47#_c_1761_n N_A_1757_47#_c_1762_n
+ N_A_1757_47#_c_1763_n PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1757_47#
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%VPWR N_VPWR_M1016_d N_VPWR_M1030_d
+ N_VPWR_M1007_d N_VPWR_M1015_d N_VPWR_M1009_s N_VPWR_M1003_d N_VPWR_M1011_d
+ N_VPWR_M1001_s N_VPWR_M1005_s N_VPWR_M1037_s N_VPWR_c_1870_n N_VPWR_c_1871_n
+ N_VPWR_c_1872_n N_VPWR_c_1873_n N_VPWR_c_1874_n N_VPWR_c_1875_n
+ N_VPWR_c_1876_n N_VPWR_c_1877_n N_VPWR_c_1878_n N_VPWR_c_1879_n
+ N_VPWR_c_1880_n N_VPWR_c_1881_n N_VPWR_c_1882_n N_VPWR_c_1883_n
+ N_VPWR_c_1884_n N_VPWR_c_1885_n N_VPWR_c_1886_n N_VPWR_c_1887_n
+ N_VPWR_c_1888_n N_VPWR_c_1889_n VPWR N_VPWR_c_1890_n N_VPWR_c_1891_n
+ N_VPWR_c_1892_n N_VPWR_c_1893_n N_VPWR_c_1894_n N_VPWR_c_1895_n
+ N_VPWR_c_1896_n N_VPWR_c_1897_n N_VPWR_c_1869_n VPWR
+ PM_SKY130_FD_SC_HDLL__SDFRTP_4%VPWR
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_700_389# N_A_700_389#_M1008_d
+ N_A_700_389#_M1010_s N_A_700_389#_M1020_d N_A_700_389#_M1025_s
+ N_A_700_389#_c_2078_n N_A_700_389#_c_2110_n N_A_700_389#_c_2086_n
+ N_A_700_389#_c_2079_n N_A_700_389#_c_2080_n N_A_700_389#_c_2081_n
+ N_A_700_389#_c_2082_n N_A_700_389#_c_2083_n N_A_700_389#_c_2123_n
+ N_A_700_389#_c_2084_n PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_700_389#
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1324_413# N_A_1324_413#_M1026_d
+ N_A_1324_413#_M1023_d N_A_1324_413#_c_2177_n N_A_1324_413#_c_2178_n
+ N_A_1324_413#_c_2179_n PM_SKY130_FD_SC_HDLL__SDFRTP_4%A_1324_413#
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%Q N_Q_M1013_s N_Q_M1019_s N_Q_M1001_d
+ N_Q_M1024_d N_Q_c_2214_n N_Q_c_2210_n N_Q_c_2212_n N_Q_c_2220_n N_Q_c_2223_n Q
+ Q Q Q PM_SKY130_FD_SC_HDLL__SDFRTP_4%Q
x_PM_SKY130_FD_SC_HDLL__SDFRTP_4%VGND N_VGND_M1031_d N_VGND_M1040_d
+ N_VGND_M1021_s N_VGND_M1038_d N_VGND_M1022_d N_VGND_M1032_d N_VGND_M1013_d
+ N_VGND_M1014_d N_VGND_M1029_d N_VGND_c_2249_n N_VGND_c_2250_n N_VGND_c_2251_n
+ N_VGND_c_2252_n N_VGND_c_2253_n N_VGND_c_2254_n N_VGND_c_2255_n
+ N_VGND_c_2256_n N_VGND_c_2257_n N_VGND_c_2258_n N_VGND_c_2259_n
+ N_VGND_c_2260_n N_VGND_c_2261_n N_VGND_c_2262_n N_VGND_c_2263_n
+ N_VGND_c_2264_n N_VGND_c_2265_n VGND N_VGND_c_2266_n N_VGND_c_2267_n
+ N_VGND_c_2268_n N_VGND_c_2269_n N_VGND_c_2270_n N_VGND_c_2271_n
+ N_VGND_c_2272_n N_VGND_c_2273_n N_VGND_c_2274_n N_VGND_c_2275_n VGND
+ PM_SKY130_FD_SC_HDLL__SDFRTP_4%VGND
cc_1 VNB N_CLK_c_266_n 0.0217391f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB CLK 0.00359948f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.105
cc_3 VNB N_CLK_c_268_n 0.0473545f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_A_27_47#_c_297_n 0.026472f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_5 VNB N_A_27_47#_c_298_n 0.0198797f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_299_n 0.0188356f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_7 VNB N_A_27_47#_c_300_n 0.00966649f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_8 VNB N_A_27_47#_c_301_n 0.0242657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_302_n 0.0184982f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.53
cc_10 VNB N_A_27_47#_M1027_g 0.0320594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_304_n 0.00710356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_305_n 0.014131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_306_n 0.011157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_307_n 0.00785455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_308_n 0.0432266f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_309_n 0.0197565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_310_n 8.25118e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_311_n 0.00234825f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_312_n 0.0152776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_313_n 6.9625e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_314_n 0.00299094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_315_n 0.0194936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_316_n 0.013946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_317_n 0.00172224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_331_66#_c_565_n 0.0202226f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_26 VNB N_A_331_66#_c_566_n 0.0150055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_331_66#_c_567_n 0.0115482f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_28 VNB N_A_331_66#_c_568_n 0.00213996f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.53
cc_29 VNB N_A_331_66#_c_569_n 0.0028631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_331_66#_c_570_n 0.00283418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_331_66#_c_571_n 0.0182067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_331_66#_c_572_n 0.00399684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_331_66#_c_573_n 0.00854157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_331_66#_c_574_n 0.00288141f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_331_66#_c_575_n 0.00659246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_331_66#_c_576_n 0.0359217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_D_M1008_g 0.0363739f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_38 VNB D 0.00422214f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.105
cc_39 VNB N_SCE_M1040_g 0.0324301f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_40 VNB N_SCE_c_753_n 0.167758f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_41 VNB N_SCE_c_754_n 0.0124454f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.105
cc_42 VNB N_SCE_c_755_n 0.033266f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.53
cc_43 VNB N_SCE_c_756_n 0.0218643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_SCE_c_757_n 0.00524045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB SCE 0.00913086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_SCD_M1038_g 0.0524162f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_47 VNB SCD 0.00510088f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_48 VNB N_A_213_47#_c_894_n 0.0185188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_213_47#_c_895_n 0.0180202f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_50 VNB N_A_213_47#_c_896_n 0.00327111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_213_47#_c_897_n 0.00493253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_213_47#_c_898_n 0.00475961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_213_47#_c_899_n 0.0364536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_213_47#_c_900_n 0.00413034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_213_47#_c_901_n 0.0107257f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_213_47#_c_902_n 0.0329211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_213_47#_c_903_n 0.00571541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1380_303#_M1000_g 0.0464983f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_59 VNB N_A_1380_303#_c_1148_n 0.00640816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_RESET_B_c_1255_n 0.00874394f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_61 VNB N_RESET_B_M1006_g 0.029376f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.202
cc_62 VNB N_RESET_B_c_1257_n 0.0054841f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_RESET_B_c_1258_n 0.00731205f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_RESET_B_c_1259_n 0.00815027f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_RESET_B_c_1260_n 0.0231888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_RESET_B_c_1261_n 0.00125033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_RESET_B_c_1262_n 9.86606e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB RESET_B 0.00541831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_RESET_B_c_1264_n 0.0338798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_RESET_B_c_1265_n 0.0180031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_RESET_B_c_1266_n 0.0242951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_RESET_B_c_1267_n 0.00381782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1202_413#_M1041_g 0.0196344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1202_413#_c_1423_n 0.00309971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1202_413#_c_1424_n 7.14483e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1202_413#_c_1425_n 0.00676602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1202_413#_c_1426_n 0.00363358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1202_413#_c_1427_n 0.00186995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1202_413#_c_1428_n 0.0311233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1972_21#_M1032_g 0.023316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1972_21#_c_1562_n 0.011426f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_82 VNB N_A_1972_21#_c_1563_n 0.0214459f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_83 VNB N_A_1972_21#_c_1564_n 0.0207077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1972_21#_c_1565_n 0.0233217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1972_21#_c_1566_n 0.0183132f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1972_21#_c_1567_n 0.0170119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1972_21#_c_1568_n 0.0224185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1972_21#_c_1569_n 0.065872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1972_21#_c_1570_n 0.00124594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1972_21#_c_1571_n 0.00503624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1972_21#_c_1572_n 0.00283498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_1972_21#_c_1573_n 4.84338e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_1972_21#_c_1574_n 0.00321973f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_1972_21#_c_1575_n 0.0107857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_1972_21#_c_1576_n 0.00822564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_1972_21#_c_1577_n 0.00380069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_1972_21#_c_1578_n 0.0513529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_1757_47#_c_1754_n 0.0290875f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_99 VNB N_A_1757_47#_c_1755_n 0.0179786f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_100 VNB N_A_1757_47#_c_1756_n 0.0136715f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_101 VNB N_A_1757_47#_c_1757_n 0.00998098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VPWR_c_1869_n 0.592346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_A_700_389#_c_2078_n 0.0083542f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=1.202
cc_104 VNB N_A_700_389#_c_2079_n 0.00717059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_A_700_389#_c_2080_n 0.00522158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_A_700_389#_c_2081_n 0.00179289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_A_700_389#_c_2082_n 0.00335972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_A_700_389#_c_2083_n 0.00550481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_A_700_389#_c_2084_n 0.00207602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_Q_c_2210_n 0.00204933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB Q 0.00217709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2249_n 0.00313571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2250_n 0.00940761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2251_n 0.00789808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2252_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2253_n 0.00502493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2254_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2255_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2256_n 0.0110259f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2257_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2258_n 0.0624319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2259_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2260_n 0.0519427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2261_n 0.00420332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2262_n 0.0389443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2263_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2264_n 0.0255501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2265_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2266_n 0.0147814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2267_n 0.0314065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2268_n 0.00610401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2269_n 0.048703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2270_n 0.0221513f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2271_n 0.0085923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2272_n 0.00503248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2273_n 0.00506042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2274_n 0.00607822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2275_n 0.674213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VPB N_CLK_c_269_n 0.0194814f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_140 VPB CLK 0.00525533f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.105
cc_141 VPB N_CLK_c_268_n 0.0183416f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_142 VPB N_A_27_47#_c_297_n 0.0299778f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_143 VPB N_A_27_47#_c_301_n 0.0255566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_320_n 0.0298423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_321_n 0.0232068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_27_47#_c_322_n 0.0296308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_27_47#_c_323_n 0.0231363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_27_47#_c_304_n 0.0101789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_27_47#_c_325_n 0.00101836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_27_47#_c_326_n 0.0273613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_27_47#_c_310_n 0.00218623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_27_47#_c_315_n 0.0151139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_331_66#_c_567_n 0.0585648f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_154 VPB N_A_331_66#_c_578_n 0.00401635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_331_66#_c_579_n 0.00499376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_331_66#_c_576_n 0.00469895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_D_c_709_n 0.0542123f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_158 VPB N_D_M1008_g 0.00190701f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_159 VPB D 0.00874572f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.105
cc_160 VPB N_SCE_c_759_n 0.00900744f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_161 VPB N_SCE_c_760_n 0.0206729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_SCE_c_761_n 0.0125604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_SCE_c_762_n 0.0193341f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.202
cc_164 VPB N_SCE_c_763_n 0.0313194f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_165 VPB N_SCE_c_764_n 0.0150959f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_166 VPB N_SCE_c_756_n 0.0234869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_SCE_c_757_n 0.00608926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_SCE_c_767_n 0.0121283f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB SCE 0.00973562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_SCD_c_857_n 0.0636323f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_171 VPB N_SCD_M1038_g 0.00409327f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_172 VPB SCD 0.00331096f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_173 VPB N_A_213_47#_c_904_n 0.0630017f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_174 VPB N_A_213_47#_c_905_n 0.057532f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_175 VPB N_A_213_47#_c_898_n 0.00259103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_213_47#_c_907_n 0.00214341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_213_47#_c_908_n 0.00150413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_213_47#_c_901_n 0.00565136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_213_47#_c_910_n 0.00417155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_213_47#_c_911_n 0.0390412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_213_47#_c_912_n 0.00294907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_213_47#_c_913_n 0.012481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_213_47#_c_914_n 0.00250224f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_213_47#_c_915_n 0.0194717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_213_47#_c_916_n 0.0010731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_213_47#_c_917_n 0.00229693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_213_47#_c_918_n 0.00501095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_213_47#_c_903_n 0.00399787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1380_303#_c_1149_n 0.0630679f $X=-0.19 $Y=1.305 $X2=0.15
+ $Y2=1.445
cc_190 VPB N_A_1380_303#_M1000_g 0.0117713f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_191 VPB N_A_1380_303#_c_1151_n 0.0130444f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.202
cc_192 VPB N_A_1380_303#_c_1152_n 0.0043592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_1380_303#_c_1148_n 0.0017978f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_RESET_B_c_1255_n 0.0372278f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_195 VPB N_RESET_B_c_1269_n 0.0280009f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_196 VPB N_RESET_B_c_1270_n 0.0333369f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_197 VPB N_RESET_B_c_1271_n 0.0241989f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_198 VPB N_RESET_B_c_1262_n 0.00114586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_RESET_B_c_1266_n 0.0033882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1202_413#_c_1429_n 0.0291803f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.202
cc_201 VPB N_A_1202_413#_c_1430_n 0.0192179f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_202 VPB N_A_1202_413#_c_1423_n 0.00279025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_1202_413#_c_1426_n 0.00529458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_1202_413#_c_1433_n 0.00464467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_1202_413#_c_1434_n 0.00144164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_1202_413#_c_1427_n 0.00126247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_1202_413#_c_1428_n 0.024381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_1972_21#_c_1562_n 0.0342287f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_209 VPB N_A_1972_21#_c_1580_n 0.0235097f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_210 VPB N_A_1972_21#_c_1581_n 0.0191571f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.53
cc_211 VPB N_A_1972_21#_c_1564_n 0.0126144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_1972_21#_c_1565_n 0.0110606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_A_1972_21#_c_1584_n 0.0169401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_1972_21#_c_1585_n 0.0165614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_A_1972_21#_c_1586_n 0.0207627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_1972_21#_c_1569_n 0.0436994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_A_1972_21#_c_1588_n 0.0109459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_1972_21#_c_1589_n 0.00320057f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_A_1972_21#_c_1590_n 0.0136633f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_1972_21#_c_1576_n 0.0071168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1972_21#_c_1577_n 5.18967e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_A_1757_47#_c_1758_n 0.0602032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_1757_47#_c_1754_n 0.0125276f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.202
cc_224 VPB N_A_1757_47#_c_1757_n 2.26879e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_1757_47#_c_1761_n 0.00207751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_1757_47#_c_1762_n 0.0151024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1757_47#_c_1763_n 0.0209467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1870_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1871_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1872_n 0.00539287f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1873_n 0.0110604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1874_n 0.00234852f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1875_n 0.014528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1876_n 0.00124395f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1877_n 0.00242779f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1878_n 0.0100141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1879_n 0.043756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1880_n 0.0462152f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1881_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1882_n 0.0485087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1883_n 0.00539544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1884_n 0.0110643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1885_n 0.0506362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1886_n 0.0461236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1887_n 0.00359646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1888_n 0.0081372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1889_n 0.00359922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1890_n 0.0149258f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1891_n 0.0190181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1892_n 0.0226378f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1893_n 0.0190731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1894_n 0.00503395f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1895_n 0.00804943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1896_n 0.00960885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1897_n 0.00359922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1869_n 0.0663855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_A_700_389#_c_2078_n 0.0104469f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.202
cc_258 VPB N_A_700_389#_c_2086_n 0.00736664f $X=-0.19 $Y=1.305 $X2=0.315
+ $Y2=1.53
cc_259 VPB N_A_700_389#_c_2079_n 0.0263997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_A_1324_413#_c_2177_n 0.00289658f $X=-0.19 $Y=1.305 $X2=0.15
+ $Y2=1.445
cc_261 VPB N_A_1324_413#_c_2178_n 0.00261635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_A_1324_413#_c_2179_n 0.0024674f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.202
cc_263 VPB N_Q_c_2212_n 0.00151409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB Q 0.00159485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 CLK N_A_27_47#_M1016_s 0.00851196f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_266 N_CLK_c_269_n N_A_27_47#_c_297_n 0.0313045f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_267 CLK N_A_27_47#_c_297_n 5.57114e-19 $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_268 N_CLK_c_268_n N_A_27_47#_c_297_n 0.0245391f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_269 N_CLK_c_266_n N_A_27_47#_c_298_n 0.0185834f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_270 N_CLK_c_266_n N_A_27_47#_c_334_n 0.0142201f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_271 CLK N_A_27_47#_c_334_n 0.00950472f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_272 N_CLK_c_268_n N_A_27_47#_c_334_n 5.397e-19 $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_273 CLK N_A_27_47#_c_307_n 0.0181733f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_274 N_CLK_c_268_n N_A_27_47#_c_307_n 0.00296057f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_275 N_CLK_c_269_n N_A_27_47#_c_339_n 0.0142887f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_276 CLK N_A_27_47#_c_339_n 0.00647421f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_277 N_CLK_c_269_n N_A_27_47#_c_325_n 0.005471f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_278 CLK N_A_27_47#_c_326_n 0.0183116f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_279 N_CLK_c_268_n N_A_27_47#_c_326_n 0.00205709f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_280 CLK N_A_27_47#_c_344_n 0.00133464f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_281 N_CLK_c_268_n N_A_27_47#_c_314_n 0.00351882f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_282 N_CLK_c_266_n N_A_27_47#_c_317_n 0.00351882f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_283 CLK N_A_27_47#_c_317_n 0.0398976f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_284 N_CLK_c_269_n N_VPWR_c_1870_n 0.0128364f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_285 N_CLK_c_269_n N_VPWR_c_1890_n 0.00367409f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_286 N_CLK_c_269_n N_VPWR_c_1869_n 0.00529727f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_287 N_CLK_c_266_n N_VGND_c_2266_n 0.00198377f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_288 N_CLK_c_266_n N_VGND_c_2271_n 0.0142867f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_289 N_CLK_c_266_n N_VGND_c_2275_n 0.00367064f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_308_n N_A_331_66#_c_565_n 0.00129888f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_308_n N_A_331_66#_c_567_n 0.00161225f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_308_n N_A_331_66#_c_568_n 0.00846126f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_308_n N_A_331_66#_c_569_n 0.0012622f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_308_n N_A_331_66#_c_579_n 0.0126167f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_308_n N_A_331_66#_c_570_n 0.0369242f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_308_n N_A_331_66#_c_571_n 0.0230746f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_308_n N_A_331_66#_c_575_n 0.0145812f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_308_n N_A_331_66#_c_576_n 0.00210964f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_308_n N_D_M1008_g 0.0110765f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_308_n D 0.0121923f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_308_n N_SCE_M1040_g 0.00137541f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_308_n N_SCE_c_760_n 0.00256503f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_308_n N_SCE_c_763_n 0.00167851f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_308_n N_SCE_c_755_n 0.00556381f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_297_n N_SCE_c_756_n 0.00765345f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_308_n N_SCE_c_756_n 0.00152301f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_308_n N_SCE_c_757_n 0.00185197f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_308_n N_SCE_c_767_n 2.97081e-19 $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_309 N_A_27_47#_c_308_n SCE 0.0337825f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_310 N_A_27_47#_c_300_n N_SCD_M1038_g 0.00608596f $X=5.72 $Y=0.745 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_308_n N_SCD_M1038_g 0.00493204f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_312 N_A_27_47#_c_315_n N_SCD_M1038_g 0.0106705f $X=5.565 $Y=1.23 $X2=0 $Y2=0
cc_313 N_A_27_47#_c_308_n SCD 0.0340088f $X=5.42 $Y=1.19 $X2=0 $Y2=0
cc_314 N_A_27_47#_c_301_n N_A_213_47#_c_904_n 0.0243425f $X=6.43 $Y=1.32 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_320_n N_A_213_47#_c_904_n 0.0139619f $X=6.53 $Y=1.89 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_321_n N_A_213_47#_c_904_n 0.0107746f $X=6.53 $Y=1.99 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_309_n N_A_213_47#_c_904_n 2.02719e-19 $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_302_n N_A_213_47#_c_894_n 0.0139156f $X=5.985 $Y=0.67 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_M1027_g N_A_213_47#_c_895_n 0.0135694f $X=9.255 $Y=0.415 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_322_n N_A_213_47#_c_905_n 0.0210549f $X=9.185 $Y=1.89 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_323_n N_A_213_47#_c_905_n 0.0165347f $X=9.185 $Y=1.99 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_299_n N_A_213_47#_c_896_n 0.0110357f $X=5.91 $Y=0.745 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_316_n N_A_213_47#_c_896_n 0.00185495f $X=5.562 $Y=1.065
+ $X2=0 $Y2=0
cc_324 N_A_27_47#_c_301_n N_A_213_47#_c_897_n 0.00591483f $X=6.43 $Y=1.32 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_309_n N_A_213_47#_c_897_n 0.019051f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_M1027_g N_A_213_47#_c_898_n 0.00239394f $X=9.255 $Y=0.415
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_304_n N_A_213_47#_c_898_n 0.00739585f $X=9.27 $Y=1.37 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_305_n N_A_213_47#_c_898_n 0.003844f $X=9.317 $Y=1.082 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_309_n N_A_213_47#_c_898_n 0.0177781f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_311_n N_A_213_47#_c_898_n 0.00254889f $X=9.32 $Y=1.19 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_313_n N_A_213_47#_c_898_n 0.0183482f $X=9.32 $Y=1.11 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_M1027_g N_A_213_47#_c_899_n 0.0215319f $X=9.255 $Y=0.415 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_309_n N_A_213_47#_c_899_n 5.39192e-19 $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_313_n N_A_213_47#_c_899_n 3.70541e-19 $X=9.32 $Y=1.11 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_322_n N_A_213_47#_c_907_n 0.00731249f $X=9.185 $Y=1.89 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_309_n N_A_213_47#_c_907_n 0.00491017f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_311_n N_A_213_47#_c_907_n 7.60662e-19 $X=9.32 $Y=1.19 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_297_n N_A_213_47#_c_900_n 2.07055e-19 $X=0.98 $Y=1.41 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_308_n N_A_213_47#_c_900_n 0.00291916f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_297_n N_A_213_47#_c_908_n 0.00608776f $X=0.98 $Y=1.41 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_339_n N_A_213_47#_c_908_n 0.00869622f $X=0.71 $Y=1.88 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_325_n N_A_213_47#_c_908_n 0.00335166f $X=0.812 $Y=1.795
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_c_308_n N_A_213_47#_c_908_n 0.00159908f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_297_n N_A_213_47#_c_901_n 0.0123414f $X=0.98 $Y=1.41 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_298_n N_A_213_47#_c_901_n 0.0064f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_325_n N_A_213_47#_c_901_n 0.0198217f $X=0.812 $Y=1.795 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_308_n N_A_213_47#_c_901_n 0.0192858f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_344_n N_A_213_47#_c_901_n 0.00240264f $X=1.085 $Y=1.19 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_314_n N_A_213_47#_c_901_n 0.0226049f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_317_n N_A_213_47#_c_901_n 0.0072771f $X=0.867 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_322_n N_A_213_47#_c_910_n 0.0119565f $X=9.185 $Y=1.89 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_323_n N_A_213_47#_c_910_n 0.00281153f $X=9.185 $Y=1.99 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_304_n N_A_213_47#_c_910_n 0.00498488f $X=9.27 $Y=1.37 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_311_n N_A_213_47#_c_910_n 0.00364468f $X=9.32 $Y=1.19 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_313_n N_A_213_47#_c_910_n 0.011998f $X=9.32 $Y=1.11 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_308_n N_A_213_47#_c_911_n 0.180893f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_309_n N_A_213_47#_c_911_n 0.00796825f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_416_p N_A_213_47#_c_911_n 0.014344f $X=5.71 $Y=1.19 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_310_n N_A_213_47#_c_911_n 0.0016551f $X=5.565 $Y=1.19 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_315_n N_A_213_47#_c_911_n 0.0025783f $X=5.565 $Y=1.23 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_297_n N_A_213_47#_c_912_n 0.00108537f $X=0.98 $Y=1.41 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_339_n N_A_213_47#_c_912_n 0.00584013f $X=0.71 $Y=1.88 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_325_n N_A_213_47#_c_912_n 0.00114159f $X=0.812 $Y=1.795
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_c_308_n N_A_213_47#_c_912_n 0.0128994f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_344_n N_A_213_47#_c_912_n 8.4505e-19 $X=1.085 $Y=1.19 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_301_n N_A_213_47#_c_913_n 0.00132845f $X=6.43 $Y=1.32 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_320_n N_A_213_47#_c_913_n 0.00262632f $X=6.53 $Y=1.89 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_321_n N_A_213_47#_c_913_n 0.00308437f $X=6.53 $Y=1.99 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_322_n N_A_213_47#_c_913_n 0.0015364f $X=9.185 $Y=1.89 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_323_n N_A_213_47#_c_913_n 0.00196843f $X=9.185 $Y=1.99 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_309_n N_A_213_47#_c_913_n 0.126539f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_311_n N_A_213_47#_c_913_n 0.013738f $X=9.32 $Y=1.19 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_313_n N_A_213_47#_c_913_n 3.77496e-19 $X=9.32 $Y=1.11 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_301_n N_A_213_47#_c_914_n 7.57971e-19 $X=6.43 $Y=1.32 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_309_n N_A_213_47#_c_914_n 0.0128756f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_323_n N_A_213_47#_c_916_n 4.6329e-19 $X=9.185 $Y=1.99 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_301_n N_A_213_47#_c_917_n 0.00183386f $X=6.43 $Y=1.32 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_c_320_n N_A_213_47#_c_917_n 4.98483e-19 $X=6.53 $Y=1.89 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_309_n N_A_213_47#_c_917_n 0.00224066f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_299_n N_A_213_47#_c_902_n 0.00668438f $X=5.91 $Y=0.745 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_301_n N_A_213_47#_c_902_n 0.0205795f $X=6.43 $Y=1.32 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_309_n N_A_213_47#_c_902_n 0.00438155f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_316_n N_A_213_47#_c_902_n 0.00171454f $X=5.562 $Y=1.065
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_322_n N_A_213_47#_c_918_n 2.44676e-19 $X=9.185 $Y=1.89 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_304_n N_A_213_47#_c_918_n 3.61623e-19 $X=9.27 $Y=1.37 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_311_n N_A_213_47#_c_918_n 5.34355e-19 $X=9.32 $Y=1.19 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_301_n N_A_213_47#_c_903_n 0.0133665f $X=6.43 $Y=1.32 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_320_n N_A_213_47#_c_903_n 0.00107722f $X=6.53 $Y=1.89 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_309_n N_A_213_47#_c_903_n 0.0215044f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_416_p N_A_213_47#_c_903_n 0.0022665f $X=5.71 $Y=1.19 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_310_n N_A_213_47#_c_903_n 0.0150534f $X=5.565 $Y=1.19 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_316_n N_A_213_47#_c_903_n 0.00254035f $X=5.562 $Y=1.065
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_320_n N_A_1380_303#_c_1149_n 0.023475f $X=6.53 $Y=1.89 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_321_n N_A_1380_303#_c_1149_n 0.0125938f $X=6.53 $Y=1.99
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_301_n N_A_1380_303#_M1000_g 0.00931633f $X=6.43 $Y=1.32
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_c_309_n N_A_1380_303#_M1000_g 0.00614226f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_320_n N_A_1380_303#_c_1151_n 5.8087e-19 $X=6.53 $Y=1.89
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_c_309_n N_A_1380_303#_c_1151_n 0.0059501f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_322_n N_A_1380_303#_c_1160_n 0.00180498f $X=9.185 $Y=1.89
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_323_n N_A_1380_303#_c_1160_n 4.15787e-19 $X=9.185 $Y=1.99
+ $X2=0 $Y2=0
cc_401 N_A_27_47#_c_309_n N_A_1380_303#_c_1160_n 0.00195566f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_323_n N_A_1380_303#_c_1163_n 0.00372111f $X=9.185 $Y=1.99
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_309_n N_A_1380_303#_c_1164_n 0.0015131f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_c_309_n N_A_1380_303#_c_1152_n 0.00397493f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_M1027_g N_A_1380_303#_c_1148_n 4.94982e-19 $X=9.255 $Y=0.415
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_309_n N_A_1380_303#_c_1148_n 0.0130718f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_309_n N_RESET_B_c_1255_n 0.00116052f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_c_309_n N_RESET_B_c_1258_n 0.0691234f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_409 N_A_27_47#_c_309_n N_RESET_B_c_1259_n 0.00371083f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_410 N_A_27_47#_M1027_g N_RESET_B_c_1260_n 0.00490692f $X=9.255 $Y=0.415 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_c_304_n N_RESET_B_c_1260_n 4.42407e-19 $X=9.27 $Y=1.37 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_c_305_n N_RESET_B_c_1260_n 8.9785e-19 $X=9.317 $Y=1.082 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_309_n N_RESET_B_c_1260_n 0.0992198f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_c_311_n N_RESET_B_c_1260_n 0.0279502f $X=9.32 $Y=1.19 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_313_n N_RESET_B_c_1260_n 0.00217385f $X=9.32 $Y=1.11 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_309_n N_RESET_B_c_1264_n 0.00296898f $X=9.155 $Y=1.19 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_322_n N_A_1202_413#_c_1429_n 0.0053475f $X=9.185 $Y=1.89
+ $X2=0 $Y2=0
cc_418 N_A_27_47#_c_309_n N_A_1202_413#_c_1429_n 0.00331303f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_419 N_A_27_47#_c_322_n N_A_1202_413#_c_1430_n 0.0151115f $X=9.185 $Y=1.89
+ $X2=0 $Y2=0
cc_420 N_A_27_47#_c_323_n N_A_1202_413#_c_1430_n 0.008324f $X=9.185 $Y=1.99
+ $X2=0 $Y2=0
cc_421 N_A_27_47#_c_301_n N_A_1202_413#_c_1423_n 0.00826718f $X=6.43 $Y=1.32
+ $X2=0 $Y2=0
cc_422 N_A_27_47#_c_309_n N_A_1202_413#_c_1423_n 0.0146704f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_423 N_A_27_47#_c_301_n N_A_1202_413#_c_1424_n 0.00451282f $X=6.43 $Y=1.32
+ $X2=0 $Y2=0
cc_424 N_A_27_47#_c_309_n N_A_1202_413#_c_1424_n 0.00696389f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_c_309_n N_A_1202_413#_c_1425_n 0.0164556f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_c_309_n N_A_1202_413#_c_1426_n 0.0304996f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_427 N_A_27_47#_c_321_n N_A_1202_413#_c_1447_n 0.00476736f $X=6.53 $Y=1.99
+ $X2=0 $Y2=0
cc_428 N_A_27_47#_c_301_n N_A_1202_413#_c_1433_n 0.0037409f $X=6.43 $Y=1.32
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_320_n N_A_1202_413#_c_1433_n 0.0154505f $X=6.53 $Y=1.89
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_321_n N_A_1202_413#_c_1433_n 0.00605858f $X=6.53 $Y=1.99
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_c_309_n N_A_1202_413#_c_1434_n 0.00403101f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_c_309_n N_A_1202_413#_c_1427_n 0.0113465f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_309_n N_A_1202_413#_c_1428_n 0.00568294f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_M1027_g N_A_1972_21#_M1032_g 0.0156688f $X=9.255 $Y=0.415
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_312_n N_A_1972_21#_c_1562_n 0.00277252f $X=9.32 $Y=1.11
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_305_n N_A_1972_21#_c_1578_n 0.00328316f $X=9.317 $Y=1.082
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_M1027_g N_A_1757_47#_c_1764_n 0.0174239f $X=9.255 $Y=0.415
+ $X2=0 $Y2=0
cc_438 N_A_27_47#_c_305_n N_A_1757_47#_c_1764_n 0.0018711f $X=9.317 $Y=1.082
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_c_313_n N_A_1757_47#_c_1764_n 0.00351567f $X=9.32 $Y=1.11
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_323_n N_A_1757_47#_c_1767_n 0.00724953f $X=9.185 $Y=1.99
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_M1027_g N_A_1757_47#_c_1757_n 0.00675244f $X=9.255 $Y=0.415
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_c_305_n N_A_1757_47#_c_1757_n 0.00325626f $X=9.317 $Y=1.082
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_c_311_n N_A_1757_47#_c_1757_n 0.00735413f $X=9.32 $Y=1.19
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_313_n N_A_1757_47#_c_1757_n 0.0177077f $X=9.32 $Y=1.11 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_c_322_n N_A_1757_47#_c_1762_n 0.00377614f $X=9.185 $Y=1.89
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_304_n N_A_1757_47#_c_1762_n 0.00144767f $X=9.27 $Y=1.37
+ $X2=0 $Y2=0
cc_447 N_A_27_47#_c_313_n N_A_1757_47#_c_1762_n 5.75024e-19 $X=9.32 $Y=1.11
+ $X2=0 $Y2=0
cc_448 N_A_27_47#_c_339_n N_VPWR_M1016_d 0.0045758f $X=0.71 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_449 N_A_27_47#_c_325_n N_VPWR_M1016_d 0.00323704f $X=0.812 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_450 N_A_27_47#_c_297_n N_VPWR_c_1870_n 0.0108218f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_451 N_A_27_47#_c_339_n N_VPWR_c_1870_n 0.0214591f $X=0.71 $Y=1.88 $X2=0 $Y2=0
cc_452 N_A_27_47#_c_326_n N_VPWR_c_1870_n 0.0237818f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_453 N_A_27_47#_c_297_n N_VPWR_c_1880_n 0.00618803f $X=0.98 $Y=1.41 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_321_n N_VPWR_c_1885_n 0.00696599f $X=6.53 $Y=1.99 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_323_n N_VPWR_c_1886_n 0.00601827f $X=9.185 $Y=1.99 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_339_n N_VPWR_c_1890_n 0.0019892f $X=0.71 $Y=1.88 $X2=0 $Y2=0
cc_457 N_A_27_47#_c_326_n N_VPWR_c_1890_n 0.0178321f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_458 N_A_27_47#_M1016_s N_VPWR_c_1869_n 0.00248688f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_297_n N_VPWR_c_1869_n 0.0114979f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_460 N_A_27_47#_c_321_n N_VPWR_c_1869_n 0.00784451f $X=6.53 $Y=1.99 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_323_n N_VPWR_c_1869_n 0.00710573f $X=9.185 $Y=1.99 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_339_n N_VPWR_c_1869_n 0.00570194f $X=0.71 $Y=1.88 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_326_n N_VPWR_c_1869_n 0.00973967f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_308_n N_A_700_389#_c_2078_n 0.0148988f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_c_308_n N_A_700_389#_c_2079_n 0.0135421f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_c_416_p N_A_700_389#_c_2079_n 0.00240264f $X=5.71 $Y=1.19
+ $X2=0 $Y2=0
cc_467 N_A_27_47#_c_310_n N_A_700_389#_c_2079_n 0.0252651f $X=5.565 $Y=1.19
+ $X2=0 $Y2=0
cc_468 N_A_27_47#_c_315_n N_A_700_389#_c_2079_n 0.00500788f $X=5.565 $Y=1.23
+ $X2=0 $Y2=0
cc_469 N_A_27_47#_c_316_n N_A_700_389#_c_2079_n 0.0017755f $X=5.562 $Y=1.065
+ $X2=0 $Y2=0
cc_470 N_A_27_47#_c_300_n N_A_700_389#_c_2080_n 0.00472302f $X=5.72 $Y=0.745
+ $X2=0 $Y2=0
cc_471 N_A_27_47#_c_308_n N_A_700_389#_c_2080_n 0.00466124f $X=5.42 $Y=1.19
+ $X2=0 $Y2=0
cc_472 N_A_27_47#_c_309_n N_A_700_389#_c_2080_n 3.78682e-19 $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_473 N_A_27_47#_c_416_p N_A_700_389#_c_2080_n 0.00657764f $X=5.71 $Y=1.19
+ $X2=0 $Y2=0
cc_474 N_A_27_47#_c_310_n N_A_700_389#_c_2080_n 0.0116936f $X=5.565 $Y=1.19
+ $X2=0 $Y2=0
cc_475 N_A_27_47#_c_315_n N_A_700_389#_c_2080_n 0.00350952f $X=5.565 $Y=1.23
+ $X2=0 $Y2=0
cc_476 N_A_27_47#_c_316_n N_A_700_389#_c_2080_n 0.00555216f $X=5.562 $Y=1.065
+ $X2=0 $Y2=0
cc_477 N_A_27_47#_c_300_n N_A_700_389#_c_2082_n 0.0051054f $X=5.72 $Y=0.745
+ $X2=0 $Y2=0
cc_478 N_A_27_47#_c_302_n N_A_700_389#_c_2082_n 0.00402367f $X=5.985 $Y=0.67
+ $X2=0 $Y2=0
cc_479 N_A_27_47#_c_308_n N_A_700_389#_c_2083_n 0.0135597f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_c_300_n N_A_700_389#_c_2084_n 0.0059572f $X=5.72 $Y=0.745
+ $X2=0 $Y2=0
cc_481 N_A_27_47#_c_309_n N_A_700_389#_c_2084_n 0.00509945f $X=9.155 $Y=1.19
+ $X2=0 $Y2=0
cc_482 N_A_27_47#_c_321_n N_A_1324_413#_c_2178_n 0.00209945f $X=6.53 $Y=1.99
+ $X2=0 $Y2=0
cc_483 N_A_27_47#_c_334_n N_VGND_M1031_d 0.00511432f $X=0.71 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_484 N_A_27_47#_c_317_n N_VGND_M1031_d 9.31974e-19 $X=0.867 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_485 N_A_27_47#_c_308_n N_VGND_c_2249_n 5.94768e-19 $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_c_308_n N_VGND_c_2250_n 0.00240425f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_c_302_n N_VGND_c_2251_n 0.0035082f $X=5.985 $Y=0.67 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_308_n N_VGND_c_2251_n 0.00519614f $X=5.42 $Y=1.19 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_c_299_n N_VGND_c_2258_n 4.41192e-19 $X=5.91 $Y=0.745 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_c_302_n N_VGND_c_2258_n 0.00434697f $X=5.985 $Y=0.67 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_M1027_g N_VGND_c_2260_n 0.00357877f $X=9.255 $Y=0.415 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_306_n N_VGND_c_2266_n 0.0107551f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_493 N_A_27_47#_c_334_n N_VGND_c_2266_n 0.00244154f $X=0.71 $Y=0.72 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_c_298_n N_VGND_c_2267_n 0.00585385f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_c_297_n N_VGND_c_2271_n 2.49184e-19 $X=0.98 $Y=1.41 $X2=0
+ $Y2=0
cc_496 N_A_27_47#_c_298_n N_VGND_c_2271_n 0.00317372f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_c_306_n N_VGND_c_2271_n 0.00921779f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_498 N_A_27_47#_c_334_n N_VGND_c_2271_n 0.0223403f $X=0.71 $Y=0.72 $X2=0 $Y2=0
cc_499 N_A_27_47#_c_344_n N_VGND_c_2271_n 3.83259e-19 $X=1.085 $Y=1.19 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_M1031_s N_VGND_c_2275_n 0.00296179f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_501 N_A_27_47#_c_298_n N_VGND_c_2275_n 0.0120602f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_502 N_A_27_47#_c_299_n N_VGND_c_2275_n 4.24653e-19 $X=5.91 $Y=0.745 $X2=0
+ $Y2=0
cc_503 N_A_27_47#_c_302_n N_VGND_c_2275_n 0.00765378f $X=5.985 $Y=0.67 $X2=0
+ $Y2=0
cc_504 N_A_27_47#_M1027_g N_VGND_c_2275_n 0.00608701f $X=9.255 $Y=0.415 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_c_306_n N_VGND_c_2275_n 0.00898615f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_c_334_n N_VGND_c_2275_n 0.00619727f $X=0.71 $Y=0.72 $X2=0
+ $Y2=0
cc_507 N_A_331_66#_c_567_n N_D_c_709_n 0.00995544f $X=4.26 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_508 N_A_331_66#_c_579_n N_D_c_709_n 8.93785e-19 $X=2.645 $Y=1.29 $X2=-0.19
+ $Y2=-0.24
cc_509 N_A_331_66#_c_570_n N_D_c_709_n 6.9685e-19 $X=3.275 $Y=1.09 $X2=-0.19
+ $Y2=-0.24
cc_510 N_A_331_66#_c_566_n N_D_M1008_g 0.0257211f $X=3.08 $Y=1.09 $X2=0 $Y2=0
cc_511 N_A_331_66#_c_567_n N_D_M1008_g 0.00677732f $X=4.26 $Y=1.87 $X2=0 $Y2=0
cc_512 N_A_331_66#_c_570_n N_D_M1008_g 0.00210251f $X=3.275 $Y=1.09 $X2=0 $Y2=0
cc_513 N_A_331_66#_c_572_n N_D_M1008_g 0.00525772f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_514 N_A_331_66#_c_573_n N_D_M1008_g 0.0037178f $X=4.265 $Y=0.34 $X2=0 $Y2=0
cc_515 N_A_331_66#_c_575_n N_D_M1008_g 0.00131275f $X=4.35 $Y=1.52 $X2=0 $Y2=0
cc_516 N_A_331_66#_c_576_n N_D_M1008_g 0.00352384f $X=2.62 $Y=1.165 $X2=0 $Y2=0
cc_517 N_A_331_66#_c_565_n D 7.28113e-19 $X=3.005 $Y=1.165 $X2=0 $Y2=0
cc_518 N_A_331_66#_c_567_n D 0.00118937f $X=4.26 $Y=1.87 $X2=0 $Y2=0
cc_519 N_A_331_66#_c_578_n D 0.00431835f $X=2.602 $Y=1.915 $X2=0 $Y2=0
cc_520 N_A_331_66#_c_579_n D 0.0239294f $X=2.645 $Y=1.29 $X2=0 $Y2=0
cc_521 N_A_331_66#_c_570_n D 0.0236451f $X=3.275 $Y=1.09 $X2=0 $Y2=0
cc_522 N_A_331_66#_c_576_n D 7.81926e-19 $X=2.62 $Y=1.165 $X2=0 $Y2=0
cc_523 N_A_331_66#_c_568_n N_SCE_M1040_g 0.0145383f $X=2.265 $Y=0.815 $X2=0
+ $Y2=0
cc_524 N_A_331_66#_c_571_n N_SCE_M1040_g 0.00748807f $X=2.73 $Y=1.09 $X2=0 $Y2=0
cc_525 N_A_331_66#_c_576_n N_SCE_M1040_g 0.0137273f $X=2.62 $Y=1.165 $X2=0 $Y2=0
cc_526 N_A_331_66#_c_566_n N_SCE_c_753_n 0.0102879f $X=3.08 $Y=1.09 $X2=0 $Y2=0
cc_527 N_A_331_66#_c_568_n N_SCE_c_753_n 2.18848e-19 $X=2.265 $Y=0.815 $X2=0
+ $Y2=0
cc_528 N_A_331_66#_c_571_n N_SCE_c_753_n 9.65915e-19 $X=2.73 $Y=1.09 $X2=0 $Y2=0
cc_529 N_A_331_66#_c_573_n N_SCE_c_753_n 0.00975092f $X=4.265 $Y=0.34 $X2=0
+ $Y2=0
cc_530 N_A_331_66#_c_574_n N_SCE_c_753_n 0.00420304f $X=3.445 $Y=0.34 $X2=0
+ $Y2=0
cc_531 N_A_331_66#_c_571_n N_SCE_c_760_n 0.0035177f $X=2.73 $Y=1.09 $X2=0 $Y2=0
cc_532 N_A_331_66#_c_578_n N_SCE_c_761_n 0.00893431f $X=2.602 $Y=1.915 $X2=0
+ $Y2=0
cc_533 N_A_331_66#_c_578_n N_SCE_c_762_n 0.010859f $X=2.602 $Y=1.915 $X2=0 $Y2=0
cc_534 N_A_331_66#_c_579_n N_SCE_c_762_n 0.00165355f $X=2.645 $Y=1.29 $X2=0
+ $Y2=0
cc_535 N_A_331_66#_c_565_n N_SCE_c_763_n 0.00935155f $X=3.005 $Y=1.165 $X2=0
+ $Y2=0
cc_536 N_A_331_66#_c_578_n N_SCE_c_763_n 5.67231e-19 $X=2.602 $Y=1.915 $X2=0
+ $Y2=0
cc_537 N_A_331_66#_c_579_n N_SCE_c_763_n 0.00714807f $X=2.645 $Y=1.29 $X2=0
+ $Y2=0
cc_538 N_A_331_66#_c_570_n N_SCE_c_763_n 0.00315696f $X=3.275 $Y=1.09 $X2=0
+ $Y2=0
cc_539 N_A_331_66#_c_578_n N_SCE_c_764_n 0.00154869f $X=2.602 $Y=1.915 $X2=0
+ $Y2=0
cc_540 N_A_331_66#_c_579_n N_SCE_c_764_n 2.87199e-19 $X=2.645 $Y=1.29 $X2=0
+ $Y2=0
cc_541 N_A_331_66#_c_567_n N_SCE_c_755_n 0.00892078f $X=4.26 $Y=1.87 $X2=0 $Y2=0
cc_542 N_A_331_66#_c_572_n N_SCE_c_755_n 0.00167135f $X=3.36 $Y=0.995 $X2=0
+ $Y2=0
cc_543 N_A_331_66#_c_573_n N_SCE_c_755_n 0.0258097f $X=4.265 $Y=0.34 $X2=0 $Y2=0
cc_544 N_A_331_66#_c_575_n N_SCE_c_755_n 0.0240247f $X=4.35 $Y=1.52 $X2=0 $Y2=0
cc_545 N_A_331_66#_c_568_n N_SCE_c_756_n 5.71498e-19 $X=2.265 $Y=0.815 $X2=0
+ $Y2=0
cc_546 N_A_331_66#_c_569_n N_SCE_c_756_n 0.00107346f $X=1.865 $Y=0.815 $X2=0
+ $Y2=0
cc_547 N_A_331_66#_c_579_n N_SCE_c_757_n 0.00135957f $X=2.645 $Y=1.29 $X2=0
+ $Y2=0
cc_548 N_A_331_66#_c_578_n N_SCE_c_767_n 4.44592e-19 $X=2.602 $Y=1.915 $X2=0
+ $Y2=0
cc_549 N_A_331_66#_c_579_n N_SCE_c_767_n 0.0109362f $X=2.645 $Y=1.29 $X2=0 $Y2=0
cc_550 N_A_331_66#_c_571_n N_SCE_c_767_n 3.29459e-19 $X=2.73 $Y=1.09 $X2=0 $Y2=0
cc_551 N_A_331_66#_c_576_n N_SCE_c_767_n 0.0249164f $X=2.62 $Y=1.165 $X2=0 $Y2=0
cc_552 N_A_331_66#_c_568_n SCE 0.0136696f $X=2.265 $Y=0.815 $X2=0 $Y2=0
cc_553 N_A_331_66#_c_569_n SCE 0.0143043f $X=1.865 $Y=0.815 $X2=0 $Y2=0
cc_554 N_A_331_66#_c_578_n SCE 0.00721995f $X=2.602 $Y=1.915 $X2=0 $Y2=0
cc_555 N_A_331_66#_c_579_n SCE 0.028953f $X=2.645 $Y=1.29 $X2=0 $Y2=0
cc_556 N_A_331_66#_c_571_n SCE 0.00523341f $X=2.73 $Y=1.09 $X2=0 $Y2=0
cc_557 N_A_331_66#_c_576_n SCE 0.00140593f $X=2.62 $Y=1.165 $X2=0 $Y2=0
cc_558 N_A_331_66#_c_567_n N_SCD_c_857_n 0.0528131f $X=4.26 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_559 N_A_331_66#_c_575_n N_SCD_c_857_n 2.98757e-19 $X=4.35 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_560 N_A_331_66#_c_567_n N_SCD_M1038_g 8.4866e-19 $X=4.26 $Y=1.87 $X2=0 $Y2=0
cc_561 N_A_331_66#_c_573_n N_SCD_M1038_g 6.01506e-19 $X=4.265 $Y=0.34 $X2=0
+ $Y2=0
cc_562 N_A_331_66#_c_575_n N_SCD_M1038_g 0.00327141f $X=4.35 $Y=1.52 $X2=0 $Y2=0
cc_563 N_A_331_66#_c_567_n SCD 0.00242948f $X=4.26 $Y=1.87 $X2=0 $Y2=0
cc_564 N_A_331_66#_c_575_n SCD 0.0730534f $X=4.35 $Y=1.52 $X2=0 $Y2=0
cc_565 N_A_331_66#_c_648_p N_A_213_47#_c_900_n 0.0157971f $X=1.78 $Y=0.56 $X2=0
+ $Y2=0
cc_566 N_A_331_66#_c_569_n N_A_213_47#_c_901_n 0.00901517f $X=1.865 $Y=0.815
+ $X2=0 $Y2=0
cc_567 N_A_331_66#_c_565_n N_A_213_47#_c_911_n 3.39815e-19 $X=3.005 $Y=1.165
+ $X2=0 $Y2=0
cc_568 N_A_331_66#_c_567_n N_A_213_47#_c_911_n 0.0076472f $X=4.26 $Y=1.87 $X2=0
+ $Y2=0
cc_569 N_A_331_66#_c_652_p N_A_213_47#_c_911_n 5.2445e-19 $X=2.295 $Y=2.22 $X2=0
+ $Y2=0
cc_570 N_A_331_66#_c_578_n N_A_213_47#_c_911_n 0.0204297f $X=2.602 $Y=1.915
+ $X2=0 $Y2=0
cc_571 N_A_331_66#_c_579_n N_A_213_47#_c_911_n 0.0155308f $X=2.645 $Y=1.29 $X2=0
+ $Y2=0
cc_572 N_A_331_66#_c_570_n N_A_213_47#_c_911_n 0.00425452f $X=3.275 $Y=1.09
+ $X2=0 $Y2=0
cc_573 N_A_331_66#_c_575_n N_A_213_47#_c_911_n 0.00219668f $X=4.35 $Y=1.52 $X2=0
+ $Y2=0
cc_574 N_A_331_66#_c_578_n N_VPWR_M1030_d 0.00225972f $X=2.602 $Y=1.915 $X2=0
+ $Y2=0
cc_575 N_A_331_66#_c_652_p N_VPWR_c_1871_n 0.00909067f $X=2.295 $Y=2.22 $X2=0
+ $Y2=0
cc_576 N_A_331_66#_c_578_n N_VPWR_c_1871_n 0.00496417f $X=2.602 $Y=1.915 $X2=0
+ $Y2=0
cc_577 N_A_331_66#_c_567_n N_VPWR_c_1872_n 0.00186755f $X=4.26 $Y=1.87 $X2=0
+ $Y2=0
cc_578 N_A_331_66#_c_652_p N_VPWR_c_1880_n 0.0125789f $X=2.295 $Y=2.22 $X2=0
+ $Y2=0
cc_579 N_A_331_66#_c_578_n N_VPWR_c_1880_n 0.00324706f $X=2.602 $Y=1.915 $X2=0
+ $Y2=0
cc_580 N_A_331_66#_c_567_n N_VPWR_c_1882_n 0.00506535f $X=4.26 $Y=1.87 $X2=0
+ $Y2=0
cc_581 N_A_331_66#_M1030_s N_VPWR_c_1869_n 0.00352874f $X=2.03 $Y=1.945 $X2=0
+ $Y2=0
cc_582 N_A_331_66#_c_567_n N_VPWR_c_1869_n 0.00739028f $X=4.26 $Y=1.87 $X2=0
+ $Y2=0
cc_583 N_A_331_66#_c_652_p N_VPWR_c_1869_n 0.00452124f $X=2.295 $Y=2.22 $X2=0
+ $Y2=0
cc_584 N_A_331_66#_c_578_n N_VPWR_c_1869_n 0.00271653f $X=2.602 $Y=1.915 $X2=0
+ $Y2=0
cc_585 N_A_331_66#_c_573_n N_A_700_389#_M1008_d 0.00378915f $X=4.265 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_586 N_A_331_66#_c_567_n N_A_700_389#_c_2078_n 0.00943309f $X=4.26 $Y=1.87
+ $X2=0 $Y2=0
cc_587 N_A_331_66#_c_570_n N_A_700_389#_c_2078_n 0.00383918f $X=3.275 $Y=1.09
+ $X2=0 $Y2=0
cc_588 N_A_331_66#_c_575_n N_A_700_389#_c_2078_n 0.035943f $X=4.35 $Y=1.52 $X2=0
+ $Y2=0
cc_589 N_A_331_66#_c_567_n N_A_700_389#_c_2110_n 0.00929615f $X=4.26 $Y=1.87
+ $X2=0 $Y2=0
cc_590 N_A_331_66#_c_567_n N_A_700_389#_c_2086_n 0.0192266f $X=4.26 $Y=1.87
+ $X2=0 $Y2=0
cc_591 N_A_331_66#_c_575_n N_A_700_389#_c_2086_n 0.00723687f $X=4.35 $Y=1.52
+ $X2=0 $Y2=0
cc_592 N_A_331_66#_c_570_n N_A_700_389#_c_2083_n 0.00433315f $X=3.275 $Y=1.09
+ $X2=0 $Y2=0
cc_593 N_A_331_66#_c_573_n N_A_700_389#_c_2083_n 0.0165664f $X=4.265 $Y=0.34
+ $X2=0 $Y2=0
cc_594 N_A_331_66#_c_575_n N_A_700_389#_c_2083_n 0.0250741f $X=4.35 $Y=1.52
+ $X2=0 $Y2=0
cc_595 N_A_331_66#_c_568_n N_VGND_M1040_d 8.82396e-19 $X=2.265 $Y=0.815 $X2=0
+ $Y2=0
cc_596 N_A_331_66#_c_571_n N_VGND_M1040_d 0.00112204f $X=2.73 $Y=1.09 $X2=0
+ $Y2=0
cc_597 N_A_331_66#_c_570_n N_VGND_M1021_s 0.00231468f $X=3.275 $Y=1.09 $X2=0
+ $Y2=0
cc_598 N_A_331_66#_c_571_n N_VGND_M1021_s 3.87318e-19 $X=2.73 $Y=1.09 $X2=0
+ $Y2=0
cc_599 N_A_331_66#_c_566_n N_VGND_c_2249_n 3.51546e-19 $X=3.08 $Y=1.09 $X2=0
+ $Y2=0
cc_600 N_A_331_66#_c_648_p N_VGND_c_2249_n 0.0123182f $X=1.78 $Y=0.56 $X2=0
+ $Y2=0
cc_601 N_A_331_66#_c_568_n N_VGND_c_2249_n 0.0125952f $X=2.265 $Y=0.815 $X2=0
+ $Y2=0
cc_602 N_A_331_66#_c_571_n N_VGND_c_2249_n 0.0122579f $X=2.73 $Y=1.09 $X2=0
+ $Y2=0
cc_603 N_A_331_66#_c_566_n N_VGND_c_2250_n 0.00772682f $X=3.08 $Y=1.09 $X2=0
+ $Y2=0
cc_604 N_A_331_66#_c_570_n N_VGND_c_2250_n 0.0185034f $X=3.275 $Y=1.09 $X2=0
+ $Y2=0
cc_605 N_A_331_66#_c_571_n N_VGND_c_2250_n 0.0134261f $X=2.73 $Y=1.09 $X2=0
+ $Y2=0
cc_606 N_A_331_66#_c_572_n N_VGND_c_2250_n 0.0232893f $X=3.36 $Y=0.995 $X2=0
+ $Y2=0
cc_607 N_A_331_66#_c_574_n N_VGND_c_2250_n 0.0119285f $X=3.445 $Y=0.34 $X2=0
+ $Y2=0
cc_608 N_A_331_66#_c_576_n N_VGND_c_2250_n 0.00205168f $X=2.62 $Y=1.165 $X2=0
+ $Y2=0
cc_609 N_A_331_66#_c_573_n N_VGND_c_2251_n 0.00499434f $X=4.265 $Y=0.34 $X2=0
+ $Y2=0
cc_610 N_A_331_66#_c_575_n N_VGND_c_2251_n 0.00303005f $X=4.35 $Y=1.52 $X2=0
+ $Y2=0
cc_611 N_A_331_66#_c_648_p N_VGND_c_2267_n 0.00604119f $X=1.78 $Y=0.56 $X2=0
+ $Y2=0
cc_612 N_A_331_66#_c_568_n N_VGND_c_2267_n 0.00196018f $X=2.265 $Y=0.815 $X2=0
+ $Y2=0
cc_613 N_A_331_66#_c_571_n N_VGND_c_2268_n 3.17207e-19 $X=2.73 $Y=1.09 $X2=0
+ $Y2=0
cc_614 N_A_331_66#_c_573_n N_VGND_c_2269_n 0.0635681f $X=4.265 $Y=0.34 $X2=0
+ $Y2=0
cc_615 N_A_331_66#_c_574_n N_VGND_c_2269_n 0.0115906f $X=3.445 $Y=0.34 $X2=0
+ $Y2=0
cc_616 N_A_331_66#_c_566_n N_VGND_c_2275_n 7.52198e-19 $X=3.08 $Y=1.09 $X2=0
+ $Y2=0
cc_617 N_A_331_66#_c_648_p N_VGND_c_2275_n 0.00591457f $X=1.78 $Y=0.56 $X2=0
+ $Y2=0
cc_618 N_A_331_66#_c_568_n N_VGND_c_2275_n 0.00497709f $X=2.265 $Y=0.815 $X2=0
+ $Y2=0
cc_619 N_A_331_66#_c_571_n N_VGND_c_2275_n 0.00112098f $X=2.73 $Y=1.09 $X2=0
+ $Y2=0
cc_620 N_A_331_66#_c_573_n N_VGND_c_2275_n 0.0328547f $X=4.265 $Y=0.34 $X2=0
+ $Y2=0
cc_621 N_A_331_66#_c_574_n N_VGND_c_2275_n 0.00576957f $X=3.445 $Y=0.34 $X2=0
+ $Y2=0
cc_622 N_A_331_66#_c_570_n A_631_119# 0.00247854f $X=3.275 $Y=1.09 $X2=-0.19
+ $Y2=-0.24
cc_623 N_A_331_66#_c_572_n A_631_119# 0.00640899f $X=3.36 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_624 N_D_M1008_g N_SCE_c_753_n 0.00882199f $X=3.54 $Y=0.805 $X2=0 $Y2=0
cc_625 N_D_c_709_n N_SCE_c_763_n 0.0153852f $X=3.41 $Y=1.87 $X2=0 $Y2=0
cc_626 D N_SCE_c_763_n 0.00279607f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_627 N_D_c_709_n N_SCE_c_764_n 0.041013f $X=3.41 $Y=1.87 $X2=0 $Y2=0
cc_628 D N_SCE_c_764_n 0.00273551f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_629 N_D_M1008_g N_SCE_c_755_n 0.010145f $X=3.54 $Y=0.805 $X2=0 $Y2=0
cc_630 D N_A_213_47#_c_911_n 0.041618f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_631 N_D_c_709_n N_VPWR_c_1871_n 0.0012639f $X=3.41 $Y=1.87 $X2=0 $Y2=0
cc_632 N_D_c_709_n N_VPWR_c_1882_n 0.00429201f $X=3.41 $Y=1.87 $X2=0 $Y2=0
cc_633 D N_VPWR_c_1882_n 0.0322181f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_634 N_D_c_709_n N_VPWR_c_1869_n 0.00661857f $X=3.41 $Y=1.87 $X2=0 $Y2=0
cc_635 D N_VPWR_c_1869_n 0.00938927f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_636 D A_618_389# 0.00113442f $X=3.355 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_637 D N_A_700_389#_M1020_d 0.0065739f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_638 N_D_c_709_n N_A_700_389#_c_2078_n 3.59695e-19 $X=3.41 $Y=1.87 $X2=0 $Y2=0
cc_639 N_D_M1008_g N_A_700_389#_c_2078_n 0.00795149f $X=3.54 $Y=0.805 $X2=0
+ $Y2=0
cc_640 D N_A_700_389#_c_2078_n 0.0388534f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_641 N_D_c_709_n N_A_700_389#_c_2110_n 0.0010492f $X=3.41 $Y=1.87 $X2=0 $Y2=0
cc_642 D N_A_700_389#_c_2110_n 0.0240011f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_643 N_D_M1008_g N_A_700_389#_c_2083_n 0.00148929f $X=3.54 $Y=0.805 $X2=0
+ $Y2=0
cc_644 N_D_c_709_n N_A_700_389#_c_2123_n 6.15237e-19 $X=3.41 $Y=1.87 $X2=0 $Y2=0
cc_645 D N_A_700_389#_c_2123_n 0.0125277f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_646 N_SCE_c_753_n N_SCD_M1038_g 0.0227157f $X=3.995 $Y=0.18 $X2=0 $Y2=0
cc_647 N_SCE_c_755_n SCD 0.00155807f $X=4.245 $Y=0.255 $X2=0 $Y2=0
cc_648 N_SCE_M1040_g N_A_213_47#_c_900_n 0.00107747f $X=2.04 $Y=0.54 $X2=0 $Y2=0
cc_649 N_SCE_c_761_n N_A_213_47#_c_908_n 0.00136539f $X=2.115 $Y=1.71 $X2=0
+ $Y2=0
cc_650 N_SCE_M1040_g N_A_213_47#_c_901_n 0.00457042f $X=2.04 $Y=0.54 $X2=0 $Y2=0
cc_651 N_SCE_c_759_n N_A_213_47#_c_901_n 4.28568e-19 $X=2.04 $Y=1.635 $X2=0
+ $Y2=0
cc_652 N_SCE_c_756_n N_A_213_47#_c_901_n 0.00273602f $X=1.965 $Y=1.31 $X2=0
+ $Y2=0
cc_653 SCE N_A_213_47#_c_901_n 0.0431784f $X=1.985 $Y=1.53 $X2=0 $Y2=0
cc_654 N_SCE_c_761_n N_A_213_47#_c_911_n 0.00863588f $X=2.115 $Y=1.71 $X2=0
+ $Y2=0
cc_655 N_SCE_c_762_n N_A_213_47#_c_911_n 7.28228e-19 $X=2.53 $Y=1.87 $X2=0 $Y2=0
cc_656 N_SCE_c_763_n N_A_213_47#_c_911_n 0.00579695f $X=2.9 $Y=1.71 $X2=0 $Y2=0
cc_657 N_SCE_c_764_n N_A_213_47#_c_911_n 0.00399739f $X=3 $Y=1.87 $X2=0 $Y2=0
cc_658 N_SCE_c_756_n N_A_213_47#_c_911_n 3.85459e-19 $X=1.965 $Y=1.31 $X2=0
+ $Y2=0
cc_659 N_SCE_c_767_n N_A_213_47#_c_911_n 0.00166507f $X=2.53 $Y=1.71 $X2=0 $Y2=0
cc_660 SCE N_A_213_47#_c_911_n 0.0234353f $X=1.985 $Y=1.53 $X2=0 $Y2=0
cc_661 N_SCE_c_761_n N_A_213_47#_c_912_n 7.16822e-19 $X=2.115 $Y=1.71 $X2=0
+ $Y2=0
cc_662 N_SCE_c_762_n N_VPWR_c_1871_n 0.0103635f $X=2.53 $Y=1.87 $X2=0 $Y2=0
cc_663 N_SCE_c_763_n N_VPWR_c_1871_n 0.00414019f $X=2.9 $Y=1.71 $X2=0 $Y2=0
cc_664 N_SCE_c_764_n N_VPWR_c_1871_n 0.00776205f $X=3 $Y=1.87 $X2=0 $Y2=0
cc_665 N_SCE_c_762_n N_VPWR_c_1880_n 0.00452725f $X=2.53 $Y=1.87 $X2=0 $Y2=0
cc_666 N_SCE_c_764_n N_VPWR_c_1882_n 0.00622633f $X=3 $Y=1.87 $X2=0 $Y2=0
cc_667 N_SCE_c_762_n N_VPWR_c_1869_n 0.00622226f $X=2.53 $Y=1.87 $X2=0 $Y2=0
cc_668 N_SCE_c_764_n N_VPWR_c_1869_n 0.00565321f $X=3 $Y=1.87 $X2=0 $Y2=0
cc_669 N_SCE_c_755_n N_A_700_389#_c_2078_n 2.17149e-19 $X=4.245 $Y=0.255 $X2=0
+ $Y2=0
cc_670 N_SCE_c_755_n N_A_700_389#_c_2083_n 0.00867384f $X=4.245 $Y=0.255 $X2=0
+ $Y2=0
cc_671 N_SCE_M1040_g N_VGND_c_2249_n 0.00911531f $X=2.04 $Y=0.54 $X2=0 $Y2=0
cc_672 N_SCE_c_753_n N_VGND_c_2249_n 0.0154857f $X=3.995 $Y=0.18 $X2=0 $Y2=0
cc_673 N_SCE_c_754_n N_VGND_c_2249_n 0.0056308f $X=2.115 $Y=0.18 $X2=0 $Y2=0
cc_674 N_SCE_M1040_g N_VGND_c_2250_n 0.00347568f $X=2.04 $Y=0.54 $X2=0 $Y2=0
cc_675 N_SCE_c_753_n N_VGND_c_2250_n 0.0261172f $X=3.995 $Y=0.18 $X2=0 $Y2=0
cc_676 N_SCE_c_753_n N_VGND_c_2251_n 0.00304147f $X=3.995 $Y=0.18 $X2=0 $Y2=0
cc_677 N_SCE_c_754_n N_VGND_c_2267_n 0.00203849f $X=2.115 $Y=0.18 $X2=0 $Y2=0
cc_678 N_SCE_c_753_n N_VGND_c_2268_n 0.00824997f $X=3.995 $Y=0.18 $X2=0 $Y2=0
cc_679 N_SCE_c_753_n N_VGND_c_2269_n 0.0360974f $X=3.995 $Y=0.18 $X2=0 $Y2=0
cc_680 N_SCE_c_753_n N_VGND_c_2275_n 0.0552579f $X=3.995 $Y=0.18 $X2=0 $Y2=0
cc_681 N_SCE_c_754_n N_VGND_c_2275_n 0.00419856f $X=2.115 $Y=0.18 $X2=0 $Y2=0
cc_682 N_SCD_c_857_n N_A_213_47#_c_904_n 0.0010218f $X=4.805 $Y=1.87 $X2=0 $Y2=0
cc_683 N_SCD_c_857_n N_A_213_47#_c_911_n 0.00826498f $X=4.805 $Y=1.87 $X2=0
+ $Y2=0
cc_684 SCD N_A_213_47#_c_911_n 0.00460548f $X=4.845 $Y=1.53 $X2=0 $Y2=0
cc_685 N_SCD_c_857_n N_VPWR_c_1872_n 0.0113733f $X=4.805 $Y=1.87 $X2=0 $Y2=0
cc_686 N_SCD_c_857_n N_VPWR_c_1882_n 0.00393283f $X=4.805 $Y=1.87 $X2=0 $Y2=0
cc_687 N_SCD_c_857_n N_VPWR_c_1869_n 0.00453105f $X=4.805 $Y=1.87 $X2=0 $Y2=0
cc_688 SCD N_A_700_389#_c_2078_n 4.80713e-19 $X=4.845 $Y=1.53 $X2=0 $Y2=0
cc_689 N_SCD_c_857_n N_A_700_389#_c_2086_n 0.0196372f $X=4.805 $Y=1.87 $X2=0
+ $Y2=0
cc_690 SCD N_A_700_389#_c_2086_n 0.0161525f $X=4.845 $Y=1.53 $X2=0 $Y2=0
cc_691 N_SCD_c_857_n N_A_700_389#_c_2079_n 0.00936494f $X=4.805 $Y=1.87 $X2=0
+ $Y2=0
cc_692 N_SCD_M1038_g N_A_700_389#_c_2079_n 0.0104512f $X=4.955 $Y=0.54 $X2=0
+ $Y2=0
cc_693 SCD N_A_700_389#_c_2079_n 0.0555582f $X=4.845 $Y=1.53 $X2=0 $Y2=0
cc_694 N_SCD_M1038_g N_A_700_389#_c_2081_n 0.00189328f $X=4.955 $Y=0.54 $X2=0
+ $Y2=0
cc_695 SCD N_A_700_389#_c_2081_n 0.0141018f $X=4.845 $Y=1.53 $X2=0 $Y2=0
cc_696 N_SCD_M1038_g N_A_700_389#_c_2082_n 0.00252094f $X=4.955 $Y=0.54 $X2=0
+ $Y2=0
cc_697 N_SCD_M1038_g N_VGND_c_2251_n 0.0114851f $X=4.955 $Y=0.54 $X2=0 $Y2=0
cc_698 N_SCD_M1038_g N_VGND_c_2269_n 0.003803f $X=4.955 $Y=0.54 $X2=0 $Y2=0
cc_699 SCD N_VGND_c_2269_n 0.00509611f $X=4.845 $Y=1.53 $X2=0 $Y2=0
cc_700 N_SCD_M1038_g N_VGND_c_2275_n 0.00593258f $X=4.955 $Y=0.54 $X2=0 $Y2=0
cc_701 SCD N_VGND_c_2275_n 0.00935171f $X=4.845 $Y=1.53 $X2=0 $Y2=0
cc_702 SCD A_899_66# 0.00441858f $X=4.845 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_703 N_A_213_47#_c_907_n N_A_1380_303#_M1009_d 4.47962e-19 $X=9.185 $Y=1.58
+ $X2=0 $Y2=0
cc_704 N_A_213_47#_c_1027_p N_A_1380_303#_M1009_d 0.00162221f $X=8.97 $Y=1.58
+ $X2=0 $Y2=0
cc_705 N_A_213_47#_c_913_n N_A_1380_303#_M1009_d 0.00213949f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_706 N_A_213_47#_c_913_n N_A_1380_303#_c_1149_n 0.00743564f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_707 N_A_213_47#_c_894_n N_A_1380_303#_M1000_g 0.0284532f $X=6.535 $Y=0.705
+ $X2=0 $Y2=0
cc_708 N_A_213_47#_c_897_n N_A_1380_303#_M1000_g 0.00103623f $X=6.425 $Y=0.87
+ $X2=0 $Y2=0
cc_709 N_A_213_47#_c_913_n N_A_1380_303#_c_1151_n 0.0215347f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_710 N_A_213_47#_c_895_n N_A_1380_303#_c_1175_n 0.00355011f $X=8.71 $Y=0.705
+ $X2=0 $Y2=0
cc_711 N_A_213_47#_c_907_n N_A_1380_303#_c_1160_n 9.4112e-19 $X=9.185 $Y=1.58
+ $X2=0 $Y2=0
cc_712 N_A_213_47#_c_1027_p N_A_1380_303#_c_1160_n 0.0153343f $X=8.97 $Y=1.58
+ $X2=0 $Y2=0
cc_713 N_A_213_47#_c_910_n N_A_1380_303#_c_1160_n 0.00698349f $X=9.315 $Y=1.58
+ $X2=0 $Y2=0
cc_714 N_A_213_47#_c_913_n N_A_1380_303#_c_1160_n 0.0191796f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_715 N_A_213_47#_c_916_n N_A_1380_303#_c_1160_n 0.00118114f $X=9.65 $Y=1.87
+ $X2=0 $Y2=0
cc_716 N_A_213_47#_c_898_n N_A_1380_303#_c_1164_n 0.0577028f $X=8.835 $Y=0.87
+ $X2=0 $Y2=0
cc_717 N_A_213_47#_c_899_n N_A_1380_303#_c_1164_n 0.00355011f $X=8.835 $Y=0.87
+ $X2=0 $Y2=0
cc_718 N_A_213_47#_c_910_n N_A_1380_303#_c_1152_n 0.00193134f $X=9.315 $Y=1.58
+ $X2=0 $Y2=0
cc_719 N_A_213_47#_c_913_n N_A_1380_303#_c_1152_n 0.0225494f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_720 N_A_213_47#_c_1027_p N_A_1380_303#_c_1148_n 0.0126476f $X=8.97 $Y=1.58
+ $X2=0 $Y2=0
cc_721 N_A_213_47#_c_913_n N_RESET_B_c_1255_n 0.00403964f $X=9.5 $Y=1.87 $X2=0
+ $Y2=0
cc_722 N_A_213_47#_c_913_n N_RESET_B_c_1269_n 0.00114418f $X=9.5 $Y=1.87 $X2=0
+ $Y2=0
cc_723 N_A_213_47#_c_898_n N_RESET_B_c_1260_n 0.017273f $X=8.835 $Y=0.87 $X2=0
+ $Y2=0
cc_724 N_A_213_47#_c_899_n N_RESET_B_c_1260_n 0.00333579f $X=8.835 $Y=0.87 $X2=0
+ $Y2=0
cc_725 N_A_213_47#_c_895_n N_A_1202_413#_M1041_g 0.0112202f $X=8.71 $Y=0.705
+ $X2=0 $Y2=0
cc_726 N_A_213_47#_c_898_n N_A_1202_413#_M1041_g 2.98198e-19 $X=8.835 $Y=0.87
+ $X2=0 $Y2=0
cc_727 N_A_213_47#_c_898_n N_A_1202_413#_c_1429_n 0.00284065f $X=8.835 $Y=0.87
+ $X2=0 $Y2=0
cc_728 N_A_213_47#_c_899_n N_A_1202_413#_c_1429_n 0.00446614f $X=8.835 $Y=0.87
+ $X2=0 $Y2=0
cc_729 N_A_213_47#_c_1027_p N_A_1202_413#_c_1429_n 0.00258112f $X=8.97 $Y=1.58
+ $X2=0 $Y2=0
cc_730 N_A_213_47#_c_1027_p N_A_1202_413#_c_1430_n 0.00299851f $X=8.97 $Y=1.58
+ $X2=0 $Y2=0
cc_731 N_A_213_47#_c_910_n N_A_1202_413#_c_1430_n 7.63882e-19 $X=9.315 $Y=1.58
+ $X2=0 $Y2=0
cc_732 N_A_213_47#_c_913_n N_A_1202_413#_c_1430_n 0.00286067f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_733 N_A_213_47#_c_894_n N_A_1202_413#_c_1462_n 0.00884831f $X=6.535 $Y=0.705
+ $X2=0 $Y2=0
cc_734 N_A_213_47#_c_896_n N_A_1202_413#_c_1462_n 4.06924e-19 $X=6.12 $Y=0.87
+ $X2=0 $Y2=0
cc_735 N_A_213_47#_c_897_n N_A_1202_413#_c_1462_n 0.026125f $X=6.425 $Y=0.87
+ $X2=0 $Y2=0
cc_736 N_A_213_47#_c_902_n N_A_1202_413#_c_1462_n 0.00351458f $X=6.535 $Y=0.87
+ $X2=0 $Y2=0
cc_737 N_A_213_47#_c_897_n N_A_1202_413#_c_1423_n 0.0116356f $X=6.425 $Y=0.87
+ $X2=0 $Y2=0
cc_738 N_A_213_47#_c_913_n N_A_1202_413#_c_1423_n 0.00602557f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_739 N_A_213_47#_c_902_n N_A_1202_413#_c_1423_n 8.05093e-19 $X=6.535 $Y=0.87
+ $X2=0 $Y2=0
cc_740 N_A_213_47#_c_897_n N_A_1202_413#_c_1424_n 0.0106449f $X=6.425 $Y=0.87
+ $X2=0 $Y2=0
cc_741 N_A_213_47#_c_902_n N_A_1202_413#_c_1424_n 8.73594e-19 $X=6.535 $Y=0.87
+ $X2=0 $Y2=0
cc_742 N_A_213_47#_c_903_n N_A_1202_413#_c_1424_n 0.0127672f $X=5.97 $Y=1.575
+ $X2=0 $Y2=0
cc_743 N_A_213_47#_c_894_n N_A_1202_413#_c_1425_n 0.0046359f $X=6.535 $Y=0.705
+ $X2=0 $Y2=0
cc_744 N_A_213_47#_c_897_n N_A_1202_413#_c_1425_n 0.0246688f $X=6.425 $Y=0.87
+ $X2=0 $Y2=0
cc_745 N_A_213_47#_c_902_n N_A_1202_413#_c_1425_n 0.00103235f $X=6.535 $Y=0.87
+ $X2=0 $Y2=0
cc_746 N_A_213_47#_c_904_n N_A_1202_413#_c_1447_n 0.00422393f $X=5.92 $Y=1.99
+ $X2=0 $Y2=0
cc_747 N_A_213_47#_c_913_n N_A_1202_413#_c_1447_n 0.00363572f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_748 N_A_213_47#_c_914_n N_A_1202_413#_c_1447_n 0.00241651f $X=6.18 $Y=1.87
+ $X2=0 $Y2=0
cc_749 N_A_213_47#_c_917_n N_A_1202_413#_c_1447_n 0.00151282f $X=5.905 $Y=1.74
+ $X2=0 $Y2=0
cc_750 N_A_213_47#_c_904_n N_A_1202_413#_c_1433_n 0.00353099f $X=5.92 $Y=1.99
+ $X2=0 $Y2=0
cc_751 N_A_213_47#_c_913_n N_A_1202_413#_c_1433_n 0.0170664f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_752 N_A_213_47#_c_914_n N_A_1202_413#_c_1433_n 0.00296099f $X=6.18 $Y=1.87
+ $X2=0 $Y2=0
cc_753 N_A_213_47#_c_903_n N_A_1202_413#_c_1433_n 0.0415032f $X=5.97 $Y=1.575
+ $X2=0 $Y2=0
cc_754 N_A_213_47#_c_913_n N_A_1202_413#_c_1434_n 0.00155738f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_755 N_A_213_47#_c_899_n N_A_1202_413#_c_1428_n 0.0112202f $X=8.835 $Y=0.87
+ $X2=0 $Y2=0
cc_756 N_A_213_47#_c_913_n N_A_1202_413#_c_1428_n 4.37453e-19 $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_757 N_A_213_47#_c_905_n N_A_1972_21#_c_1562_n 0.0164563f $X=9.665 $Y=1.99
+ $X2=0 $Y2=0
cc_758 N_A_213_47#_c_910_n N_A_1972_21#_c_1562_n 4.60638e-19 $X=9.315 $Y=1.58
+ $X2=0 $Y2=0
cc_759 N_A_213_47#_c_918_n N_A_1972_21#_c_1562_n 0.0010053f $X=9.63 $Y=1.745
+ $X2=0 $Y2=0
cc_760 N_A_213_47#_c_905_n N_A_1972_21#_c_1580_n 0.0262728f $X=9.665 $Y=1.99
+ $X2=0 $Y2=0
cc_761 N_A_213_47#_c_895_n N_A_1757_47#_c_1764_n 0.00279863f $X=8.71 $Y=0.705
+ $X2=0 $Y2=0
cc_762 N_A_213_47#_c_898_n N_A_1757_47#_c_1764_n 0.0116575f $X=8.835 $Y=0.87
+ $X2=0 $Y2=0
cc_763 N_A_213_47#_c_899_n N_A_1757_47#_c_1764_n 0.00120647f $X=8.835 $Y=0.87
+ $X2=0 $Y2=0
cc_764 N_A_213_47#_c_905_n N_A_1757_47#_c_1767_n 0.0149309f $X=9.665 $Y=1.99
+ $X2=0 $Y2=0
cc_765 N_A_213_47#_c_910_n N_A_1757_47#_c_1767_n 0.0160793f $X=9.315 $Y=1.58
+ $X2=0 $Y2=0
cc_766 N_A_213_47#_c_913_n N_A_1757_47#_c_1767_n 0.00142849f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_767 N_A_213_47#_c_916_n N_A_1757_47#_c_1767_n 0.00316956f $X=9.65 $Y=1.87
+ $X2=0 $Y2=0
cc_768 N_A_213_47#_c_918_n N_A_1757_47#_c_1767_n 0.0230959f $X=9.63 $Y=1.745
+ $X2=0 $Y2=0
cc_769 N_A_213_47#_c_905_n N_A_1757_47#_c_1761_n 0.00282444f $X=9.665 $Y=1.99
+ $X2=0 $Y2=0
cc_770 N_A_213_47#_c_916_n N_A_1757_47#_c_1761_n 0.00266839f $X=9.65 $Y=1.87
+ $X2=0 $Y2=0
cc_771 N_A_213_47#_c_918_n N_A_1757_47#_c_1761_n 0.013964f $X=9.63 $Y=1.745
+ $X2=0 $Y2=0
cc_772 N_A_213_47#_c_905_n N_A_1757_47#_c_1762_n 0.00534461f $X=9.665 $Y=1.99
+ $X2=0 $Y2=0
cc_773 N_A_213_47#_c_910_n N_A_1757_47#_c_1762_n 0.00576712f $X=9.315 $Y=1.58
+ $X2=0 $Y2=0
cc_774 N_A_213_47#_c_916_n N_A_1757_47#_c_1762_n 8.39805e-19 $X=9.65 $Y=1.87
+ $X2=0 $Y2=0
cc_775 N_A_213_47#_c_918_n N_A_1757_47#_c_1762_n 0.0203823f $X=9.63 $Y=1.745
+ $X2=0 $Y2=0
cc_776 N_A_213_47#_c_913_n N_VPWR_M1009_s 3.30587e-19 $X=9.5 $Y=1.87 $X2=0 $Y2=0
cc_777 N_A_213_47#_c_915_n N_VPWR_c_1870_n 0.0203051f $X=1.22 $Y=1.87 $X2=0
+ $Y2=0
cc_778 N_A_213_47#_c_911_n N_VPWR_c_1871_n 0.00655717f $X=5.89 $Y=1.87 $X2=0
+ $Y2=0
cc_779 N_A_213_47#_c_904_n N_VPWR_c_1872_n 0.00247711f $X=5.92 $Y=1.99 $X2=0
+ $Y2=0
cc_780 N_A_213_47#_c_911_n N_VPWR_c_1872_n 0.00124277f $X=5.89 $Y=1.87 $X2=0
+ $Y2=0
cc_781 N_A_213_47#_c_913_n N_VPWR_c_1873_n 0.00271934f $X=9.5 $Y=1.87 $X2=0
+ $Y2=0
cc_782 N_A_213_47#_c_915_n N_VPWR_c_1880_n 0.0160592f $X=1.22 $Y=1.87 $X2=0
+ $Y2=0
cc_783 N_A_213_47#_c_913_n N_VPWR_c_1884_n 0.00131844f $X=9.5 $Y=1.87 $X2=0
+ $Y2=0
cc_784 N_A_213_47#_c_904_n N_VPWR_c_1885_n 0.00691661f $X=5.92 $Y=1.99 $X2=0
+ $Y2=0
cc_785 N_A_213_47#_c_905_n N_VPWR_c_1886_n 0.00429453f $X=9.665 $Y=1.99 $X2=0
+ $Y2=0
cc_786 N_A_213_47#_M1033_d N_VPWR_c_1869_n 0.00224123f $X=1.07 $Y=1.485 $X2=0
+ $Y2=0
cc_787 N_A_213_47#_c_904_n N_VPWR_c_1869_n 0.0083956f $X=5.92 $Y=1.99 $X2=0
+ $Y2=0
cc_788 N_A_213_47#_c_905_n N_VPWR_c_1869_n 0.00611502f $X=9.665 $Y=1.99 $X2=0
+ $Y2=0
cc_789 N_A_213_47#_c_910_n N_VPWR_c_1869_n 6.28369e-19 $X=9.315 $Y=1.58 $X2=0
+ $Y2=0
cc_790 N_A_213_47#_c_911_n N_VPWR_c_1869_n 0.213784f $X=5.89 $Y=1.87 $X2=0 $Y2=0
cc_791 N_A_213_47#_c_912_n N_VPWR_c_1869_n 0.0154857f $X=1.37 $Y=1.87 $X2=0
+ $Y2=0
cc_792 N_A_213_47#_c_913_n N_VPWR_c_1869_n 0.1524f $X=9.5 $Y=1.87 $X2=0 $Y2=0
cc_793 N_A_213_47#_c_914_n N_VPWR_c_1869_n 0.0160418f $X=6.18 $Y=1.87 $X2=0
+ $Y2=0
cc_794 N_A_213_47#_c_915_n N_VPWR_c_1869_n 0.0039866f $X=1.22 $Y=1.87 $X2=0
+ $Y2=0
cc_795 N_A_213_47#_c_916_n N_VPWR_c_1869_n 0.0158166f $X=9.65 $Y=1.87 $X2=0
+ $Y2=0
cc_796 N_A_213_47#_c_917_n N_VPWR_c_1869_n 0.00320789f $X=5.905 $Y=1.74 $X2=0
+ $Y2=0
cc_797 N_A_213_47#_c_911_n N_A_700_389#_c_2078_n 0.013705f $X=5.89 $Y=1.87 $X2=0
+ $Y2=0
cc_798 N_A_213_47#_c_911_n N_A_700_389#_c_2086_n 0.0401661f $X=5.89 $Y=1.87
+ $X2=0 $Y2=0
cc_799 N_A_213_47#_c_904_n N_A_700_389#_c_2079_n 0.01374f $X=5.92 $Y=1.99 $X2=0
+ $Y2=0
cc_800 N_A_213_47#_c_896_n N_A_700_389#_c_2079_n 0.00490452f $X=6.12 $Y=0.87
+ $X2=0 $Y2=0
cc_801 N_A_213_47#_c_911_n N_A_700_389#_c_2079_n 0.0386379f $X=5.89 $Y=1.87
+ $X2=0 $Y2=0
cc_802 N_A_213_47#_c_914_n N_A_700_389#_c_2079_n 0.00129231f $X=6.18 $Y=1.87
+ $X2=0 $Y2=0
cc_803 N_A_213_47#_c_917_n N_A_700_389#_c_2079_n 0.0123086f $X=5.905 $Y=1.74
+ $X2=0 $Y2=0
cc_804 N_A_213_47#_c_903_n N_A_700_389#_c_2079_n 0.00675181f $X=5.97 $Y=1.575
+ $X2=0 $Y2=0
cc_805 N_A_213_47#_c_896_n N_A_700_389#_c_2080_n 0.0146758f $X=6.12 $Y=0.87
+ $X2=0 $Y2=0
cc_806 N_A_213_47#_c_902_n N_A_700_389#_c_2080_n 2.12824e-19 $X=6.535 $Y=0.87
+ $X2=0 $Y2=0
cc_807 N_A_213_47#_c_896_n N_A_700_389#_c_2082_n 6.94909e-19 $X=6.12 $Y=0.87
+ $X2=0 $Y2=0
cc_808 N_A_213_47#_c_911_n N_A_700_389#_c_2123_n 0.00501633f $X=5.89 $Y=1.87
+ $X2=0 $Y2=0
cc_809 N_A_213_47#_c_913_n N_A_1324_413#_c_2177_n 0.0251636f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_810 N_A_213_47#_c_913_n N_A_1324_413#_c_2178_n 0.00701432f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_811 N_A_213_47#_c_913_n N_A_1324_413#_c_2179_n 0.00567047f $X=9.5 $Y=1.87
+ $X2=0 $Y2=0
cc_812 N_A_213_47#_c_900_n N_VGND_c_2249_n 0.00137385f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_813 N_A_213_47#_c_894_n N_VGND_c_2258_n 0.00368123f $X=6.535 $Y=0.705 $X2=0
+ $Y2=0
cc_814 N_A_213_47#_c_896_n N_VGND_c_2258_n 0.00333937f $X=6.12 $Y=0.87 $X2=0
+ $Y2=0
cc_815 N_A_213_47#_c_895_n N_VGND_c_2260_n 0.0050861f $X=8.71 $Y=0.705 $X2=0
+ $Y2=0
cc_816 N_A_213_47#_c_898_n N_VGND_c_2260_n 0.00106209f $X=8.835 $Y=0.87 $X2=0
+ $Y2=0
cc_817 N_A_213_47#_c_900_n N_VGND_c_2267_n 0.0107699f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_818 N_A_213_47#_M1002_d N_VGND_c_2275_n 0.00394021f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_819 N_A_213_47#_c_894_n N_VGND_c_2275_n 0.00584426f $X=6.535 $Y=0.705 $X2=0
+ $Y2=0
cc_820 N_A_213_47#_c_895_n N_VGND_c_2275_n 0.00639584f $X=8.71 $Y=0.705 $X2=0
+ $Y2=0
cc_821 N_A_213_47#_c_896_n N_VGND_c_2275_n 0.00520195f $X=6.12 $Y=0.87 $X2=0
+ $Y2=0
cc_822 N_A_213_47#_c_898_n N_VGND_c_2275_n 0.00110317f $X=8.835 $Y=0.87 $X2=0
+ $Y2=0
cc_823 N_A_213_47#_c_900_n N_VGND_c_2275_n 0.00903594f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_824 N_A_1380_303#_c_1149_n N_RESET_B_c_1255_n 0.0272425f $X=7 $Y=1.99 $X2=0
+ $Y2=0
cc_825 N_A_1380_303#_M1000_g N_RESET_B_c_1255_n 0.0133987f $X=7.065 $Y=0.445
+ $X2=0 $Y2=0
cc_826 N_A_1380_303#_c_1151_n N_RESET_B_c_1255_n 0.0140624f $X=8.23 $Y=1.68
+ $X2=0 $Y2=0
cc_827 N_A_1380_303#_c_1152_n N_RESET_B_c_1255_n 0.00346452f $X=8.385 $Y=1.68
+ $X2=0 $Y2=0
cc_828 N_A_1380_303#_c_1148_n N_RESET_B_c_1255_n 4.85413e-19 $X=8.385 $Y=1.595
+ $X2=0 $Y2=0
cc_829 N_A_1380_303#_c_1149_n N_RESET_B_c_1269_n 0.0155095f $X=7 $Y=1.99 $X2=0
+ $Y2=0
cc_830 N_A_1380_303#_M1000_g N_RESET_B_c_1258_n 0.00499546f $X=7.065 $Y=0.445
+ $X2=0 $Y2=0
cc_831 N_A_1380_303#_M1000_g N_RESET_B_c_1259_n 0.00200402f $X=7.065 $Y=0.445
+ $X2=0 $Y2=0
cc_832 N_A_1380_303#_c_1164_n N_RESET_B_c_1259_n 0.00174508f $X=8.385 $Y=0.835
+ $X2=0 $Y2=0
cc_833 N_A_1380_303#_c_1148_n N_RESET_B_c_1259_n 0.00296076f $X=8.385 $Y=1.595
+ $X2=0 $Y2=0
cc_834 N_A_1380_303#_c_1196_p N_RESET_B_c_1260_n 0.00176185f $X=8.445 $Y=0.36
+ $X2=0 $Y2=0
cc_835 N_A_1380_303#_c_1164_n N_RESET_B_c_1260_n 0.0145363f $X=8.385 $Y=0.835
+ $X2=0 $Y2=0
cc_836 N_A_1380_303#_c_1148_n N_RESET_B_c_1260_n 0.00587291f $X=8.385 $Y=1.595
+ $X2=0 $Y2=0
cc_837 N_A_1380_303#_c_1164_n N_RESET_B_c_1261_n 0.00178696f $X=8.385 $Y=0.835
+ $X2=0 $Y2=0
cc_838 N_A_1380_303#_c_1148_n N_RESET_B_c_1261_n 0.00124848f $X=8.385 $Y=1.595
+ $X2=0 $Y2=0
cc_839 N_A_1380_303#_M1000_g N_RESET_B_c_1265_n 0.0491516f $X=7.065 $Y=0.445
+ $X2=0 $Y2=0
cc_840 N_A_1380_303#_c_1196_p N_RESET_B_c_1265_n 9.53262e-19 $X=8.445 $Y=0.36
+ $X2=0 $Y2=0
cc_841 N_A_1380_303#_c_1175_n N_A_1202_413#_M1041_g 0.00639817f $X=8.385 $Y=0.68
+ $X2=0 $Y2=0
cc_842 N_A_1380_303#_c_1196_p N_A_1202_413#_M1041_g 0.00331537f $X=8.445 $Y=0.36
+ $X2=0 $Y2=0
cc_843 N_A_1380_303#_c_1164_n N_A_1202_413#_M1041_g 0.00652415f $X=8.385
+ $Y=0.835 $X2=0 $Y2=0
cc_844 N_A_1380_303#_c_1148_n N_A_1202_413#_M1041_g 0.0115826f $X=8.385 $Y=1.595
+ $X2=0 $Y2=0
cc_845 N_A_1380_303#_c_1160_n N_A_1202_413#_c_1429_n 6.65821e-19 $X=8.815
+ $Y=1.92 $X2=0 $Y2=0
cc_846 N_A_1380_303#_c_1164_n N_A_1202_413#_c_1429_n 8.88512e-19 $X=8.385
+ $Y=0.835 $X2=0 $Y2=0
cc_847 N_A_1380_303#_c_1148_n N_A_1202_413#_c_1429_n 0.0144528f $X=8.385
+ $Y=1.595 $X2=0 $Y2=0
cc_848 N_A_1380_303#_c_1160_n N_A_1202_413#_c_1430_n 0.0149935f $X=8.815 $Y=1.92
+ $X2=0 $Y2=0
cc_849 N_A_1380_303#_c_1163_n N_A_1202_413#_c_1430_n 0.00489841f $X=8.9 $Y=2.3
+ $X2=0 $Y2=0
cc_850 N_A_1380_303#_c_1152_n N_A_1202_413#_c_1430_n 0.00197846f $X=8.385
+ $Y=1.68 $X2=0 $Y2=0
cc_851 N_A_1380_303#_c_1148_n N_A_1202_413#_c_1430_n 0.00574694f $X=8.385
+ $Y=1.595 $X2=0 $Y2=0
cc_852 N_A_1380_303#_M1000_g N_A_1202_413#_c_1462_n 0.005989f $X=7.065 $Y=0.445
+ $X2=0 $Y2=0
cc_853 N_A_1380_303#_M1000_g N_A_1202_413#_c_1425_n 0.0190937f $X=7.065 $Y=0.445
+ $X2=0 $Y2=0
cc_854 N_A_1380_303#_c_1149_n N_A_1202_413#_c_1426_n 0.00410583f $X=7 $Y=1.99
+ $X2=0 $Y2=0
cc_855 N_A_1380_303#_M1000_g N_A_1202_413#_c_1426_n 0.00957327f $X=7.065
+ $Y=0.445 $X2=0 $Y2=0
cc_856 N_A_1380_303#_c_1151_n N_A_1202_413#_c_1426_n 0.0498518f $X=8.23 $Y=1.68
+ $X2=0 $Y2=0
cc_857 N_A_1380_303#_c_1149_n N_A_1202_413#_c_1433_n 0.00235419f $X=7 $Y=1.99
+ $X2=0 $Y2=0
cc_858 N_A_1380_303#_M1000_g N_A_1202_413#_c_1433_n 5.64424e-19 $X=7.065
+ $Y=0.445 $X2=0 $Y2=0
cc_859 N_A_1380_303#_c_1151_n N_A_1202_413#_c_1433_n 0.00529221f $X=8.23 $Y=1.68
+ $X2=0 $Y2=0
cc_860 N_A_1380_303#_c_1149_n N_A_1202_413#_c_1434_n 0.00292203f $X=7 $Y=1.99
+ $X2=0 $Y2=0
cc_861 N_A_1380_303#_M1000_g N_A_1202_413#_c_1434_n 0.00334413f $X=7.065
+ $Y=0.445 $X2=0 $Y2=0
cc_862 N_A_1380_303#_c_1151_n N_A_1202_413#_c_1434_n 0.00280794f $X=8.23 $Y=1.68
+ $X2=0 $Y2=0
cc_863 N_A_1380_303#_c_1151_n N_A_1202_413#_c_1427_n 0.0096056f $X=8.23 $Y=1.68
+ $X2=0 $Y2=0
cc_864 N_A_1380_303#_c_1148_n N_A_1202_413#_c_1427_n 0.0213978f $X=8.385
+ $Y=1.595 $X2=0 $Y2=0
cc_865 N_A_1380_303#_c_1151_n N_A_1202_413#_c_1428_n 0.00617564f $X=8.23 $Y=1.68
+ $X2=0 $Y2=0
cc_866 N_A_1380_303#_c_1152_n N_A_1202_413#_c_1428_n 0.00687455f $X=8.385
+ $Y=1.68 $X2=0 $Y2=0
cc_867 N_A_1380_303#_c_1175_n N_A_1757_47#_c_1764_n 0.00556097f $X=8.385 $Y=0.68
+ $X2=0 $Y2=0
cc_868 N_A_1380_303#_c_1163_n N_A_1757_47#_c_1767_n 0.0225461f $X=8.9 $Y=2.3
+ $X2=0 $Y2=0
cc_869 N_A_1380_303#_c_1152_n N_VPWR_M1009_s 0.00479206f $X=8.385 $Y=1.68 $X2=0
+ $Y2=0
cc_870 N_A_1380_303#_c_1151_n N_VPWR_c_1873_n 0.00180429f $X=8.23 $Y=1.68 $X2=0
+ $Y2=0
cc_871 N_A_1380_303#_c_1163_n N_VPWR_c_1873_n 0.017731f $X=8.9 $Y=2.3 $X2=0
+ $Y2=0
cc_872 N_A_1380_303#_c_1152_n N_VPWR_c_1873_n 0.0219424f $X=8.385 $Y=1.68 $X2=0
+ $Y2=0
cc_873 N_A_1380_303#_c_1149_n N_VPWR_c_1884_n 0.00401376f $X=7 $Y=1.99 $X2=0
+ $Y2=0
cc_874 N_A_1380_303#_c_1149_n N_VPWR_c_1885_n 0.00513013f $X=7 $Y=1.99 $X2=0
+ $Y2=0
cc_875 N_A_1380_303#_c_1160_n N_VPWR_c_1886_n 0.00301931f $X=8.815 $Y=1.92 $X2=0
+ $Y2=0
cc_876 N_A_1380_303#_c_1163_n N_VPWR_c_1886_n 0.0117479f $X=8.9 $Y=2.3 $X2=0
+ $Y2=0
cc_877 N_A_1380_303#_M1009_d N_VPWR_c_1869_n 0.00327123f $X=8.75 $Y=1.645 $X2=0
+ $Y2=0
cc_878 N_A_1380_303#_c_1149_n N_VPWR_c_1869_n 0.0067254f $X=7 $Y=1.99 $X2=0
+ $Y2=0
cc_879 N_A_1380_303#_c_1160_n N_VPWR_c_1869_n 0.00245611f $X=8.815 $Y=1.92 $X2=0
+ $Y2=0
cc_880 N_A_1380_303#_c_1163_n N_VPWR_c_1869_n 0.00306902f $X=8.9 $Y=2.3 $X2=0
+ $Y2=0
cc_881 N_A_1380_303#_c_1152_n N_VPWR_c_1869_n 8.41228e-19 $X=8.385 $Y=1.68 $X2=0
+ $Y2=0
cc_882 N_A_1380_303#_c_1149_n N_A_1324_413#_c_2177_n 0.0168268f $X=7 $Y=1.99
+ $X2=0 $Y2=0
cc_883 N_A_1380_303#_c_1151_n N_A_1324_413#_c_2177_n 0.0496655f $X=8.23 $Y=1.68
+ $X2=0 $Y2=0
cc_884 N_A_1380_303#_c_1149_n N_A_1324_413#_c_2178_n 2.52506e-19 $X=7 $Y=1.99
+ $X2=0 $Y2=0
cc_885 N_A_1380_303#_c_1151_n N_A_1324_413#_c_2179_n 0.011083f $X=8.23 $Y=1.68
+ $X2=0 $Y2=0
cc_886 N_A_1380_303#_c_1152_n N_A_1324_413#_c_2179_n 0.00375057f $X=8.385
+ $Y=1.68 $X2=0 $Y2=0
cc_887 N_A_1380_303#_c_1196_p N_VGND_c_2252_n 0.0178713f $X=8.445 $Y=0.36 $X2=0
+ $Y2=0
cc_888 N_A_1380_303#_M1000_g N_VGND_c_2258_n 0.0055639f $X=7.065 $Y=0.445 $X2=0
+ $Y2=0
cc_889 N_A_1380_303#_c_1196_p N_VGND_c_2260_n 0.0203886f $X=8.445 $Y=0.36 $X2=0
+ $Y2=0
cc_890 N_A_1380_303#_M1041_d N_VGND_c_2275_n 0.00233415f $X=8.31 $Y=0.235 $X2=0
+ $Y2=0
cc_891 N_A_1380_303#_M1000_g N_VGND_c_2275_n 0.0103614f $X=7.065 $Y=0.445 $X2=0
+ $Y2=0
cc_892 N_A_1380_303#_c_1196_p N_VGND_c_2275_n 0.00654291f $X=8.445 $Y=0.36 $X2=0
+ $Y2=0
cc_893 N_RESET_B_c_1259_n N_A_1202_413#_M1041_g 0.00200706f $X=7.7 $Y=0.85 $X2=0
+ $Y2=0
cc_894 N_RESET_B_c_1260_n N_A_1202_413#_M1041_g 0.00452207f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_895 N_RESET_B_c_1261_n N_A_1202_413#_M1041_g 0.00174935f $X=7.9 $Y=0.85 $X2=0
+ $Y2=0
cc_896 N_RESET_B_c_1264_n N_A_1202_413#_M1041_g 0.0062745f $X=7.535 $Y=0.96
+ $X2=0 $Y2=0
cc_897 N_RESET_B_c_1265_n N_A_1202_413#_M1041_g 0.00995576f $X=7.56 $Y=0.755
+ $X2=0 $Y2=0
cc_898 N_RESET_B_c_1265_n N_A_1202_413#_c_1462_n 8.20253e-19 $X=7.56 $Y=0.755
+ $X2=0 $Y2=0
cc_899 N_RESET_B_c_1255_n N_A_1202_413#_c_1425_n 5.71854e-19 $X=7.62 $Y=1.89
+ $X2=0 $Y2=0
cc_900 N_RESET_B_c_1258_n N_A_1202_413#_c_1425_n 0.00850069f $X=7.785 $Y=0.85
+ $X2=0 $Y2=0
cc_901 N_RESET_B_c_1259_n N_A_1202_413#_c_1425_n 0.0148433f $X=7.7 $Y=0.85 $X2=0
+ $Y2=0
cc_902 N_RESET_B_c_1264_n N_A_1202_413#_c_1425_n 6.64193e-19 $X=7.535 $Y=0.96
+ $X2=0 $Y2=0
cc_903 N_RESET_B_c_1265_n N_A_1202_413#_c_1425_n 0.00140348f $X=7.56 $Y=0.755
+ $X2=0 $Y2=0
cc_904 N_RESET_B_c_1255_n N_A_1202_413#_c_1426_n 0.0118406f $X=7.62 $Y=1.89
+ $X2=0 $Y2=0
cc_905 N_RESET_B_c_1258_n N_A_1202_413#_c_1426_n 0.00117441f $X=7.785 $Y=0.85
+ $X2=0 $Y2=0
cc_906 N_RESET_B_c_1259_n N_A_1202_413#_c_1426_n 0.0374317f $X=7.7 $Y=0.85 $X2=0
+ $Y2=0
cc_907 N_RESET_B_c_1260_n N_A_1202_413#_c_1426_n 4.29892e-19 $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_908 N_RESET_B_c_1261_n N_A_1202_413#_c_1426_n 3.52736e-19 $X=7.9 $Y=0.85
+ $X2=0 $Y2=0
cc_909 N_RESET_B_c_1264_n N_A_1202_413#_c_1426_n 0.00251038f $X=7.535 $Y=0.96
+ $X2=0 $Y2=0
cc_910 N_RESET_B_c_1259_n N_A_1202_413#_c_1427_n 0.00316807f $X=7.7 $Y=0.85
+ $X2=0 $Y2=0
cc_911 N_RESET_B_c_1260_n N_A_1202_413#_c_1427_n 0.00429153f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_912 N_RESET_B_c_1264_n N_A_1202_413#_c_1427_n 0.00141794f $X=7.535 $Y=0.96
+ $X2=0 $Y2=0
cc_913 N_RESET_B_c_1255_n N_A_1202_413#_c_1428_n 0.00859083f $X=7.62 $Y=1.89
+ $X2=0 $Y2=0
cc_914 N_RESET_B_c_1259_n N_A_1202_413#_c_1428_n 2.69296e-19 $X=7.7 $Y=0.85
+ $X2=0 $Y2=0
cc_915 N_RESET_B_c_1260_n N_A_1202_413#_c_1428_n 0.00102675f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_916 N_RESET_B_c_1264_n N_A_1202_413#_c_1428_n 0.0221169f $X=7.535 $Y=0.96
+ $X2=0 $Y2=0
cc_917 N_RESET_B_c_1267_n N_A_1972_21#_M1012_d 7.28066e-19 $X=11.26 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_918 N_RESET_B_M1006_g N_A_1972_21#_M1032_g 0.00764787f $X=10.71 $Y=0.445
+ $X2=0 $Y2=0
cc_919 N_RESET_B_c_1260_n N_A_1972_21#_M1032_g 0.00240753f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_920 N_RESET_B_c_1257_n N_A_1972_21#_c_1562_n 0.00307301f $X=11.065 $Y=1.17
+ $X2=0 $Y2=0
cc_921 N_RESET_B_c_1266_n N_A_1972_21#_c_1562_n 0.0138081f $X=10.77 $Y=1.15
+ $X2=0 $Y2=0
cc_922 N_RESET_B_c_1270_n N_A_1972_21#_c_1580_n 0.0138081f $X=10.735 $Y=1.89
+ $X2=0 $Y2=0
cc_923 N_RESET_B_c_1271_n N_A_1972_21#_c_1580_n 0.0132989f $X=10.735 $Y=1.99
+ $X2=0 $Y2=0
cc_924 N_RESET_B_M1006_g N_A_1972_21#_c_1570_n 0.00140538f $X=10.71 $Y=0.445
+ $X2=0 $Y2=0
cc_925 N_RESET_B_c_1257_n N_A_1972_21#_c_1570_n 0.00478211f $X=11.065 $Y=1.17
+ $X2=0 $Y2=0
cc_926 N_RESET_B_c_1260_n N_A_1972_21#_c_1570_n 0.00933039f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_927 N_RESET_B_c_1262_n N_A_1972_21#_c_1570_n 3.71404e-19 $X=10.92 $Y=1.17
+ $X2=0 $Y2=0
cc_928 RESET_B N_A_1972_21#_c_1570_n 0.00483613f $X=11.185 $Y=0.765 $X2=0 $Y2=0
cc_929 N_RESET_B_M1006_g N_A_1972_21#_c_1571_n 0.00629891f $X=10.71 $Y=0.445
+ $X2=0 $Y2=0
cc_930 N_RESET_B_c_1257_n N_A_1972_21#_c_1571_n 0.00682325f $X=11.065 $Y=1.17
+ $X2=0 $Y2=0
cc_931 N_RESET_B_c_1260_n N_A_1972_21#_c_1571_n 0.0179653f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_932 RESET_B N_A_1972_21#_c_1571_n 2.94839e-19 $X=11.185 $Y=0.765 $X2=0 $Y2=0
cc_933 N_RESET_B_c_1267_n N_A_1972_21#_c_1571_n 0.00669372f $X=11.26 $Y=0.85
+ $X2=0 $Y2=0
cc_934 N_RESET_B_c_1260_n N_A_1972_21#_c_1572_n 0.00679872f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_935 N_RESET_B_M1006_g N_A_1972_21#_c_1573_n 0.00756196f $X=10.71 $Y=0.445
+ $X2=0 $Y2=0
cc_936 N_RESET_B_c_1267_n N_A_1972_21#_c_1573_n 0.00216331f $X=11.26 $Y=0.85
+ $X2=0 $Y2=0
cc_937 N_RESET_B_M1006_g N_A_1972_21#_c_1574_n 0.00502769f $X=10.71 $Y=0.445
+ $X2=0 $Y2=0
cc_938 N_RESET_B_c_1257_n N_A_1972_21#_c_1574_n 0.00379117f $X=11.065 $Y=1.17
+ $X2=0 $Y2=0
cc_939 N_RESET_B_c_1260_n N_A_1972_21#_c_1574_n 0.00469044f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_940 RESET_B N_A_1972_21#_c_1574_n 0.00195155f $X=11.185 $Y=0.765 $X2=0 $Y2=0
cc_941 N_RESET_B_c_1266_n N_A_1972_21#_c_1574_n 0.00163075f $X=10.77 $Y=1.15
+ $X2=0 $Y2=0
cc_942 N_RESET_B_c_1267_n N_A_1972_21#_c_1574_n 0.0132934f $X=11.26 $Y=0.85
+ $X2=0 $Y2=0
cc_943 N_RESET_B_M1006_g N_A_1972_21#_c_1626_n 0.00441127f $X=10.71 $Y=0.445
+ $X2=0 $Y2=0
cc_944 N_RESET_B_c_1271_n N_A_1972_21#_c_1589_n 0.00522156f $X=10.735 $Y=1.99
+ $X2=0 $Y2=0
cc_945 RESET_B N_A_1972_21#_c_1575_n 0.00762142f $X=11.185 $Y=0.765 $X2=0 $Y2=0
cc_946 N_RESET_B_c_1267_n N_A_1972_21#_c_1575_n 0.0219708f $X=11.26 $Y=0.85
+ $X2=0 $Y2=0
cc_947 N_RESET_B_c_1257_n N_A_1972_21#_c_1577_n 0.0163069f $X=11.065 $Y=1.17
+ $X2=0 $Y2=0
cc_948 N_RESET_B_c_1262_n N_A_1972_21#_c_1577_n 0.0023744f $X=10.92 $Y=1.17
+ $X2=0 $Y2=0
cc_949 N_RESET_B_c_1267_n N_A_1972_21#_c_1577_n 0.00506212f $X=11.26 $Y=0.85
+ $X2=0 $Y2=0
cc_950 N_RESET_B_M1006_g N_A_1972_21#_c_1578_n 0.0209838f $X=10.71 $Y=0.445
+ $X2=0 $Y2=0
cc_951 N_RESET_B_c_1257_n N_A_1972_21#_c_1578_n 5.583e-19 $X=11.065 $Y=1.17
+ $X2=0 $Y2=0
cc_952 N_RESET_B_c_1260_n N_A_1972_21#_c_1578_n 0.00636935f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_953 RESET_B N_A_1972_21#_c_1578_n 7.17527e-19 $X=11.185 $Y=0.765 $X2=0 $Y2=0
cc_954 N_RESET_B_c_1270_n N_A_1757_47#_c_1758_n 0.0296859f $X=10.735 $Y=1.89
+ $X2=0 $Y2=0
cc_955 N_RESET_B_c_1271_n N_A_1757_47#_c_1758_n 0.0110716f $X=10.735 $Y=1.99
+ $X2=0 $Y2=0
cc_956 N_RESET_B_c_1257_n N_A_1757_47#_c_1758_n 0.0023746f $X=11.065 $Y=1.17
+ $X2=0 $Y2=0
cc_957 N_RESET_B_c_1262_n N_A_1757_47#_c_1758_n 5.7962e-19 $X=10.92 $Y=1.17
+ $X2=0 $Y2=0
cc_958 N_RESET_B_M1006_g N_A_1757_47#_c_1754_n 0.00423781f $X=10.71 $Y=0.445
+ $X2=0 $Y2=0
cc_959 N_RESET_B_c_1270_n N_A_1757_47#_c_1754_n 0.00796937f $X=10.735 $Y=1.89
+ $X2=0 $Y2=0
cc_960 N_RESET_B_c_1257_n N_A_1757_47#_c_1754_n 0.0108565f $X=11.065 $Y=1.17
+ $X2=0 $Y2=0
cc_961 N_RESET_B_c_1262_n N_A_1757_47#_c_1754_n 5.5375e-19 $X=10.92 $Y=1.17
+ $X2=0 $Y2=0
cc_962 RESET_B N_A_1757_47#_c_1754_n 0.00121136f $X=11.185 $Y=0.765 $X2=0 $Y2=0
cc_963 N_RESET_B_c_1266_n N_A_1757_47#_c_1754_n 0.018989f $X=10.77 $Y=1.15 $X2=0
+ $Y2=0
cc_964 N_RESET_B_c_1267_n N_A_1757_47#_c_1754_n 0.00609004f $X=11.26 $Y=0.85
+ $X2=0 $Y2=0
cc_965 N_RESET_B_M1006_g N_A_1757_47#_c_1755_n 0.028267f $X=10.71 $Y=0.445 $X2=0
+ $Y2=0
cc_966 N_RESET_B_c_1267_n N_A_1757_47#_c_1755_n 0.0055381f $X=11.26 $Y=0.85
+ $X2=0 $Y2=0
cc_967 RESET_B N_A_1757_47#_c_1756_n 9.94285e-19 $X=11.185 $Y=0.765 $X2=0 $Y2=0
cc_968 N_RESET_B_c_1267_n N_A_1757_47#_c_1756_n 0.00643617f $X=11.26 $Y=0.85
+ $X2=0 $Y2=0
cc_969 N_RESET_B_c_1260_n N_A_1757_47#_c_1764_n 0.0185721f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_970 N_RESET_B_c_1271_n N_A_1757_47#_c_1767_n 2.91724e-19 $X=10.735 $Y=1.99
+ $X2=0 $Y2=0
cc_971 N_RESET_B_c_1260_n N_A_1757_47#_c_1757_n 0.0278903f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_972 N_RESET_B_c_1270_n N_A_1757_47#_c_1761_n 0.00133935f $X=10.735 $Y=1.89
+ $X2=0 $Y2=0
cc_973 N_RESET_B_c_1271_n N_A_1757_47#_c_1761_n 7.30168e-19 $X=10.735 $Y=1.99
+ $X2=0 $Y2=0
cc_974 N_RESET_B_c_1270_n N_A_1757_47#_c_1762_n 0.00550928f $X=10.735 $Y=1.89
+ $X2=0 $Y2=0
cc_975 N_RESET_B_c_1260_n N_A_1757_47#_c_1762_n 0.00960106f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_976 N_RESET_B_c_1270_n N_A_1757_47#_c_1763_n 0.0188936f $X=10.735 $Y=1.89
+ $X2=0 $Y2=0
cc_977 N_RESET_B_c_1257_n N_A_1757_47#_c_1763_n 0.0318741f $X=11.065 $Y=1.17
+ $X2=0 $Y2=0
cc_978 N_RESET_B_c_1262_n N_A_1757_47#_c_1763_n 0.00809733f $X=10.92 $Y=1.17
+ $X2=0 $Y2=0
cc_979 RESET_B N_A_1757_47#_c_1763_n 0.00111646f $X=11.185 $Y=0.765 $X2=0 $Y2=0
cc_980 N_RESET_B_c_1266_n N_A_1757_47#_c_1763_n 0.00225267f $X=10.77 $Y=1.15
+ $X2=0 $Y2=0
cc_981 N_RESET_B_c_1269_n N_VPWR_c_1873_n 0.0055115f $X=7.62 $Y=1.99 $X2=0 $Y2=0
cc_982 N_RESET_B_c_1271_n N_VPWR_c_1874_n 0.00839123f $X=10.735 $Y=1.99 $X2=0
+ $Y2=0
cc_983 N_RESET_B_c_1271_n N_VPWR_c_1875_n 0.00643335f $X=10.735 $Y=1.99 $X2=0
+ $Y2=0
cc_984 N_RESET_B_c_1269_n N_VPWR_c_1884_n 0.00639631f $X=7.62 $Y=1.99 $X2=0
+ $Y2=0
cc_985 N_RESET_B_c_1269_n N_VPWR_c_1891_n 0.00512994f $X=7.62 $Y=1.99 $X2=0
+ $Y2=0
cc_986 N_RESET_B_c_1271_n N_VPWR_c_1896_n 7.66292e-19 $X=10.735 $Y=1.99 $X2=0
+ $Y2=0
cc_987 N_RESET_B_c_1269_n N_VPWR_c_1869_n 0.00808107f $X=7.62 $Y=1.99 $X2=0
+ $Y2=0
cc_988 N_RESET_B_c_1271_n N_VPWR_c_1869_n 0.0108488f $X=10.735 $Y=1.99 $X2=0
+ $Y2=0
cc_989 N_RESET_B_c_1269_n N_A_1324_413#_c_2177_n 0.0133899f $X=7.62 $Y=1.99
+ $X2=0 $Y2=0
cc_990 N_RESET_B_c_1269_n N_A_1324_413#_c_2179_n 0.00113575f $X=7.62 $Y=1.99
+ $X2=0 $Y2=0
cc_991 N_RESET_B_c_1260_n N_VGND_M1022_d 0.00359137f $X=10.775 $Y=0.85 $X2=0
+ $Y2=0
cc_992 N_RESET_B_c_1261_n N_VGND_M1022_d 7.69682e-19 $X=7.9 $Y=0.85 $X2=0 $Y2=0
cc_993 N_RESET_B_c_1258_n N_VGND_c_2252_n 0.00321159f $X=7.785 $Y=0.85 $X2=0
+ $Y2=0
cc_994 N_RESET_B_c_1259_n N_VGND_c_2252_n 0.00640958f $X=7.7 $Y=0.85 $X2=0 $Y2=0
cc_995 N_RESET_B_c_1260_n N_VGND_c_2252_n 0.00202686f $X=10.775 $Y=0.85 $X2=0
+ $Y2=0
cc_996 N_RESET_B_c_1264_n N_VGND_c_2252_n 5.41848e-19 $X=7.535 $Y=0.96 $X2=0
+ $Y2=0
cc_997 N_RESET_B_c_1265_n N_VGND_c_2252_n 0.0112955f $X=7.56 $Y=0.755 $X2=0
+ $Y2=0
cc_998 N_RESET_B_M1006_g N_VGND_c_2253_n 0.00398835f $X=10.71 $Y=0.445 $X2=0
+ $Y2=0
cc_999 N_RESET_B_c_1260_n N_VGND_c_2253_n 0.00211161f $X=10.775 $Y=0.85 $X2=0
+ $Y2=0
cc_1000 N_RESET_B_c_1264_n N_VGND_c_2258_n 0.00173251f $X=7.535 $Y=0.96 $X2=0
+ $Y2=0
cc_1001 N_RESET_B_c_1265_n N_VGND_c_2258_n 0.00585385f $X=7.56 $Y=0.755 $X2=0
+ $Y2=0
cc_1002 N_RESET_B_M1006_g N_VGND_c_2262_n 0.00365983f $X=10.71 $Y=0.445 $X2=0
+ $Y2=0
cc_1003 N_RESET_B_M1006_g N_VGND_c_2275_n 0.00609608f $X=10.71 $Y=0.445 $X2=0
+ $Y2=0
cc_1004 N_RESET_B_c_1258_n N_VGND_c_2275_n 0.0413117f $X=7.785 $Y=0.85 $X2=0
+ $Y2=0
cc_1005 N_RESET_B_c_1259_n N_VGND_c_2275_n 0.00508167f $X=7.7 $Y=0.85 $X2=0
+ $Y2=0
cc_1006 N_RESET_B_c_1260_n N_VGND_c_2275_n 0.155008f $X=10.775 $Y=0.85 $X2=0
+ $Y2=0
cc_1007 RESET_B N_VGND_c_2275_n 0.0145638f $X=11.185 $Y=0.765 $X2=0 $Y2=0
cc_1008 N_RESET_B_c_1264_n N_VGND_c_2275_n 8.48191e-19 $X=7.535 $Y=0.96 $X2=0
+ $Y2=0
cc_1009 N_RESET_B_c_1265_n N_VGND_c_2275_n 0.00637693f $X=7.56 $Y=0.755 $X2=0
+ $Y2=0
cc_1010 N_A_1202_413#_c_1429_n N_VPWR_c_1873_n 5.18369e-19 $X=8.57 $Y=1.495
+ $X2=0 $Y2=0
cc_1011 N_A_1202_413#_c_1430_n N_VPWR_c_1873_n 0.00509065f $X=8.66 $Y=1.57 $X2=0
+ $Y2=0
cc_1012 N_A_1202_413#_c_1428_n N_VPWR_c_1873_n 4.68276e-19 $X=8.065 $Y=1.17
+ $X2=0 $Y2=0
cc_1013 N_A_1202_413#_c_1447_n N_VPWR_c_1885_n 0.0227799f $X=6.295 $Y=2.33 $X2=0
+ $Y2=0
cc_1014 N_A_1202_413#_c_1430_n N_VPWR_c_1886_n 0.00522999f $X=8.66 $Y=1.57 $X2=0
+ $Y2=0
cc_1015 N_A_1202_413#_M1025_d N_VPWR_c_1869_n 0.00305741f $X=6.01 $Y=2.065 $X2=0
+ $Y2=0
cc_1016 N_A_1202_413#_c_1430_n N_VPWR_c_1869_n 0.00772129f $X=8.66 $Y=1.57 $X2=0
+ $Y2=0
cc_1017 N_A_1202_413#_c_1447_n N_VPWR_c_1869_n 0.00637846f $X=6.295 $Y=2.33
+ $X2=0 $Y2=0
cc_1018 N_A_1202_413#_c_1447_n N_A_700_389#_c_2079_n 0.0168471f $X=6.295 $Y=2.33
+ $X2=0 $Y2=0
cc_1019 N_A_1202_413#_c_1433_n N_A_700_389#_c_2079_n 0.00498523f $X=6.277
+ $Y=2.135 $X2=0 $Y2=0
cc_1020 N_A_1202_413#_c_1434_n N_A_1324_413#_c_2177_n 0.00204762f $X=6.925
+ $Y=1.3 $X2=0 $Y2=0
cc_1021 N_A_1202_413#_c_1423_n N_A_1324_413#_c_2178_n 0.00297929f $X=6.84 $Y=1.3
+ $X2=0 $Y2=0
cc_1022 N_A_1202_413#_c_1433_n N_A_1324_413#_c_2178_n 0.0260688f $X=6.277
+ $Y=2.135 $X2=0 $Y2=0
cc_1023 N_A_1202_413#_c_1430_n N_A_1324_413#_c_2179_n 0.00360997f $X=8.66
+ $Y=1.57 $X2=0 $Y2=0
cc_1024 N_A_1202_413#_M1041_g N_VGND_c_2252_n 0.00655088f $X=8.235 $Y=0.555
+ $X2=0 $Y2=0
cc_1025 N_A_1202_413#_c_1426_n N_VGND_c_2252_n 0.00205385f $X=7.98 $Y=1.3 $X2=0
+ $Y2=0
cc_1026 N_A_1202_413#_c_1427_n N_VGND_c_2252_n 6.81471e-19 $X=8.065 $Y=1.17
+ $X2=0 $Y2=0
cc_1027 N_A_1202_413#_c_1428_n N_VGND_c_2252_n 0.00132464f $X=8.065 $Y=1.17
+ $X2=0 $Y2=0
cc_1028 N_A_1202_413#_c_1462_n N_VGND_c_2258_n 0.0398571f $X=6.84 $Y=0.39 $X2=0
+ $Y2=0
cc_1029 N_A_1202_413#_M1041_g N_VGND_c_2260_n 0.00467644f $X=8.235 $Y=0.555
+ $X2=0 $Y2=0
cc_1030 N_A_1202_413#_M1010_d N_VGND_c_2275_n 0.00348136f $X=6.06 $Y=0.235 $X2=0
+ $Y2=0
cc_1031 N_A_1202_413#_M1041_g N_VGND_c_2275_n 0.00659132f $X=8.235 $Y=0.555
+ $X2=0 $Y2=0
cc_1032 N_A_1202_413#_c_1462_n N_VGND_c_2275_n 0.0318737f $X=6.84 $Y=0.39 $X2=0
+ $Y2=0
cc_1033 N_A_1202_413#_c_1462_n A_1322_47# 0.00955634f $X=6.84 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_1034 N_A_1202_413#_c_1425_n A_1322_47# 0.00216963f $X=6.925 $Y=1.215
+ $X2=-0.19 $Y2=-0.24
cc_1035 N_A_1972_21#_c_1588_n N_A_1757_47#_c_1758_n 0.0170837f $X=11.56 $Y=2
+ $X2=0 $Y2=0
cc_1036 N_A_1972_21#_c_1589_n N_A_1757_47#_c_1758_n 8.84497e-19 $X=11.08 $Y=2
+ $X2=0 $Y2=0
cc_1037 N_A_1972_21#_c_1590_n N_A_1757_47#_c_1758_n 0.0029852f $X=11.645
+ $Y=1.915 $X2=0 $Y2=0
cc_1038 N_A_1972_21#_c_1565_n N_A_1757_47#_c_1754_n 0.00408921f $X=12.325
+ $Y=1.16 $X2=0 $Y2=0
cc_1039 N_A_1972_21#_c_1590_n N_A_1757_47#_c_1754_n 0.0156075f $X=11.645
+ $Y=1.915 $X2=0 $Y2=0
cc_1040 N_A_1972_21#_c_1577_n N_A_1757_47#_c_1754_n 0.00426472f $X=11.647
+ $Y=1.16 $X2=0 $Y2=0
cc_1041 N_A_1972_21#_c_1571_n N_A_1757_47#_c_1755_n 2.25605e-19 $X=10.56 $Y=0.78
+ $X2=0 $Y2=0
cc_1042 N_A_1972_21#_c_1573_n N_A_1757_47#_c_1755_n 9.93751e-19 $X=10.645
+ $Y=0.695 $X2=0 $Y2=0
cc_1043 N_A_1972_21#_c_1574_n N_A_1757_47#_c_1755_n 0.00813009f $X=11.56 $Y=0.38
+ $X2=0 $Y2=0
cc_1044 N_A_1972_21#_c_1575_n N_A_1757_47#_c_1755_n 0.00397992f $X=11.647
+ $Y=0.995 $X2=0 $Y2=0
cc_1045 N_A_1972_21#_c_1574_n N_A_1757_47#_c_1756_n 6.86779e-19 $X=11.56 $Y=0.38
+ $X2=0 $Y2=0
cc_1046 N_A_1972_21#_c_1575_n N_A_1757_47#_c_1756_n 0.00441406f $X=11.647
+ $Y=0.995 $X2=0 $Y2=0
cc_1047 N_A_1972_21#_M1032_g N_A_1757_47#_c_1764_n 0.00892221f $X=9.935 $Y=0.445
+ $X2=0 $Y2=0
cc_1048 N_A_1972_21#_c_1573_n N_A_1757_47#_c_1764_n 2.62721e-19 $X=10.645
+ $Y=0.695 $X2=0 $Y2=0
cc_1049 N_A_1972_21#_c_1580_n N_A_1757_47#_c_1767_n 0.0128301f $X=10.175 $Y=1.99
+ $X2=0 $Y2=0
cc_1050 N_A_1972_21#_M1032_g N_A_1757_47#_c_1757_n 0.00864444f $X=9.935 $Y=0.445
+ $X2=0 $Y2=0
cc_1051 N_A_1972_21#_c_1570_n N_A_1757_47#_c_1757_n 0.0142137f $X=10.235 $Y=0.98
+ $X2=0 $Y2=0
cc_1052 N_A_1972_21#_c_1572_n N_A_1757_47#_c_1757_n 0.00860636f $X=10.37 $Y=0.78
+ $X2=0 $Y2=0
cc_1053 N_A_1972_21#_c_1573_n N_A_1757_47#_c_1757_n 0.00389347f $X=10.645
+ $Y=0.695 $X2=0 $Y2=0
cc_1054 N_A_1972_21#_c_1578_n N_A_1757_47#_c_1757_n 0.0111004f $X=10.175 $Y=0.98
+ $X2=0 $Y2=0
cc_1055 N_A_1972_21#_c_1562_n N_A_1757_47#_c_1761_n 0.00450023f $X=10.175
+ $Y=1.89 $X2=0 $Y2=0
cc_1056 N_A_1972_21#_c_1580_n N_A_1757_47#_c_1761_n 0.00777832f $X=10.175
+ $Y=1.99 $X2=0 $Y2=0
cc_1057 N_A_1972_21#_c_1562_n N_A_1757_47#_c_1762_n 0.0235271f $X=10.175 $Y=1.89
+ $X2=0 $Y2=0
cc_1058 N_A_1972_21#_c_1570_n N_A_1757_47#_c_1762_n 0.0102912f $X=10.235 $Y=0.98
+ $X2=0 $Y2=0
cc_1059 N_A_1972_21#_c_1578_n N_A_1757_47#_c_1762_n 0.0062359f $X=10.175 $Y=0.98
+ $X2=0 $Y2=0
cc_1060 N_A_1972_21#_c_1570_n N_A_1757_47#_c_1763_n 0.00321233f $X=10.235
+ $Y=0.98 $X2=0 $Y2=0
cc_1061 N_A_1972_21#_c_1588_n N_A_1757_47#_c_1763_n 0.019955f $X=11.56 $Y=2
+ $X2=0 $Y2=0
cc_1062 N_A_1972_21#_c_1589_n N_A_1757_47#_c_1763_n 0.0134565f $X=11.08 $Y=2
+ $X2=0 $Y2=0
cc_1063 N_A_1972_21#_c_1590_n N_A_1757_47#_c_1763_n 0.0123382f $X=11.645
+ $Y=1.915 $X2=0 $Y2=0
cc_1064 N_A_1972_21#_c_1578_n N_A_1757_47#_c_1763_n 0.00193244f $X=10.175
+ $Y=0.98 $X2=0 $Y2=0
cc_1065 N_A_1972_21#_c_1588_n N_VPWR_M1011_d 0.00226776f $X=11.56 $Y=2 $X2=0
+ $Y2=0
cc_1066 N_A_1972_21#_c_1580_n N_VPWR_c_1874_n 0.0049242f $X=10.175 $Y=1.99 $X2=0
+ $Y2=0
cc_1067 N_A_1972_21#_c_1669_p N_VPWR_c_1874_n 0.00982513f $X=10.995 $Y=2.21
+ $X2=0 $Y2=0
cc_1068 N_A_1972_21#_c_1669_p N_VPWR_c_1875_n 0.00725596f $X=10.995 $Y=2.21
+ $X2=0 $Y2=0
cc_1069 N_A_1972_21#_c_1588_n N_VPWR_c_1875_n 0.00248346f $X=11.56 $Y=2 $X2=0
+ $Y2=0
cc_1070 N_A_1972_21#_c_1581_n N_VPWR_c_1876_n 0.0196928f $X=12.225 $Y=1.41 $X2=0
+ $Y2=0
cc_1071 N_A_1972_21#_c_1565_n N_VPWR_c_1876_n 0.00311818f $X=12.325 $Y=1.16
+ $X2=0 $Y2=0
cc_1072 N_A_1972_21#_c_1584_n N_VPWR_c_1876_n 0.00183303f $X=12.76 $Y=1.41 $X2=0
+ $Y2=0
cc_1073 N_A_1972_21#_c_1588_n N_VPWR_c_1876_n 0.0141977f $X=11.56 $Y=2 $X2=0
+ $Y2=0
cc_1074 N_A_1972_21#_c_1590_n N_VPWR_c_1876_n 0.0312705f $X=11.645 $Y=1.915
+ $X2=0 $Y2=0
cc_1075 N_A_1972_21#_c_1576_n N_VPWR_c_1876_n 0.018152f $X=12.12 $Y=1.16 $X2=0
+ $Y2=0
cc_1076 N_A_1972_21#_c_1584_n N_VPWR_c_1877_n 0.0130562f $X=12.76 $Y=1.41 $X2=0
+ $Y2=0
cc_1077 N_A_1972_21#_c_1585_n N_VPWR_c_1877_n 0.0174189f $X=13.295 $Y=1.41 $X2=0
+ $Y2=0
cc_1078 N_A_1972_21#_c_1586_n N_VPWR_c_1877_n 0.00192429f $X=13.765 $Y=1.41
+ $X2=0 $Y2=0
cc_1079 N_A_1972_21#_c_1569_n N_VPWR_c_1877_n 0.00523068f $X=13.765 $Y=1.202
+ $X2=0 $Y2=0
cc_1080 N_A_1972_21#_c_1586_n N_VPWR_c_1879_n 0.0109796f $X=13.765 $Y=1.41 $X2=0
+ $Y2=0
cc_1081 N_A_1972_21#_c_1580_n N_VPWR_c_1886_n 0.00528089f $X=10.175 $Y=1.99
+ $X2=0 $Y2=0
cc_1082 N_A_1972_21#_c_1588_n N_VPWR_c_1888_n 0.00192891f $X=11.56 $Y=2 $X2=0
+ $Y2=0
cc_1083 N_A_1972_21#_c_1581_n N_VPWR_c_1892_n 0.00622633f $X=12.225 $Y=1.41
+ $X2=0 $Y2=0
cc_1084 N_A_1972_21#_c_1584_n N_VPWR_c_1892_n 0.00590376f $X=12.76 $Y=1.41 $X2=0
+ $Y2=0
cc_1085 N_A_1972_21#_c_1585_n N_VPWR_c_1893_n 0.00622633f $X=13.295 $Y=1.41
+ $X2=0 $Y2=0
cc_1086 N_A_1972_21#_c_1586_n N_VPWR_c_1893_n 0.00677109f $X=13.765 $Y=1.41
+ $X2=0 $Y2=0
cc_1087 N_A_1972_21#_c_1581_n N_VPWR_c_1896_n 9.66739e-19 $X=12.225 $Y=1.41
+ $X2=0 $Y2=0
cc_1088 N_A_1972_21#_c_1669_p N_VPWR_c_1896_n 0.00875981f $X=10.995 $Y=2.21
+ $X2=0 $Y2=0
cc_1089 N_A_1972_21#_c_1588_n N_VPWR_c_1896_n 0.0247989f $X=11.56 $Y=2 $X2=0
+ $Y2=0
cc_1090 N_A_1972_21#_M1004_d N_VPWR_c_1869_n 0.00560711f $X=10.825 $Y=2.065
+ $X2=0 $Y2=0
cc_1091 N_A_1972_21#_c_1580_n N_VPWR_c_1869_n 0.00858035f $X=10.175 $Y=1.99
+ $X2=0 $Y2=0
cc_1092 N_A_1972_21#_c_1581_n N_VPWR_c_1869_n 0.0106417f $X=12.225 $Y=1.41 $X2=0
+ $Y2=0
cc_1093 N_A_1972_21#_c_1584_n N_VPWR_c_1869_n 0.0100476f $X=12.76 $Y=1.41 $X2=0
+ $Y2=0
cc_1094 N_A_1972_21#_c_1585_n N_VPWR_c_1869_n 0.010479f $X=13.295 $Y=1.41 $X2=0
+ $Y2=0
cc_1095 N_A_1972_21#_c_1586_n N_VPWR_c_1869_n 0.0128111f $X=13.765 $Y=1.41 $X2=0
+ $Y2=0
cc_1096 N_A_1972_21#_c_1669_p N_VPWR_c_1869_n 0.00608739f $X=10.995 $Y=2.21
+ $X2=0 $Y2=0
cc_1097 N_A_1972_21#_c_1588_n N_VPWR_c_1869_n 0.0090279f $X=11.56 $Y=2 $X2=0
+ $Y2=0
cc_1098 N_A_1972_21#_c_1569_n N_Q_c_2214_n 0.0692163f $X=13.765 $Y=1.202 $X2=0
+ $Y2=0
cc_1099 N_A_1972_21#_c_1567_n N_Q_c_2210_n 0.0039527f $X=13.32 $Y=0.995 $X2=0
+ $Y2=0
cc_1100 N_A_1972_21#_c_1568_n N_Q_c_2210_n 0.00413525f $X=13.79 $Y=0.995 $X2=0
+ $Y2=0
cc_1101 N_A_1972_21#_c_1585_n N_Q_c_2212_n 0.00592525f $X=13.295 $Y=1.41 $X2=0
+ $Y2=0
cc_1102 N_A_1972_21#_c_1586_n N_Q_c_2212_n 0.0160608f $X=13.765 $Y=1.41 $X2=0
+ $Y2=0
cc_1103 N_A_1972_21#_c_1569_n N_Q_c_2212_n 0.00679626f $X=13.765 $Y=1.202 $X2=0
+ $Y2=0
cc_1104 N_A_1972_21#_c_1564_n N_Q_c_2220_n 0.0242284f $X=12.66 $Y=1.16 $X2=0
+ $Y2=0
cc_1105 N_A_1972_21#_c_1569_n N_Q_c_2220_n 0.00332539f $X=13.765 $Y=1.202 $X2=0
+ $Y2=0
cc_1106 N_A_1972_21#_c_1576_n N_Q_c_2220_n 0.022453f $X=12.12 $Y=1.16 $X2=0
+ $Y2=0
cc_1107 N_A_1972_21#_c_1569_n N_Q_c_2223_n 0.0316582f $X=13.765 $Y=1.202 $X2=0
+ $Y2=0
cc_1108 N_A_1972_21#_c_1563_n Q 0.0147804f $X=12.2 $Y=0.995 $X2=0 $Y2=0
cc_1109 N_A_1972_21#_c_1566_n Q 0.00798032f $X=12.84 $Y=0.995 $X2=0 $Y2=0
cc_1110 N_A_1972_21#_c_1581_n Q 0.00650237f $X=12.225 $Y=1.41 $X2=0 $Y2=0
cc_1111 N_A_1972_21#_c_1565_n Q 0.00223846f $X=12.325 $Y=1.16 $X2=0 $Y2=0
cc_1112 N_A_1972_21#_c_1584_n Q 0.0191366f $X=12.76 $Y=1.41 $X2=0 $Y2=0
cc_1113 N_A_1972_21#_c_1585_n Q 4.00483e-19 $X=13.295 $Y=1.41 $X2=0 $Y2=0
cc_1114 N_A_1972_21#_c_1569_n Q 0.00368786f $X=13.765 $Y=1.202 $X2=0 $Y2=0
cc_1115 N_A_1972_21#_c_1573_n N_VGND_M1032_d 0.00294039f $X=10.645 $Y=0.695
+ $X2=0 $Y2=0
cc_1116 N_A_1972_21#_c_1626_n N_VGND_M1032_d 0.00211963f $X=10.73 $Y=0.38 $X2=0
+ $Y2=0
cc_1117 N_A_1972_21#_M1032_g N_VGND_c_2253_n 0.00417329f $X=9.935 $Y=0.445 $X2=0
+ $Y2=0
cc_1118 N_A_1972_21#_c_1572_n N_VGND_c_2253_n 0.0139752f $X=10.37 $Y=0.78 $X2=0
+ $Y2=0
cc_1119 N_A_1972_21#_c_1573_n N_VGND_c_2253_n 0.00352582f $X=10.645 $Y=0.695
+ $X2=0 $Y2=0
cc_1120 N_A_1972_21#_c_1626_n N_VGND_c_2253_n 0.0112461f $X=10.73 $Y=0.38 $X2=0
+ $Y2=0
cc_1121 N_A_1972_21#_c_1578_n N_VGND_c_2253_n 0.00234391f $X=10.175 $Y=0.98
+ $X2=0 $Y2=0
cc_1122 N_A_1972_21#_c_1563_n N_VGND_c_2254_n 0.00438629f $X=12.2 $Y=0.995 $X2=0
+ $Y2=0
cc_1123 N_A_1972_21#_c_1565_n N_VGND_c_2254_n 0.00169434f $X=12.325 $Y=1.16
+ $X2=0 $Y2=0
cc_1124 N_A_1972_21#_c_1574_n N_VGND_c_2254_n 0.0141315f $X=11.56 $Y=0.38 $X2=0
+ $Y2=0
cc_1125 N_A_1972_21#_c_1575_n N_VGND_c_2254_n 0.00589269f $X=11.647 $Y=0.995
+ $X2=0 $Y2=0
cc_1126 N_A_1972_21#_c_1576_n N_VGND_c_2254_n 0.00669683f $X=12.12 $Y=1.16 $X2=0
+ $Y2=0
cc_1127 N_A_1972_21#_c_1566_n N_VGND_c_2255_n 0.00423308f $X=12.84 $Y=0.995
+ $X2=0 $Y2=0
cc_1128 N_A_1972_21#_c_1567_n N_VGND_c_2255_n 0.00421175f $X=13.32 $Y=0.995
+ $X2=0 $Y2=0
cc_1129 N_A_1972_21#_c_1569_n N_VGND_c_2255_n 0.00268604f $X=13.765 $Y=1.202
+ $X2=0 $Y2=0
cc_1130 N_A_1972_21#_c_1568_n N_VGND_c_2257_n 0.00438629f $X=13.79 $Y=0.995
+ $X2=0 $Y2=0
cc_1131 N_A_1972_21#_M1032_g N_VGND_c_2260_n 0.00539841f $X=9.935 $Y=0.445 $X2=0
+ $Y2=0
cc_1132 N_A_1972_21#_c_1571_n N_VGND_c_2262_n 0.00305478f $X=10.56 $Y=0.78 $X2=0
+ $Y2=0
cc_1133 N_A_1972_21#_c_1572_n N_VGND_c_2262_n 6.89658e-19 $X=10.37 $Y=0.78 $X2=0
+ $Y2=0
cc_1134 N_A_1972_21#_c_1574_n N_VGND_c_2262_n 0.0477747f $X=11.56 $Y=0.38 $X2=0
+ $Y2=0
cc_1135 N_A_1972_21#_c_1626_n N_VGND_c_2262_n 0.00769222f $X=10.73 $Y=0.38 $X2=0
+ $Y2=0
cc_1136 N_A_1972_21#_c_1563_n N_VGND_c_2264_n 0.00585385f $X=12.2 $Y=0.995 $X2=0
+ $Y2=0
cc_1137 N_A_1972_21#_c_1566_n N_VGND_c_2264_n 0.00585385f $X=12.84 $Y=0.995
+ $X2=0 $Y2=0
cc_1138 N_A_1972_21#_c_1567_n N_VGND_c_2270_n 0.00585385f $X=13.32 $Y=0.995
+ $X2=0 $Y2=0
cc_1139 N_A_1972_21#_c_1568_n N_VGND_c_2270_n 0.00585385f $X=13.79 $Y=0.995
+ $X2=0 $Y2=0
cc_1140 N_A_1972_21#_M1012_d N_VGND_c_2275_n 0.00242029f $X=11.265 $Y=0.235
+ $X2=0 $Y2=0
cc_1141 N_A_1972_21#_M1032_g N_VGND_c_2275_n 0.00738016f $X=9.935 $Y=0.445 $X2=0
+ $Y2=0
cc_1142 N_A_1972_21#_c_1563_n N_VGND_c_2275_n 0.0124353f $X=12.2 $Y=0.995 $X2=0
+ $Y2=0
cc_1143 N_A_1972_21#_c_1566_n N_VGND_c_2275_n 0.0112853f $X=12.84 $Y=0.995 $X2=0
+ $Y2=0
cc_1144 N_A_1972_21#_c_1567_n N_VGND_c_2275_n 0.0110185f $X=13.32 $Y=0.995 $X2=0
+ $Y2=0
cc_1145 N_A_1972_21#_c_1568_n N_VGND_c_2275_n 0.011699f $X=13.79 $Y=0.995 $X2=0
+ $Y2=0
cc_1146 N_A_1972_21#_c_1571_n N_VGND_c_2275_n 0.00219209f $X=10.56 $Y=0.78 $X2=0
+ $Y2=0
cc_1147 N_A_1972_21#_c_1572_n N_VGND_c_2275_n 0.00103135f $X=10.37 $Y=0.78 $X2=0
+ $Y2=0
cc_1148 N_A_1972_21#_c_1574_n N_VGND_c_2275_n 0.0227282f $X=11.56 $Y=0.38 $X2=0
+ $Y2=0
cc_1149 N_A_1972_21#_c_1626_n N_VGND_c_2275_n 0.0028133f $X=10.73 $Y=0.38 $X2=0
+ $Y2=0
cc_1150 N_A_1972_21#_c_1578_n N_VGND_c_2275_n 5.84978e-19 $X=10.175 $Y=0.98
+ $X2=0 $Y2=0
cc_1151 N_A_1972_21#_c_1574_n A_2157_47# 0.00572931f $X=11.56 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_1152 N_A_1757_47#_c_1758_n N_VPWR_c_1874_n 7.07177e-19 $X=11.235 $Y=1.99
+ $X2=0 $Y2=0
cc_1153 N_A_1757_47#_c_1767_n N_VPWR_c_1874_n 0.019222f $X=10.04 $Y=2.295 $X2=0
+ $Y2=0
cc_1154 N_A_1757_47#_c_1763_n N_VPWR_c_1874_n 0.0086938f $X=11.18 $Y=1.66 $X2=0
+ $Y2=0
cc_1155 N_A_1757_47#_c_1758_n N_VPWR_c_1875_n 0.00315029f $X=11.235 $Y=1.99
+ $X2=0 $Y2=0
cc_1156 N_A_1757_47#_c_1758_n N_VPWR_c_1876_n 0.00425257f $X=11.235 $Y=1.99
+ $X2=0 $Y2=0
cc_1157 N_A_1757_47#_c_1767_n N_VPWR_c_1886_n 0.0603021f $X=10.04 $Y=2.295 $X2=0
+ $Y2=0
cc_1158 N_A_1757_47#_c_1758_n N_VPWR_c_1896_n 0.0113143f $X=11.235 $Y=1.99 $X2=0
+ $Y2=0
cc_1159 N_A_1757_47#_M1035_d N_VPWR_c_1869_n 0.00194481f $X=9.275 $Y=2.065 $X2=0
+ $Y2=0
cc_1160 N_A_1757_47#_c_1758_n N_VPWR_c_1869_n 0.00385472f $X=11.235 $Y=1.99
+ $X2=0 $Y2=0
cc_1161 N_A_1757_47#_c_1767_n N_VPWR_c_1869_n 0.0251419f $X=10.04 $Y=2.295 $X2=0
+ $Y2=0
cc_1162 N_A_1757_47#_c_1767_n A_1951_413# 0.00596016f $X=10.04 $Y=2.295
+ $X2=-0.19 $Y2=-0.24
cc_1163 N_A_1757_47#_c_1764_n N_VGND_c_2253_n 0.0176949f $X=9.67 $Y=0.395 $X2=0
+ $Y2=0
cc_1164 N_A_1757_47#_c_1755_n N_VGND_c_2254_n 0.00215654f $X=11.245 $Y=0.73
+ $X2=0 $Y2=0
cc_1165 N_A_1757_47#_c_1764_n N_VGND_c_2260_n 0.0662357f $X=9.67 $Y=0.395 $X2=0
+ $Y2=0
cc_1166 N_A_1757_47#_c_1755_n N_VGND_c_2262_n 0.00366111f $X=11.245 $Y=0.73
+ $X2=0 $Y2=0
cc_1167 N_A_1757_47#_M1028_d N_VGND_c_2275_n 0.00259616f $X=8.785 $Y=0.235 $X2=0
+ $Y2=0
cc_1168 N_A_1757_47#_c_1755_n N_VGND_c_2275_n 0.0066353f $X=11.245 $Y=0.73 $X2=0
+ $Y2=0
cc_1169 N_A_1757_47#_c_1764_n N_VGND_c_2275_n 0.0191758f $X=9.67 $Y=0.395 $X2=0
+ $Y2=0
cc_1170 N_A_1757_47#_c_1764_n A_1866_47# 0.0102613f $X=9.67 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_1171 N_A_1757_47#_c_1757_n A_1866_47# 0.00169576f $X=9.78 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_1172 N_VPWR_c_1869_n A_618_389# 0.00173928f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1173 N_VPWR_c_1869_n N_A_700_389#_M1020_d 0.00642194f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1174 N_VPWR_c_1869_n N_A_700_389#_M1025_s 0.00256642f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1175 N_VPWR_c_1882_n N_A_700_389#_c_2110_n 0.0118139f $X=4.855 $Y=2.72 $X2=0
+ $Y2=0
cc_1176 N_VPWR_c_1869_n N_A_700_389#_c_2110_n 0.00308197f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1177 N_VPWR_M1007_d N_A_700_389#_c_2086_n 0.00246822f $X=4.895 $Y=1.945 $X2=0
+ $Y2=0
cc_1178 N_VPWR_c_1872_n N_A_700_389#_c_2086_n 0.015761f $X=5.04 $Y=2.36 $X2=0
+ $Y2=0
cc_1179 N_VPWR_c_1882_n N_A_700_389#_c_2086_n 0.0130728f $X=4.855 $Y=2.72 $X2=0
+ $Y2=0
cc_1180 N_VPWR_c_1869_n N_A_700_389#_c_2086_n 0.0101862f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1181 N_VPWR_M1007_d N_A_700_389#_c_2079_n 8.75701e-19 $X=4.895 $Y=1.945 $X2=0
+ $Y2=0
cc_1182 N_VPWR_c_1872_n N_A_700_389#_c_2079_n 0.0145016f $X=5.04 $Y=2.36 $X2=0
+ $Y2=0
cc_1183 N_VPWR_c_1885_n N_A_700_389#_c_2079_n 0.0247694f $X=7.135 $Y=2.72 $X2=0
+ $Y2=0
cc_1184 N_VPWR_c_1869_n N_A_700_389#_c_2079_n 0.0102483f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1185 N_VPWR_c_1869_n A_870_389# 0.00314879f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1186 N_VPWR_c_1869_n N_A_1324_413#_M1026_d 0.00251718f $X=14.03 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_1187 N_VPWR_c_1869_n N_A_1324_413#_M1023_d 0.00226832f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1188 N_VPWR_M1015_d N_A_1324_413#_c_2177_n 0.00406748f $X=7.09 $Y=2.065 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1884_n N_A_1324_413#_c_2177_n 0.0148301f $X=7.3 $Y=2.44 $X2=0
+ $Y2=0
cc_1190 N_VPWR_c_1885_n N_A_1324_413#_c_2177_n 0.00418739f $X=7.135 $Y=2.72
+ $X2=0 $Y2=0
cc_1191 N_VPWR_c_1891_n N_A_1324_413#_c_2177_n 0.0044576f $X=8.15 $Y=2.72 $X2=0
+ $Y2=0
cc_1192 N_VPWR_c_1869_n N_A_1324_413#_c_2177_n 0.00777578f $X=14.03 $Y=2.72
+ $X2=0 $Y2=0
cc_1193 N_VPWR_c_1885_n N_A_1324_413#_c_2178_n 0.00723406f $X=7.135 $Y=2.72
+ $X2=0 $Y2=0
cc_1194 N_VPWR_c_1869_n N_A_1324_413#_c_2178_n 0.00284468f $X=14.03 $Y=2.72
+ $X2=0 $Y2=0
cc_1195 N_VPWR_c_1873_n N_A_1324_413#_c_2179_n 0.013659f $X=8.425 $Y=2.34 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1884_n N_A_1324_413#_c_2179_n 9.9383e-19 $X=7.3 $Y=2.44 $X2=0
+ $Y2=0
cc_1197 N_VPWR_c_1891_n N_A_1324_413#_c_2179_n 0.00723406f $X=8.15 $Y=2.72 $X2=0
+ $Y2=0
cc_1198 N_VPWR_c_1869_n N_A_1324_413#_c_2179_n 0.00284468f $X=14.03 $Y=2.72
+ $X2=0 $Y2=0
cc_1199 N_VPWR_c_1869_n A_1951_413# 0.00258386f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1200 N_VPWR_c_1869_n N_Q_M1001_d 0.00687494f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1201 N_VPWR_c_1869_n N_Q_M1024_d 0.0046067f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1202 N_VPWR_c_1877_n N_Q_c_2214_n 0.0178273f $X=13.06 $Y=1.66 $X2=0 $Y2=0
cc_1203 N_VPWR_c_1877_n N_Q_c_2212_n 0.0506754f $X=13.06 $Y=1.66 $X2=0 $Y2=0
cc_1204 N_VPWR_c_1879_n N_Q_c_2212_n 0.0506754f $X=14 $Y=1.66 $X2=0 $Y2=0
cc_1205 N_VPWR_c_1893_n N_Q_c_2212_n 0.00807743f $X=13.915 $Y=2.72 $X2=0 $Y2=0
cc_1206 N_VPWR_c_1869_n N_Q_c_2212_n 0.00871977f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1207 N_VPWR_c_1876_n Q 0.0442947f $X=11.99 $Y=1.66 $X2=0 $Y2=0
cc_1208 N_VPWR_c_1877_n Q 0.0517323f $X=13.06 $Y=1.66 $X2=0 $Y2=0
cc_1209 N_VPWR_c_1892_n Q 0.0109048f $X=12.975 $Y=2.72 $X2=0 $Y2=0
cc_1210 N_VPWR_c_1869_n Q 0.011248f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1211 N_A_700_389#_c_2086_n A_870_389# 0.00431971f $X=5.14 $Y=2.02 $X2=-0.19
+ $Y2=-0.24
cc_1212 N_A_700_389#_c_2080_n N_VGND_M1038_d 2.35236e-19 $X=5.55 $Y=0.805 $X2=0
+ $Y2=0
cc_1213 N_A_700_389#_c_2081_n N_VGND_M1038_d 0.00246715f $X=5.31 $Y=0.805 $X2=0
+ $Y2=0
cc_1214 N_A_700_389#_c_2080_n N_VGND_c_2251_n 0.0029069f $X=5.55 $Y=0.805 $X2=0
+ $Y2=0
cc_1215 N_A_700_389#_c_2081_n N_VGND_c_2251_n 0.0138829f $X=5.31 $Y=0.805 $X2=0
+ $Y2=0
cc_1216 N_A_700_389#_c_2082_n N_VGND_c_2251_n 0.00248453f $X=5.635 $Y=0.715
+ $X2=0 $Y2=0
cc_1217 N_A_700_389#_c_2084_n N_VGND_c_2251_n 0.0126008f $X=5.725 $Y=0.42 $X2=0
+ $Y2=0
cc_1218 N_A_700_389#_c_2080_n N_VGND_c_2258_n 0.00310525f $X=5.55 $Y=0.805 $X2=0
+ $Y2=0
cc_1219 N_A_700_389#_c_2084_n N_VGND_c_2258_n 0.0136647f $X=5.725 $Y=0.42 $X2=0
+ $Y2=0
cc_1220 N_A_700_389#_M1010_s N_VGND_c_2275_n 0.00273547f $X=5.6 $Y=0.235 $X2=0
+ $Y2=0
cc_1221 N_A_700_389#_c_2080_n N_VGND_c_2275_n 0.00552288f $X=5.55 $Y=0.805 $X2=0
+ $Y2=0
cc_1222 N_A_700_389#_c_2081_n N_VGND_c_2275_n 7.57107e-19 $X=5.31 $Y=0.805 $X2=0
+ $Y2=0
cc_1223 N_A_700_389#_c_2084_n N_VGND_c_2275_n 0.0120347f $X=5.725 $Y=0.42 $X2=0
+ $Y2=0
cc_1224 N_Q_c_2214_n N_VGND_c_2255_n 0.00649431f $X=13.445 $Y=1.16 $X2=0 $Y2=0
cc_1225 Q N_VGND_c_2264_n 0.0201753f $X=12.565 $Y=0.425 $X2=0 $Y2=0
cc_1226 N_Q_c_2210_n N_VGND_c_2270_n 0.0150193f $X=13.53 $Y=0.63 $X2=0 $Y2=0
cc_1227 N_Q_M1013_s N_VGND_c_2275_n 0.00958453f $X=12.275 $Y=0.235 $X2=0 $Y2=0
cc_1228 N_Q_M1019_s N_VGND_c_2275_n 0.00507218f $X=13.395 $Y=0.235 $X2=0 $Y2=0
cc_1229 N_Q_c_2210_n N_VGND_c_2275_n 0.00950576f $X=13.53 $Y=0.63 $X2=0 $Y2=0
cc_1230 Q N_VGND_c_2275_n 0.0125721f $X=12.565 $Y=0.425 $X2=0 $Y2=0
cc_1231 N_VGND_c_2275_n A_1322_47# 0.00309919f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1232 N_VGND_c_2275_n A_1428_47# 0.00297921f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1233 N_VGND_c_2275_n A_1866_47# 0.00352964f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1234 N_VGND_c_2275_n A_2157_47# 0.0021994f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
