* File: sky130_fd_sc_hdll__muxb4to1_1.spice
* Created: Thu Aug 27 19:11:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__muxb4to1_1.pex.spice"
.subckt sky130_fd_sc_hdll__muxb4to1_1  VNB VPB D[0] S[0] S[1] D[1] D[2] S[2]
+ S[3] D[3] VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* D[3]	D[3]
* S[3]	S[3]
* S[2]	S[2]
* D[2]	D[2]
* D[1]	D[1]
* S[1]	S[1]
* S[0]	S[0]
* D[0]	D[0]
* VPB	VPB
* VNB	VNB
MM1021 A_109_47# N_D[0]_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.169 PD=1.08333 PS=1.82 NRD=21.636 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1023 N_Z_M1023_d N_S[0]_M1023_g A_109_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75000.7
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1017 N_VGND_M1017_d N_S[0]_M1017_g N_A_184_265#_M1017_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1016 N_A_533_47#_M1016_d N_S[1]_M1016_g N_VGND_M1017_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1006 A_746_47# N_S[1]_M1006_g N_Z_M1006_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1018 N_VGND_M1018_d N_D[1]_M1018_g A_746_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1000 A_937_47# N_D[2]_M1000_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_Z_M1004_d N_S[2]_M1004_g A_937_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1022 N_VGND_M1022_d N_S[2]_M1022_g N_A_1012_265#_M1022_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1015 N_A_1361_47#_M1015_d N_S[3]_M1015_g N_VGND_M1022_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1002 A_1574_47# N_S[3]_M1002_g N_Z_M1002_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.7 A=0.078 P=1.34 MULT=1
MM1020 N_VGND_M1020_d N_D[3]_M1020_g A_1574_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.111944 PD=1.82 PS=1.08333 NRD=0 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 A_117_297# N_D[0]_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.27 PD=1.47802 PS=2.54 NRD=24.8417 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_Z_M1009_d N_A_184_265#_M1009_g A_117_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90000.7 SB=90000.2 A=0.1476 P=2 MULT=1
MM1013 N_VPWR_M1013_d N_S[0]_M1013_g N_A_184_265#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1010 N_A_533_47#_M1010_d N_S[1]_M1010_g N_VPWR_M1013_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 A_734_333# N_A_533_47#_M1003_g N_Z_M1003_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1019 N_VPWR_M1019_d N_D[1]_M1019_g A_734_333# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1011 A_945_297# N_D[2]_M1011_g N_VPWR_M1019_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1012 N_Z_M1012_d N_A_1012_265#_M1012_g A_945_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1014 N_VPWR_M1014_d N_S[2]_M1014_g N_A_1012_265#_M1014_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1001 N_A_1361_47#_M1001_d N_S[3]_M1001_g N_VPWR_M1014_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 A_1562_333# N_A_1361_47#_M1005_g N_Z_M1005_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.7 A=0.1476 P=2 MULT=1
MM1008 N_VPWR_M1008_d N_D[3]_M1008_g A_1562_333# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.181154 PD=2.54 PS=1.47802 NRD=0.9653 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=14.6376 P=21.45
*
.include "sky130_fd_sc_hdll__muxb4to1_1.pxi.spice"
*
.ends
*
*
