* File: sky130_fd_sc_hdll__mux2i_2.spice
* Created: Thu Aug 27 19:11:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__mux2i_2.pex.spice"
.subckt sky130_fd_sc_hdll__mux2i_2  VNB VPB S A0 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_S_M1011_g N_A_27_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1002 N_A_213_47#_M1002_d N_S_M1002_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1016 N_A_213_47#_M1002_d N_S_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1016_s N_A_27_47#_M1008_g N_A_401_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_27_47#_M1012_g N_A_401_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_A0_M1000_g N_A_401_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_A0_M1003_g N_A_401_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.104 PD=0.96 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1007 N_A_213_47#_M1007_d N_A1_M1007_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.10075 PD=0.975 PS=0.96 NRD=8.304 NRS=6.456 M=1 R=4.33333
+ SA=75001.2 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1017 N_A_213_47#_M1007_d N_A1_M1017_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.32825 PD=0.975 PS=2.31 NRD=0 NRS=44.304 M=1 R=4.33333
+ SA=75001.6 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_S_M1005_g N_A_27_47#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1001 N_A_211_297#_M1001_d N_S_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1014 N_A_211_297#_M1001_d N_S_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1014_s N_A_27_47#_M1006_g N_A_399_297#_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_27_47#_M1009_g N_A_399_297#_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1004 N_A_211_297#_M1004_d N_A0_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1015 N_A_211_297#_M1004_d N_A0_M1015_g N_Y_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.165 PD=1.29 PS=1.33 NRD=0.9653 NRS=4.9053 M=1 R=5.55556
+ SA=90000.6 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1010 N_Y_M1015_s N_A1_M1010_g N_A_399_297#_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.165 AS=0.1475 PD=1.33 PS=1.295 NRD=4.9053 NRS=1.9503 M=1 R=5.55556
+ SA=90001.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1013 N_Y_M1013_d N_A1_M1013_g N_A_399_297#_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.465 AS=0.1475 PD=2.93 PS=1.295 NRD=1.9503 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.4 A=0.18 P=2.36 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.4695 P=15.01
c_43 VNB 0 1.34758e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hdll__mux2i_2.pxi.spice"
*
.ends
*
*
