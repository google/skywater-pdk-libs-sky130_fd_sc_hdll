* File: sky130_fd_sc_hdll__or4bb_4.pex.spice
* Created: Thu Aug 27 19:25:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%C_N 2 3 5 8 9 10 14 15 16
r35 14 17 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.16
+ $X2=0.535 $Y2=1.325
r36 14 16 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.16
+ $X2=0.535 $Y2=0.995
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.52
+ $Y=1.16 $X2=0.52 $Y2=1.16
r38 9 10 10.0469 $w=3.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.63 $Y=1.19 $X2=0.63
+ $Y2=1.53
r39 9 15 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=0.63 $Y=1.19 $X2=0.63
+ $Y2=1.16
r40 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.555 $Y=0.675
+ $X2=0.555 $Y2=0.995
r41 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.975
+ $X2=0.495 $Y2=2.26
r42 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.875 $X2=0.495
+ $Y2=1.975
r43 2 17 182.367 $w=2e-07 $l=5.5e-07 $layer=POLY_cond $X=0.495 $Y=1.875
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%D_N 1 3 4 6 7
r31 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.16 $X2=1.08 $Y2=1.16
r32 4 10 38.6069 $w=3.31e-07 $l=1.93533e-07 $layer=POLY_cond $X=1.05 $Y=0.995
+ $X2=1.112 $Y2=1.16
r33 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.05 $Y=0.995 $X2=1.05
+ $Y2=0.675
r34 1 10 46.3664 $w=3.31e-07 $l=2.88097e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.112 $Y2=1.16
r35 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.03 $Y=1.41 $X2=1.03
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%A_224_297# 1 2 7 9 10 12 13 14 15 22 24 27
+ 29
r65 27 30 7.92688 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=1.16
+ $X2=1.65 $Y2=1.325
r66 27 29 7.92688 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=1.16
+ $X2=1.65 $Y2=0.995
r67 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.16 $X2=1.71 $Y2=1.16
r68 24 25 17.5021 $w=2.37e-07 $l=3.4e-07 $layer=LI1_cond $X=1.26 $Y=0.655
+ $X2=1.6 $Y2=0.655
r69 22 30 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=1.6 $Y=1.56 $X2=1.6
+ $Y2=1.325
r70 19 25 2.03416 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=1.6 $Y=0.825 $X2=1.6
+ $Y2=0.655
r71 19 29 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=1.6 $Y=0.825 $X2=1.6
+ $Y2=0.995
r72 15 22 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.505 $Y=1.645
+ $X2=1.6 $Y2=1.56
r73 15 17 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.505 $Y=1.645
+ $X2=1.265 $Y2=1.645
r74 13 28 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.935 $Y=1.16
+ $X2=1.71 $Y2=1.16
r75 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.935 $Y=1.16
+ $X2=2.035 $Y2=1.202
r76 10 14 34.7346 $w=1.65e-07 $l=2.09485e-07 $layer=POLY_cond $X=2.04 $Y=0.995
+ $X2=2.035 $Y2=1.202
r77 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.04 $Y=0.995
+ $X2=2.04 $Y2=0.56
r78 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=2.035 $Y=1.41
+ $X2=2.035 $Y2=1.202
r79 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.035 $Y=1.41
+ $X2=2.035 $Y2=1.985
r80 2 17 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.645
r81 1 24 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.465 $X2=1.26 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%A_27_410# 1 2 7 9 10 12 14 17 19 22 23 24
+ 27 33 35
r81 30 33 3.53416 $w=3.73e-07 $l=1.15e-07 $layer=LI1_cond $X=0.18 $Y=0.637
+ $X2=0.295 $Y2=0.637
r82 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.16 $X2=2.48 $Y2=1.16
r83 25 27 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.48 $Y=2.295
+ $X2=2.48 $Y2=1.16
r84 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.395 $Y=2.38
+ $X2=2.48 $Y2=2.295
r85 23 24 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=2.395 $Y=2.38
+ $X2=1.395 $Y2=2.38
r86 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.31 $Y=2.295
+ $X2=1.395 $Y2=2.38
r87 21 22 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.31 $Y=2.07
+ $X2=1.31 $Y2=2.295
r88 20 35 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.345 $Y=1.985
+ $X2=0.22 $Y2=1.985
r89 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.225 $Y=1.985
+ $X2=1.31 $Y2=2.07
r90 19 20 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.225 $Y=1.985
+ $X2=0.345 $Y2=1.985
r91 15 35 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.22 $Y=2.07 $X2=0.22
+ $Y2=1.985
r92 15 17 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=0.22 $Y=2.07
+ $X2=0.22 $Y2=2.29
r93 14 35 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.18 $Y=1.9
+ $X2=0.22 $Y2=1.985
r94 13 30 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.18 $Y=0.825
+ $X2=0.18 $Y2=0.637
r95 13 14 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=0.18 $Y=0.825
+ $X2=0.18 $Y2=1.9
r96 10 28 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.505 $Y2=1.16
r97 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=0.56
r98 7 28 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.565 $Y=1.41
+ $X2=2.505 $Y2=1.16
r99 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.565 $Y=1.41
+ $X2=2.565 $Y2=1.985
r100 2 17 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r101 1 33 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.465 $X2=0.295 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%B 1 3 4 6 7 8 13
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.01
+ $Y=1.16 $X2=3.01 $Y2=1.16
r32 7 8 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=2.995 $Y=1.87 $X2=2.995
+ $Y2=2.21
r33 7 13 27.2745 $w=2.98e-07 $l=7.1e-07 $layer=LI1_cond $X=2.995 $Y=1.87
+ $X2=2.995 $Y2=1.16
r34 4 12 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.06 $Y=0.995
+ $X2=3.035 $Y2=1.16
r35 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.06 $Y=0.995 $X2=3.06
+ $Y2=0.56
r36 1 12 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.035 $Y=1.41
+ $X2=3.035 $Y2=1.16
r37 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.035 $Y=1.41
+ $X2=3.035 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%A 1 3 4 6 7 9 12 18
c38 7 0 1.93999e-19 $X=3.565 $Y=1.4
r39 12 18 1.07204 $w=2.13e-07 $l=2e-08 $layer=LI1_cond $X=3.45 $Y=1.507 $X2=3.47
+ $Y2=1.507
r40 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.54
+ $Y=1.16 $X2=3.54 $Y2=1.16
r41 7 18 5.09219 $w=2.13e-07 $l=9.5e-08 $layer=LI1_cond $X=3.565 $Y=1.507
+ $X2=3.47 $Y2=1.507
r42 7 9 12.5721 $w=2.18e-07 $l=2.4e-07 $layer=LI1_cond $X=3.565 $Y=1.4 $X2=3.565
+ $Y2=1.16
r43 4 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=3.505 $Y=1.41
+ $X2=3.565 $Y2=1.16
r44 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.505 $Y=1.41
+ $X2=3.505 $Y2=1.985
r45 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.48 $Y=0.995
+ $X2=3.565 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.48 $Y=0.995 $X2=3.48
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%A_335_297# 1 2 3 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 33 34 39 42 44 45 48 50 53 54 59 65 74
c148 74 0 1.93999e-19 $X=5.485 $Y=1.202
r149 74 75 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.485 $Y=1.202
+ $X2=5.51 $Y2=1.202
r150 71 72 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.99 $Y=1.202
+ $X2=5.015 $Y2=1.202
r151 70 71 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.545 $Y=1.202
+ $X2=4.99 $Y2=1.202
r152 69 70 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.52 $Y=1.202
+ $X2=4.545 $Y2=1.202
r153 66 67 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.05 $Y=1.202
+ $X2=4.075 $Y2=1.202
r154 62 64 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.13 $Y=0.74 $X2=2.33
+ $Y2=0.74
r155 60 74 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=5.28 $Y=1.202
+ $X2=5.485 $Y2=1.202
r156 60 72 34.336 $w=3.72e-07 $l=2.65e-07 $layer=POLY_cond $X=5.28 $Y=1.202
+ $X2=5.015 $Y2=1.202
r157 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.28
+ $Y=1.16 $X2=5.28 $Y2=1.16
r158 57 69 53.1237 $w=3.72e-07 $l=4.1e-07 $layer=POLY_cond $X=4.11 $Y=1.202
+ $X2=4.52 $Y2=1.202
r159 57 67 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=4.11 $Y=1.202
+ $X2=4.075 $Y2=1.202
r160 56 59 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.11 $Y=1.16
+ $X2=5.28 $Y2=1.16
r161 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.11
+ $Y=1.16 $X2=4.11 $Y2=1.16
r162 54 56 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.015 $Y=1.16
+ $X2=4.11 $Y2=1.16
r163 53 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.93 $Y=1.075
+ $X2=4.015 $Y2=1.16
r164 52 53 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.93 $Y=0.825
+ $X2=3.93 $Y2=1.075
r165 51 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=0.74
+ $X2=3.27 $Y2=0.74
r166 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.845 $Y=0.74
+ $X2=3.93 $Y2=0.825
r167 50 51 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.845 $Y=0.74
+ $X2=3.355 $Y2=0.74
r168 46 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.655
+ $X2=3.27 $Y2=0.74
r169 46 48 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.27 $Y=0.655
+ $X2=3.27 $Y2=0.49
r170 45 64 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=0.74
+ $X2=2.33 $Y2=0.74
r171 44 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0.74
+ $X2=3.27 $Y2=0.74
r172 44 45 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.185 $Y=0.74
+ $X2=2.415 $Y2=0.74
r173 40 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.33 $Y=0.655
+ $X2=2.33 $Y2=0.74
r174 40 42 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0.655
+ $X2=2.33 $Y2=0.49
r175 38 62 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=0.825
+ $X2=2.13 $Y2=0.74
r176 38 39 65.9617 $w=1.88e-07 $l=1.13e-06 $layer=LI1_cond $X=2.13 $Y=0.825
+ $X2=2.13 $Y2=1.955
r177 34 39 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.035 $Y=2.04
+ $X2=2.13 $Y2=1.955
r178 34 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.035 $Y=2.04
+ $X2=1.8 $Y2=2.04
r179 31 75 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.51 $Y=0.995
+ $X2=5.51 $Y2=1.202
r180 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.51 $Y=0.995
+ $X2=5.51 $Y2=0.56
r181 28 74 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.485 $Y=1.41
+ $X2=5.485 $Y2=1.202
r182 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.485 $Y=1.41
+ $X2=5.485 $Y2=1.985
r183 25 72 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.015 $Y=1.41
+ $X2=5.015 $Y2=1.202
r184 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.015 $Y=1.41
+ $X2=5.015 $Y2=1.985
r185 22 71 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.99 $Y=0.995
+ $X2=4.99 $Y2=1.202
r186 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.99 $Y=0.995
+ $X2=4.99 $Y2=0.56
r187 19 70 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.545 $Y=1.41
+ $X2=4.545 $Y2=1.202
r188 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.545 $Y=1.41
+ $X2=4.545 $Y2=1.985
r189 16 69 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.52 $Y=0.995
+ $X2=4.52 $Y2=1.202
r190 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.52 $Y=0.995
+ $X2=4.52 $Y2=0.56
r191 13 67 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.075 $Y=1.41
+ $X2=4.075 $Y2=1.202
r192 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.075 $Y=1.41
+ $X2=4.075 $Y2=1.985
r193 10 66 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.05 $Y=0.995
+ $X2=4.05 $Y2=1.202
r194 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.05 $Y=0.995
+ $X2=4.05 $Y2=0.56
r195 3 36 600 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=1 $X=1.675
+ $Y=1.485 $X2=1.8 $Y2=2.04
r196 2 48 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=3.135
+ $Y=0.235 $X2=3.27 $Y2=0.49
r197 1 42 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.235 $X2=2.33 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%VPWR 1 2 3 4 15 19 23 25 27 30 31 33 34 35
+ 37 52 57 61
r73 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r74 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 55 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r76 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r77 52 60 3.98688 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=5.787 $Y2=2.72
r78 52 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=5.29 $Y2=2.72
r79 51 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r80 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r81 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r82 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 45 48 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r84 45 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r85 44 47 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r86 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r87 42 57 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r88 42 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r89 37 57 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r90 37 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r91 35 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r92 35 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r93 33 50 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.655 $Y=2.72
+ $X2=4.37 $Y2=2.72
r94 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.655 $Y=2.72
+ $X2=4.78 $Y2=2.72
r95 32 54 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.905 $Y=2.72
+ $X2=5.29 $Y2=2.72
r96 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.905 $Y=2.72
+ $X2=4.78 $Y2=2.72
r97 30 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.66 $Y=2.72
+ $X2=3.45 $Y2=2.72
r98 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.66 $Y=2.72
+ $X2=3.785 $Y2=2.72
r99 29 50 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r100 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=3.785 $Y2=2.72
r101 25 60 3.15628 $w=2.5e-07 $l=1.13666e-07 $layer=LI1_cond $X=5.72 $Y=2.635
+ $X2=5.787 $Y2=2.72
r102 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.72 $Y=2.635
+ $X2=5.72 $Y2=1.96
r103 21 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=2.635
+ $X2=4.78 $Y2=2.72
r104 21 23 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.78 $Y=2.635
+ $X2=4.78 $Y2=1.96
r105 17 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=2.635
+ $X2=3.785 $Y2=2.72
r106 17 19 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.785 $Y=2.635
+ $X2=3.785 $Y2=1.96
r107 13 57 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r108 13 15 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.325
r109 4 27 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.575
+ $Y=1.485 $X2=5.72 $Y2=1.96
r110 3 23 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.635
+ $Y=1.485 $X2=4.78 $Y2=1.96
r111 2 19 300 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_PDIFF $count=2 $X=3.595
+ $Y=1.485 $X2=3.785 $Y2=1.96
r112 1 15 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.05 $X2=0.73 $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%X 1 2 3 4 13 15 19 21 23 24 27 31 33 35 39
+ 41 43 46
r77 43 46 3.05086 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=5.74 $Y=0.815 $X2=5.74
+ $Y2=0.905
r78 43 46 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.74 $Y=0.92
+ $X2=5.74 $Y2=0.905
r79 42 43 26.8068 $w=2.28e-07 $l=5.35e-07 $layer=LI1_cond $X=5.74 $Y=1.455
+ $X2=5.74 $Y2=0.92
r80 36 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.415 $Y=0.815
+ $X2=5.225 $Y2=0.815
r81 35 43 3.89832 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=5.625 $Y=0.815
+ $X2=5.74 $Y2=0.815
r82 35 36 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=5.625 $Y=0.815
+ $X2=5.415 $Y2=0.815
r83 34 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.375 $Y=1.54
+ $X2=5.25 $Y2=1.54
r84 33 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.625 $Y=1.54
+ $X2=5.74 $Y2=1.455
r85 33 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.625 $Y=1.54
+ $X2=5.375 $Y2=1.54
r86 29 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.25 $Y=1.625
+ $X2=5.25 $Y2=1.54
r87 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.25 $Y=1.625
+ $X2=5.25 $Y2=2.3
r88 25 39 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.225 $Y=0.725
+ $X2=5.225 $Y2=0.815
r89 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.225 $Y=0.725
+ $X2=5.225 $Y2=0.39
r90 23 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.035 $Y=0.815
+ $X2=5.225 $Y2=0.815
r91 23 24 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.035 $Y=0.815
+ $X2=4.475 $Y2=0.815
r92 22 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=1.54
+ $X2=4.31 $Y2=1.54
r93 21 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.125 $Y=1.54
+ $X2=5.25 $Y2=1.54
r94 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.125 $Y=1.54
+ $X2=4.435 $Y2=1.54
r95 17 24 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=4.35 $Y=0.725
+ $X2=4.475 $Y2=0.815
r96 17 19 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=4.35 $Y=0.725
+ $X2=4.35 $Y2=0.485
r97 13 38 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=1.625
+ $X2=4.31 $Y2=1.54
r98 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.31 $Y=1.625
+ $X2=4.31 $Y2=2.3
r99 4 41 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.105
+ $Y=1.485 $X2=5.25 $Y2=1.62
r100 4 31 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.105
+ $Y=1.485 $X2=5.25 $Y2=2.3
r101 3 38 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.165
+ $Y=1.485 $X2=4.31 $Y2=1.62
r102 3 15 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.165
+ $Y=1.485 $X2=4.31 $Y2=2.3
r103 2 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.065
+ $Y=0.235 $X2=5.25 $Y2=0.39
r104 1 19 182 $w=1.7e-07 $l=3.29773e-07 $layer=licon1_NDIFF $count=1 $X=4.125
+ $Y=0.235 $X2=4.31 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4BB_4%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44
+ 45 47 48 50 51 53 54 55 67 75 80 84
r102 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r103 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r104 78 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r105 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r106 75 83 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=5.635 $Y=0
+ $X2=5.807 $Y2=0
r107 75 77 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.635 $Y=0 $X2=5.29
+ $Y2=0
r108 74 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r109 74 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r110 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r111 71 80 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.805
+ $Y2=0
r112 71 73 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.995 $Y=0
+ $X2=4.37 $Y2=0
r113 70 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r114 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r115 67 80 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.805
+ $Y2=0
r116 67 69 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0
+ $X2=3.45 $Y2=0
r117 66 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r118 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r119 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r120 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r121 59 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r122 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r123 55 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r124 53 73 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.695 $Y=0
+ $X2=4.37 $Y2=0
r125 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=0 $X2=4.78
+ $Y2=0
r126 52 77 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.865 $Y=0
+ $X2=5.29 $Y2=0
r127 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=0 $X2=4.78
+ $Y2=0
r128 50 65 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.53
+ $Y2=0
r129 50 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.775
+ $Y2=0
r130 49 69 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.965 $Y=0
+ $X2=3.45 $Y2=0
r131 49 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.775
+ $Y2=0
r132 47 62 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.61
+ $Y2=0
r133 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.78
+ $Y2=0
r134 46 65 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.945 $Y=0
+ $X2=2.53 $Y2=0
r135 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.78
+ $Y2=0
r136 44 58 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.69
+ $Y2=0
r137 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.79
+ $Y2=0
r138 43 62 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=1.61 $Y2=0
r139 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.79
+ $Y2=0
r140 39 83 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=5.72 $Y=0.085
+ $X2=5.807 $Y2=0
r141 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.72 $Y=0.085
+ $X2=5.72 $Y2=0.39
r142 35 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=0.085
+ $X2=4.78 $Y2=0
r143 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.78 $Y=0.085
+ $X2=4.78 $Y2=0.39
r144 31 80 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0
r145 31 33 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0.4
r146 27 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=0.085
+ $X2=2.775 $Y2=0
r147 27 29 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.775 $Y=0.085
+ $X2=2.775 $Y2=0.4
r148 23 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r149 23 25 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.395
r150 19 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r151 19 21 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.66
r152 6 41 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.39
r153 5 37 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.595
+ $Y=0.235 $X2=4.78 $Y2=0.39
r154 4 33 182 $w=1.7e-07 $l=3.47851e-07 $layer=licon1_NDIFF $count=1 $X=3.555
+ $Y=0.235 $X2=3.83 $Y2=0.4
r155 3 29 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.4
r156 2 25 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.235 $X2=1.78 $Y2=0.395
r157 1 21 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.465 $X2=0.79 $Y2=0.66
.ends

