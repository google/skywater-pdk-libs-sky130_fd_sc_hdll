* File: sky130_fd_sc_hdll__a22oi_1.spice
* Created: Wed Sep  2 08:18:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a22oi_1.pex.spice"
.subckt sky130_fd_sc_hdll__a22oi_1  VNB VPB B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1007 A_119_47# N_B2_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.2015 PD=0.92 PS=1.92 NRD=14.76 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g A_119_47# VNB NSHORT L=0.15 W=0.65 AD=0.1755
+ AS=0.08775 PD=1.84 PS=0.92 NRD=0.912 NRS=14.76 M=1 R=4.33333 SA=75000.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 A_411_47# N_A1_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.2015 PD=0.92 PS=1.92 NRD=14.76 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g A_411_47# VNB NSHORT L=0.15 W=0.65 AD=0.2275
+ AS=0.08775 PD=2 PS=0.92 NRD=10.152 NRS=14.76 M=1 R=4.33333 SA=75000.7
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1002 N_A_117_297#_M1002_d N_B2_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_A_117_297#_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_117_297#_M1005_d N_A1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_117_297#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.31 AS=0.145 PD=2.62 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.778 P=10.41
pX9_noxref noxref_13 B1 B1 PROBETYPE=1
pX10_noxref noxref_14 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a22oi_1.pxi.spice"
*
.ends
*
*
