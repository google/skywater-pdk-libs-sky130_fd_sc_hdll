* File: sky130_fd_sc_hdll__inv_2.pxi.spice
* Created: Thu Aug 27 19:09:18 2020
* 
x_PM_SKY130_FD_SC_HDLL__INV_2%A N_A_c_30_n N_A_M1000_g N_A_c_26_n N_A_M1001_g
+ N_A_c_31_n N_A_M1003_g N_A_c_27_n N_A_M1002_g A N_A_c_29_n
+ PM_SKY130_FD_SC_HDLL__INV_2%A
x_PM_SKY130_FD_SC_HDLL__INV_2%VPWR N_VPWR_M1000_s N_VPWR_M1003_s N_VPWR_c_62_n
+ N_VPWR_c_63_n N_VPWR_c_64_n N_VPWR_c_65_n VPWR N_VPWR_c_66_n N_VPWR_c_61_n
+ N_VPWR_c_68_n PM_SKY130_FD_SC_HDLL__INV_2%VPWR
x_PM_SKY130_FD_SC_HDLL__INV_2%Y N_Y_M1001_s N_Y_M1000_d N_Y_c_85_n N_Y_c_86_n Y
+ Y Y Y Y PM_SKY130_FD_SC_HDLL__INV_2%Y
x_PM_SKY130_FD_SC_HDLL__INV_2%VGND N_VGND_M1001_d N_VGND_M1002_d N_VGND_c_107_n
+ N_VGND_c_108_n N_VGND_c_109_n N_VGND_c_110_n VGND N_VGND_c_111_n
+ N_VGND_c_112_n N_VGND_c_113_n PM_SKY130_FD_SC_HDLL__INV_2%VGND
cc_1 VNB N_A_c_26_n 0.0218806f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.995
cc_2 VNB N_A_c_27_n 0.0219019f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.995
cc_3 VNB A 0.00854082f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_c_29_n 0.0757777f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.202
cc_5 VNB N_VPWR_c_61_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB Y 0.00198623f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.202
cc_7 VNB N_VGND_c_107_n 0.010609f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_8 VNB N_VGND_c_108_n 0.0308509f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_9 VNB N_VGND_c_109_n 0.0207407f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.56
cc_10 VNB N_VGND_c_110_n 0.00930828f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.202
cc_11 VNB N_VGND_c_111_n 0.0182134f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.202
cc_12 VNB N_VGND_c_112_n 0.140956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_113_n 0.0040393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VPB N_A_c_30_n 0.0210369f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.41
cc_15 VPB N_A_c_31_n 0.0207627f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_16 VPB A 7.08627e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_17 VPB N_A_c_29_n 0.0365523f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.202
cc_18 VPB N_VPWR_c_62_n 0.0105831f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_19 VPB N_VPWR_c_63_n 0.0410274f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_20 VPB N_VPWR_c_64_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_21 VPB N_VPWR_c_65_n 0.00496839f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_22 VPB N_VPWR_c_66_n 0.0182134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_23 VPB N_VPWR_c_61_n 0.0609911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_68_n 0.00401341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB Y 0.00153746f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.202
cc_26 N_A_c_30_n N_VPWR_c_63_n 0.00766668f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_27 A N_VPWR_c_63_n 0.0185036f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_28 N_A_c_29_n N_VPWR_c_63_n 0.00531141f $X=0.975 $Y=1.202 $X2=0 $Y2=0
cc_29 N_A_c_30_n N_VPWR_c_64_n 0.00597712f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_30 N_A_c_31_n N_VPWR_c_64_n 0.00673617f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_31 N_A_c_31_n N_VPWR_c_65_n 0.00831232f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_32 N_A_c_30_n N_VPWR_c_61_n 0.0109152f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_33 N_A_c_31_n N_VPWR_c_61_n 0.0131262f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_34 N_A_c_26_n N_Y_c_85_n 0.00695889f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_35 N_A_c_30_n N_Y_c_86_n 0.0120229f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_36 N_A_c_31_n N_Y_c_86_n 0.00989133f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_37 N_A_c_30_n Y 0.00210513f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_38 N_A_c_26_n Y 0.00759593f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_39 N_A_c_31_n Y 0.00388655f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_40 N_A_c_27_n Y 0.00273168f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_41 A Y 0.0185726f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_42 N_A_c_29_n Y 0.0473428f $X=0.975 $Y=1.202 $X2=0 $Y2=0
cc_43 N_A_c_30_n Y 0.0049031f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_44 N_A_c_31_n Y 0.00266144f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_45 N_A_c_26_n N_VGND_c_108_n 0.00659294f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_46 A N_VGND_c_108_n 0.0188678f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_47 N_A_c_29_n N_VGND_c_108_n 0.00585411f $X=0.975 $Y=1.202 $X2=0 $Y2=0
cc_48 N_A_c_26_n N_VGND_c_109_n 0.00465454f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_49 N_A_c_27_n N_VGND_c_109_n 0.00585385f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_50 N_A_c_27_n N_VGND_c_110_n 0.00490145f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_51 N_A_c_26_n N_VGND_c_112_n 0.00890904f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_52 N_A_c_27_n N_VGND_c_112_n 0.0119902f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_53 N_VPWR_c_61_n N_Y_M1000_d 0.00231261f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_54 N_VPWR_c_64_n N_Y_c_86_n 0.0223557f $X=1.125 $Y=2.72 $X2=0 $Y2=0
cc_55 N_VPWR_c_61_n N_Y_c_86_n 0.0140101f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_56 N_VPWR_c_63_n Y 0.0740092f $X=0.27 $Y=1.66 $X2=0 $Y2=0
cc_57 N_VPWR_c_65_n Y 0.0602777f $X=1.21 $Y=1.66 $X2=0 $Y2=0
cc_58 N_VPWR_c_65_n N_VGND_c_110_n 0.00776079f $X=1.21 $Y=1.66 $X2=0 $Y2=0
cc_59 N_Y_c_85_n N_VGND_c_108_n 0.0480547f $X=0.74 $Y=0.38 $X2=0 $Y2=0
cc_60 Y N_VGND_c_108_n 0.00119665f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_61 N_Y_c_85_n N_VGND_c_109_n 0.0231099f $X=0.74 $Y=0.38 $X2=0 $Y2=0
cc_62 Y N_VGND_c_110_n 0.00126619f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_63 N_Y_M1001_s N_VGND_c_112_n 0.00324782f $X=0.605 $Y=0.235 $X2=0 $Y2=0
cc_64 N_Y_c_85_n N_VGND_c_112_n 0.0141178f $X=0.74 $Y=0.38 $X2=0 $Y2=0
