* File: sky130_fd_sc_hdll__a32oi_4.spice
* Created: Wed Sep  2 08:21:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a32oi_4.pex.spice"
.subckt sky130_fd_sc_hdll__a32oi_4  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1002 N_A_27_47#_M1002_d N_B2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1024 N_A_27_47#_M1024_d N_B2_M1024_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1025 N_A_27_47#_M1024_d N_B2_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1039 N_A_27_47#_M1039_d N_B2_M1039_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1010 N_A_27_47#_M1039_d N_B1_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1017 N_A_27_47#_M1017_d N_B1_M1017_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1030 N_A_27_47#_M1017_d N_B1_M1030_g N_Y_M1030_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1033 N_A_27_47#_M1033_d N_B1_M1033_g N_Y_M1030_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_893_47#_M1007_d N_A1_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1013 N_A_893_47#_M1013_d N_A1_M1013_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1031 N_A_893_47#_M1013_d N_A1_M1031_g N_Y_M1031_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1034 N_A_893_47#_M1034_d N_A1_M1034_g N_Y_M1031_s VNB NSHORT L=0.15 W=0.65
+ AD=0.13325 AS=0.104 PD=1.06 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_893_47#_M1034_d N_A2_M1003_g N_A_1379_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.13325 AS=0.104 PD=1.06 PS=0.97 NRD=24.912 NRS=8.304 M=1 R=4.33333
+ SA=75002.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1018 N_A_893_47#_M1018_d N_A2_M1018_g N_A_1379_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1020 N_A_893_47#_M1018_d N_A2_M1020_g N_A_1379_47#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1036 N_A_893_47#_M1036_d N_A2_M1036_g N_A_1379_47#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1015 N_A_1379_47#_M1015_d N_A3_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1022 N_A_1379_47#_M1015_d N_A3_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1037 N_A_1379_47#_M1037_d N_A3_M1037_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1038 N_A_1379_47#_M1037_d N_A3_M1038_g N_VGND_M1038_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.182 PD=1.02 PS=1.86 NRD=8.304 NRS=0.912 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_297#_M1001_d N_B2_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90010.3 A=0.18 P=2.36 MULT=1
MM1012 N_A_27_297#_M1012_d N_B2_M1012_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90009.9 A=0.18 P=2.36 MULT=1
MM1021 N_A_27_297#_M1012_d N_B2_M1021_g N_Y_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90009.4 A=0.18 P=2.36 MULT=1
MM1035 N_A_27_297#_M1035_d N_B2_M1035_g N_Y_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90008.9 A=0.18 P=2.36 MULT=1
MM1000 N_A_27_297#_M1035_d N_B1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90008.5 A=0.18 P=2.36 MULT=1
MM1004 N_A_27_297#_M1004_d N_B1_M1004_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90008 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1004_d N_B1_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90007.5 A=0.18 P=2.36 MULT=1
MM1016 N_A_27_297#_M1016_d N_B1_M1016_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.155 AS=0.145 PD=1.31 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90007 A=0.18 P=2.36 MULT=1
MM1005 N_A_27_297#_M1016_d N_A1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.155 AS=0.145 PD=1.31 PS=1.29 NRD=4.9053 NRS=0.9653 M=1 R=5.55556 SA=90004
+ SB=90006.6 A=0.18 P=2.36 MULT=1
MM1011 N_A_27_297#_M1011_d N_A1_M1011_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90006.1 A=0.18 P=2.36 MULT=1
MM1026 N_A_27_297#_M1011_d N_A1_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.3725 PD=1.29 PS=1.745 NRD=0.9653 NRS=7.8603 M=1 R=5.55556
+ SA=90004.9 SB=90005.6 A=0.18 P=2.36 MULT=1
MM1029 N_A_27_297#_M1029_d N_A1_M1029_g N_VPWR_M1026_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2625 AS=0.3725 PD=1.525 PS=1.745 NRD=0.9653 NRS=16.7253 M=1 R=5.55556
+ SA=90005.8 SB=90004.7 A=0.18 P=2.36 MULT=1
MM1008 N_A_27_297#_M1029_d N_A2_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2625 AS=0.145 PD=1.525 PS=1.29 NRD=47.2603 NRS=0.9653 M=1 R=5.55556
+ SA=90006.5 SB=90004 A=0.18 P=2.36 MULT=1
MM1014 N_A_27_297#_M1014_d N_A2_M1014_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90007
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1019 N_A_27_297#_M1014_d N_A2_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.5 SB=90003 A=0.18 P=2.36 MULT=1
MM1027 N_A_27_297#_M1027_d N_A2_M1027_g N_VPWR_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.405 AS=0.145 PD=1.81 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.9 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A3_M1006_g N_A_27_297#_M1027_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.405 PD=1.29 PS=1.81 NRD=0.9653 NRS=103.405 M=1 R=5.55556
+ SA=90008.9 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1006_d N_A3_M1023_g N_A_27_297#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90009.4 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1028 N_VPWR_M1028_d N_A3_M1028_g N_A_27_297#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90009.9 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1032 N_VPWR_M1028_d N_A3_M1032_g N_A_27_297#_M1032_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90010.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.0674 P=26.97
pX41_noxref noxref_15 Y Y PROBETYPE=1
pX42_noxref noxref_16 Y Y PROBETYPE=1
pX43_noxref noxref_17 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a32oi_4.pxi.spice"
*
.ends
*
*
