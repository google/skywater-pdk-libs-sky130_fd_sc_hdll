* File: sky130_fd_sc_hdll__o221ai_1.pex.spice
* Created: Thu Aug 27 19:20:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%C1 1 3 4 6 7 11
r25 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.38
+ $Y=1.16 $X2=0.38 $Y2=1.16
r26 7 11 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.23 $Y=1.16 $X2=0.38
+ $Y2=1.16
r27 4 10 38.6365 $w=3.35e-07 $l=2.13014e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.43 $Y2=1.16
r28 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r29 1 10 46.2237 $w=3.35e-07 $l=2.89396e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.43 $Y2=1.16
r30 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%B1 1 3 4 6 7 11 13
r25 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.51
+ $Y=1.16 $X2=1.51 $Y2=1.16
r26 7 11 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=1.51 $Y2=1.16
r27 7 13 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.155 $Y=1.16 $X2=1.15
+ $Y2=1.16
r28 4 10 38.7956 $w=3.51e-07 $l=2.16852e-07 $layer=POLY_cond $X=1.69 $Y=0.995
+ $X2=1.57 $Y2=1.16
r29 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.69 $Y=0.995 $X2=1.69
+ $Y2=0.56
r30 1 10 45.736 $w=3.51e-07 $l=2.93684e-07 $layer=POLY_cond $X=1.665 $Y=1.41
+ $X2=1.57 $Y2=1.16
r31 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.665 $Y=1.41
+ $X2=1.665 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%B2 1 3 4 6 7 13
r34 7 13 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.08 $Y=1.16 $X2=1.98
+ $Y2=1.16
r35 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.16 $X2=2.14 $Y2=1.16
r36 4 10 38.578 $w=2.95e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.16 $Y=0.995
+ $X2=2.165 $Y2=1.16
r37 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.16 $Y=0.995 $X2=2.16
+ $Y2=0.56
r38 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.165 $Y2=1.16
r39 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.105 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%A2 1 3 4 6 8 10 17 19
r46 17 19 11.5222 $w=2.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.99 $Y=1.615
+ $X2=2.99 $Y2=1.87
r47 10 13 3.79523 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=1.16 $X2=2.7
+ $Y2=1.245
r48 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.16 $X2=2.67 $Y2=1.16
r49 8 17 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.765 $Y=1.53
+ $X2=2.99 $Y2=1.53
r50 8 13 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=2.765 $Y=1.445
+ $X2=2.765 $Y2=1.245
r51 4 11 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.755 $Y=1.41
+ $X2=2.695 $Y2=1.16
r52 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.755 $Y=1.41
+ $X2=2.755 $Y2=1.985
r53 1 11 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=2.72 $Y=0.995
+ $X2=2.695 $Y2=1.16
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.72 $Y=0.995 $X2=2.72
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%A1 1 3 4 6 7 14
r24 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.375
+ $Y=1.16 $X2=3.375 $Y2=1.16
r25 7 14 3.05 $w=1.98e-07 $l=5.5e-08 $layer=LI1_cond $X=3.43 $Y=1.175 $X2=3.375
+ $Y2=1.175
r26 4 10 44.7611 $w=4.18e-07 $l=3.11047e-07 $layer=POLY_cond $X=3.165 $Y=1.41
+ $X2=3.302 $Y2=1.16
r27 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.165 $Y=1.41
+ $X2=3.165 $Y2=1.985
r28 1 10 39.9551 $w=4.18e-07 $l=2.32282e-07 $layer=POLY_cond $X=3.14 $Y=0.995
+ $X2=3.302 $Y2=1.16
r29 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.14 $Y=0.995 $X2=3.14
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%Y 1 2 3 10 13 15 17 18 19 22 23 27 28 31
+ 32 41
r63 41 42 0.662163 $w=6.03e-07 $l=3e-08 $layer=LI1_cond $X=2.202 $Y=2.21
+ $X2=2.202 $Y2=2.18
r64 32 45 2.0363 $w=6.03e-07 $l=1.03e-07 $layer=LI1_cond $X=2.202 $Y=2.237
+ $X2=2.202 $Y2=2.34
r65 32 41 0.533787 $w=6.03e-07 $l=2.7e-08 $layer=LI1_cond $X=2.202 $Y=2.237
+ $X2=2.202 $Y2=2.21
r66 32 42 0.592747 $w=5.63e-07 $l=2.8e-08 $layer=LI1_cond $X=2.182 $Y=2.152
+ $X2=2.182 $Y2=2.18
r67 31 32 5.96981 $w=5.63e-07 $l=2.82e-07 $layer=LI1_cond $X=2.182 $Y=1.87
+ $X2=2.182 $Y2=2.152
r68 28 31 3.49297 $w=5.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.182 $Y=1.705
+ $X2=2.182 $Y2=1.87
r69 28 30 2.40612 $w=5.65e-07 $l=1.05e-07 $layer=LI1_cond $X=2.182 $Y=1.705
+ $X2=2.182 $Y2=1.6
r70 24 27 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=1.6 $X2=0.76
+ $Y2=1.6
r71 23 30 6.46215 $w=2.1e-07 $l=2.82e-07 $layer=LI1_cond $X=1.9 $Y=1.6 $X2=2.182
+ $Y2=1.6
r72 23 24 55.7186 $w=2.08e-07 $l=1.055e-06 $layer=LI1_cond $X=1.9 $Y=1.6
+ $X2=0.845 $Y2=1.6
r73 22 27 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.76 $Y=1.495
+ $X2=0.76 $Y2=1.6
r74 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.76 $Y=0.825
+ $X2=0.76 $Y2=1.495
r75 20 26 3.99943 $w=2.1e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=1.6
+ $X2=0.225 $Y2=1.6
r76 19 27 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=1.6 $X2=0.76
+ $Y2=1.6
r77 19 20 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=0.675 $Y=1.6
+ $X2=0.365 $Y2=1.6
r78 17 21 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.675 $Y=0.735
+ $X2=0.76 $Y2=0.825
r79 17 18 20.3333 $w=1.78e-07 $l=3.3e-07 $layer=LI1_cond $X=0.675 $Y=0.735
+ $X2=0.345 $Y2=0.735
r80 13 26 2.99957 $w=2.8e-07 $l=1.05e-07 $layer=LI1_cond $X=0.225 $Y=1.705
+ $X2=0.225 $Y2=1.6
r81 13 15 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.225 $Y=1.705
+ $X2=0.225 $Y2=1.96
r82 10 18 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=0.215 $Y=0.645
+ $X2=0.345 $Y2=0.735
r83 10 12 2.34615 $w=2.6e-07 $l=5e-08 $layer=LI1_cond $X=0.215 $Y=0.645
+ $X2=0.215 $Y2=0.595
r84 3 45 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.195
+ $Y=1.485 $X2=2.34 $Y2=2.34
r85 3 30 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=2.195
+ $Y=1.485 $X2=2.34 $Y2=1.66
r86 2 26 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r87 2 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.96
r88 1 12 182 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%VPWR 1 2 7 9 13 20 31 34 37
r43 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 33 34 12.4498 $w=9.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=2.34
+ $X2=1.58 $Y2=2.34
r45 29 33 3.47634 $w=9.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.15 $Y=2.34
+ $X2=1.415 $Y2=2.34
r46 29 31 17.5003 $w=9.28e-07 $l=5.5e-07 $layer=LI1_cond $X=1.15 $Y=2.34 $X2=0.6
+ $Y2=2.34
r47 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r49 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 24 27 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 23 26 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 23 34 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.61 $Y=2.72 $X2=1.58
+ $Y2=2.72
r54 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 20 36 4.11481 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.315 $Y=2.72
+ $X2=3.497 $Y2=2.72
r56 20 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.315 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 17 31 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=0.6
+ $Y2=2.72
r58 13 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 13 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r60 9 12 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=3.445 $Y=1.66
+ $X2=3.445 $Y2=2.34
r61 7 36 3.09741 $w=2.6e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.445 $Y=2.635
+ $X2=3.497 $Y2=2.72
r62 7 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.445 $Y=2.635
+ $X2=3.445 $Y2=2.34
r63 2 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=1.485 $X2=3.4 $Y2=2.34
r64 2 9 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=1.485 $X2=3.4 $Y2=1.66
r65 1 33 150 $w=1.7e-07 $l=1.02022e-06 $layer=licon1_PDIFF $count=4 $X=0.605
+ $Y=1.485 $X2=1.415 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%A_123_47# 1 2 11
r15 8 11 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=0.75 $Y=0.39 $X2=1.9
+ $Y2=0.39
r16 2 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.235 $X2=1.9 $Y2=0.39
r17 1 8 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%A_261_47# 1 2 3 10 16 20 23
r45 18 20 9.0127 $w=3.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.38 $Y=0.695
+ $X2=3.38 $Y2=0.39
r46 17 23 7.38875 $w=1.75e-07 $l=3.35783e-07 $layer=LI1_cond $X=2.56 $Y=0.78
+ $X2=2.285 $Y2=0.645
r47 16 18 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=3.185 $Y=0.78
+ $X2=3.38 $Y2=0.695
r48 16 17 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.185 $Y=0.78
+ $X2=2.56 $Y2=0.78
r49 10 23 7.38875 $w=1.75e-07 $l=9e-08 $layer=LI1_cond $X=2.285 $Y=0.735
+ $X2=2.285 $Y2=0.645
r50 10 12 52.6818 $w=1.78e-07 $l=8.55e-07 $layer=LI1_cond $X=2.285 $Y=0.735
+ $X2=1.43 $Y2=0.735
r51 3 20 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.215
+ $Y=0.235 $X2=3.4 $Y2=0.39
r52 2 23 182 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.235 $X2=2.37 $Y2=0.66
r53 1 12 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=1.305
+ $Y=0.235 $X2=1.43 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_1%VGND 1 6 9 10 11 21 22
r40 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r41 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r42 18 19 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r43 14 18 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r44 11 19 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r45 11 14 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r46 9 18 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.53
+ $Y2=0
r47 9 10 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.93
+ $Y2=0
r48 8 21 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.45
+ $Y2=0
r49 8 10 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=2.93
+ $Y2=0
r50 4 10 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=0.085 $X2=2.93
+ $Y2=0
r51 4 6 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.93 $Y=0.085
+ $X2=2.93 $Y2=0.36
r52 1 6 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.235 $X2=2.93 $Y2=0.36
.ends

