* File: sky130_fd_sc_hdll__a2bb2o_4.pxi.spice
* Created: Wed Sep  2 08:19:25 2020
* 
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%B1 N_B1_c_126_n N_B1_M1009_g N_B1_c_127_n
+ N_B1_M1018_g N_B1_c_128_n N_B1_M1015_g N_B1_c_129_n N_B1_M1019_g N_B1_c_135_n
+ N_B1_c_130_n N_B1_c_131_n B1 N_B1_c_132_n PM_SKY130_FD_SC_HDLL__A2BB2O_4%B1
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%B2 N_B2_c_208_n N_B2_M1006_g N_B2_c_212_n
+ N_B2_M1001_g N_B2_c_213_n N_B2_M1023_g N_B2_c_209_n N_B2_M1027_g B2
+ N_B2_c_210_n B2 PM_SKY130_FD_SC_HDLL__A2BB2O_4%B2
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_455_21# N_A_455_21#_M1000_d
+ N_A_455_21#_M1025_d N_A_455_21#_M1013_s N_A_455_21#_c_254_n
+ N_A_455_21#_M1014_g N_A_455_21#_c_265_n N_A_455_21#_M1005_g
+ N_A_455_21#_c_266_n N_A_455_21#_M1011_g N_A_455_21#_c_255_n
+ N_A_455_21#_M1022_g N_A_455_21#_c_256_n N_A_455_21#_c_257_n
+ N_A_455_21#_c_258_n N_A_455_21#_c_259_n N_A_455_21#_c_260_n
+ N_A_455_21#_c_277_p N_A_455_21#_c_283_p N_A_455_21#_c_261_n
+ N_A_455_21#_c_300_p N_A_455_21#_c_262_n N_A_455_21#_c_263_n
+ N_A_455_21#_c_291_p N_A_455_21#_c_264_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_455_21#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%A1_N N_A1_N_c_391_n N_A1_N_M1004_g
+ N_A1_N_c_392_n N_A1_N_M1000_g N_A1_N_c_393_n N_A1_N_M1026_g N_A1_N_c_394_n
+ N_A1_N_M1010_g N_A1_N_c_399_n N_A1_N_c_395_n A1_N
+ PM_SKY130_FD_SC_HDLL__A2BB2O_4%A1_N
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%A2_N N_A2_N_c_477_n N_A2_N_M1017_g
+ N_A2_N_c_481_n N_A2_N_M1013_g N_A2_N_c_482_n N_A2_N_M1020_g N_A2_N_c_478_n
+ N_A2_N_M1025_g A2_N N_A2_N_c_479_n N_A2_N_c_480_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_4%A2_N
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_203_47# N_A_203_47#_M1006_d
+ N_A_203_47#_M1014_s N_A_203_47#_M1005_s N_A_203_47#_c_526_n
+ N_A_203_47#_M1002_g N_A_203_47#_c_535_n N_A_203_47#_M1003_g
+ N_A_203_47#_c_527_n N_A_203_47#_M1007_g N_A_203_47#_c_536_n
+ N_A_203_47#_M1012_g N_A_203_47#_c_528_n N_A_203_47#_M1008_g
+ N_A_203_47#_c_537_n N_A_203_47#_M1016_g N_A_203_47#_c_538_n
+ N_A_203_47#_M1024_g N_A_203_47#_c_529_n N_A_203_47#_M1021_g
+ N_A_203_47#_c_530_n N_A_203_47#_c_549_n N_A_203_47#_c_531_n
+ N_A_203_47#_c_636_p N_A_203_47#_c_532_n N_A_203_47#_c_533_n
+ N_A_203_47#_c_540_n N_A_203_47#_c_541_n N_A_203_47#_c_596_n
+ N_A_203_47#_c_534_n N_A_203_47#_c_543_n N_A_203_47#_c_544_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_203_47#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_27_297# N_A_27_297#_M1009_s
+ N_A_27_297#_M1001_d N_A_27_297#_M1015_s N_A_27_297#_M1011_d
+ N_A_27_297#_c_736_p N_A_27_297#_c_699_n N_A_27_297#_c_695_n
+ N_A_27_297#_c_730_p N_A_27_297#_c_704_n N_A_27_297#_c_696_n
+ N_A_27_297#_c_716_n N_A_27_297#_c_734_p N_A_27_297#_c_710_n
+ N_A_27_297#_c_711_n N_A_27_297#_c_725_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%VPWR N_VPWR_M1009_d N_VPWR_M1023_s
+ N_VPWR_M1004_d N_VPWR_M1026_d N_VPWR_M1012_s N_VPWR_M1024_s N_VPWR_c_749_n
+ N_VPWR_c_750_n N_VPWR_c_751_n N_VPWR_c_752_n N_VPWR_c_753_n N_VPWR_c_754_n
+ N_VPWR_c_755_n N_VPWR_c_756_n N_VPWR_c_757_n N_VPWR_c_758_n N_VPWR_c_759_n
+ N_VPWR_c_760_n N_VPWR_c_761_n N_VPWR_c_762_n N_VPWR_c_763_n VPWR
+ N_VPWR_c_764_n N_VPWR_c_765_n N_VPWR_c_748_n N_VPWR_c_767_n N_VPWR_c_768_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_785_297# N_A_785_297#_M1004_s
+ N_A_785_297#_M1020_d N_A_785_297#_c_867_n N_A_785_297#_c_874_n
+ N_A_785_297#_c_870_n PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_785_297#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%X N_X_M1002_d N_X_M1008_d N_X_M1003_d
+ N_X_M1016_d N_X_c_897_n N_X_c_936_n N_X_c_900_n N_X_c_904_n N_X_c_885_n
+ N_X_c_886_n N_X_c_918_n N_X_c_941_n N_X_c_890_n N_X_c_887_n N_X_c_888_n
+ N_X_c_891_n X X N_X_c_893_n PM_SKY130_FD_SC_HDLL__A2BB2O_4%X
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%VGND N_VGND_M1018_s N_VGND_M1019_s
+ N_VGND_M1022_d N_VGND_M1017_s N_VGND_M1010_s N_VGND_M1007_s N_VGND_M1021_s
+ N_VGND_c_965_n N_VGND_c_966_n N_VGND_c_967_n N_VGND_c_968_n N_VGND_c_969_n
+ N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n N_VGND_c_974_n
+ N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n N_VGND_c_978_n N_VGND_c_979_n
+ VGND N_VGND_c_980_n N_VGND_c_981_n N_VGND_c_982_n N_VGND_c_983_n
+ N_VGND_c_984_n N_VGND_c_985_n PM_SKY130_FD_SC_HDLL__A2BB2O_4%VGND
x_PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_119_47# N_A_119_47#_M1018_d
+ N_A_119_47#_M1027_s N_A_119_47#_c_1091_n N_A_119_47#_c_1090_n
+ N_A_119_47#_c_1095_n PM_SKY130_FD_SC_HDLL__A2BB2O_4%A_119_47#
cc_1 VNB N_B1_c_126_n 0.0326155f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_B1_c_127_n 0.0218318f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_B1_c_128_n 0.022322f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_4 VNB N_B1_c_129_n 0.0166635f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_B1_c_130_n 7.01377e-19 $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.445
cc_6 VNB N_B1_c_131_n 0.00400122f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_7 VNB N_B1_c_132_n 0.015702f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_8 VNB N_B2_c_208_n 0.0170472f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_B2_c_209_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_10 VNB N_B2_c_210_n 0.0364409f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_11 VNB B2 0.00165109f $X=-0.19 $Y=-0.24 $X2=0.435 $Y2=1.16
cc_12 VNB N_A_455_21#_c_254_n 0.0168842f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_13 VNB N_A_455_21#_c_255_n 0.0203913f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_14 VNB N_A_455_21#_c_256_n 2.36777e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_455_21#_c_257_n 0.00342205f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_16 VNB N_A_455_21#_c_258_n 8.98821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_455_21#_c_259_n 0.00316518f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.19
cc_18 VNB N_A_455_21#_c_260_n 2.73823e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_455_21#_c_261_n 0.00603069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_455_21#_c_262_n 0.00108975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_455_21#_c_263_n 0.00323152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_455_21#_c_264_n 0.0583828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A1_N_c_391_n 0.0272393f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_24 VNB N_A1_N_c_392_n 0.0196954f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_25 VNB N_A1_N_c_393_n 0.0254053f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_26 VNB N_A1_N_c_394_n 0.0169367f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_27 VNB N_A1_N_c_395_n 0.00325404f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.445
cc_28 VNB A1_N 0.00194469f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_29 VNB N_A2_N_c_477_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_30 VNB N_A2_N_c_478_n 0.0173889f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_31 VNB N_A2_N_c_479_n 0.00318801f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_32 VNB N_A2_N_c_480_n 0.0343033f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_33 VNB N_A_203_47#_c_526_n 0.016627f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_34 VNB N_A_203_47#_c_527_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.445
cc_35 VNB N_A_203_47#_c_528_n 0.0171989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_203_47#_c_529_n 0.0200861f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.19
cc_37 VNB N_A_203_47#_c_530_n 0.00707111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_203_47#_c_531_n 0.00163384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_203_47#_c_532_n 0.00266295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_203_47#_c_533_n 0.00344627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_203_47#_c_534_n 0.0769623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_748_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_X_c_885_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_44 VNB N_X_c_886_n 0.00240962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_X_c_887_n 0.0127057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_X_c_888_n 0.00261326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB X 0.0229789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_965_n 0.0110494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_966_n 0.00651836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_967_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_51 VNB N_VGND_c_968_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_969_n 0.00741231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_970_n 0.00468725f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_971_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_972_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_973_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_974_n 0.0201004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_975_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_976_n 0.0201935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_977_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_978_n 0.0195532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_979_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_980_n 0.0407345f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_981_n 0.0132245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_982_n 0.3766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_983_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_984_n 0.0201295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_985_n 0.0208882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_119_47#_c_1090_n 0.00331877f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_70 VPB N_B1_c_126_n 0.0301878f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_71 VPB N_B1_c_128_n 0.0257974f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_72 VPB N_B1_c_135_n 0.00820796f $X=-0.19 $Y=1.305 $X2=1.665 $Y2=1.53
cc_73 VPB N_B1_c_130_n 0.00130348f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.445
cc_74 VPB N_B1_c_132_n 0.0162013f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_75 VPB N_B2_c_212_n 0.0159799f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_76 VPB N_B2_c_213_n 0.0159754f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_77 VPB N_B2_c_210_n 0.0193472f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_78 VPB N_A_455_21#_c_265_n 0.0163347f $X=-0.19 $Y=1.305 $X2=1.665 $Y2=1.53
cc_79 VPB N_A_455_21#_c_266_n 0.019515f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.445
cc_80 VPB N_A_455_21#_c_258_n 0.0181321f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_455_21#_c_264_n 0.0333895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A1_N_c_391_n 0.0313923f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_83 VPB N_A1_N_c_393_n 0.0248459f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_84 VPB N_A1_N_c_399_n 0.0077654f $X=-0.19 $Y=1.305 $X2=1.665 $Y2=1.53
cc_85 VPB N_A1_N_c_395_n 0.00283438f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.445
cc_86 VPB A1_N 0.00232579f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_87 VPB N_A2_N_c_481_n 0.0159773f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_88 VPB N_A2_N_c_482_n 0.0159792f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_89 VPB N_A2_N_c_480_n 0.0192755f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_90 VPB N_A_203_47#_c_535_n 0.0159538f $X=-0.19 $Y=1.305 $X2=1.665 $Y2=1.53
cc_91 VPB N_A_203_47#_c_536_n 0.0160946f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_92 VPB N_A_203_47#_c_537_n 0.0160765f $X=-0.19 $Y=1.305 $X2=0.435 $Y2=1.16
cc_93 VPB N_A_203_47#_c_538_n 0.0191635f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.16
cc_94 VPB N_A_203_47#_c_531_n 0.00155612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_203_47#_c_540_n 0.00962913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_203_47#_c_541_n 0.00137626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_203_47#_c_534_n 0.0484324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_203_47#_c_543_n 0.00103996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_203_47#_c_544_n 0.00161355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_27_297#_c_695_n 0.00692367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_27_297#_c_696_n 0.00358759f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.19
cc_102 VPB N_VPWR_c_749_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_103 VPB N_VPWR_c_750_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_104 VPB N_VPWR_c_751_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_105 VPB N_VPWR_c_752_n 0.00518f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.19
cc_106 VPB N_VPWR_c_753_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_754_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_755_n 0.00518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_756_n 0.041786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_757_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_758_n 0.0395589f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_759_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_760_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_761_n 0.00478125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_762_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_763_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_764_n 0.0190625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_765_n 0.0128037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_748_n 0.0654928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_767_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_768_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_X_c_890_n 0.00140119f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.53
cc_123 VPB N_X_c_891_n 0.00245799f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB X 0.00629494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_X_c_893_n 0.0192751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 N_B1_c_127_n N_B2_c_208_n 0.0165098f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_127 N_B1_c_126_n N_B2_c_212_n 0.0371597f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B1_c_135_n N_B2_c_212_n 0.0114861f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_129 N_B1_c_132_n N_B2_c_212_n 9.80334e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B1_c_128_n N_B2_c_213_n 0.0364057f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_131 N_B1_c_135_n N_B2_c_213_n 0.0128234f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_132 N_B1_c_130_n N_B2_c_213_n 7.38573e-19 $X=1.75 $Y=1.445 $X2=0 $Y2=0
cc_133 N_B1_c_129_n N_B2_c_209_n 0.0224097f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B1_c_126_n N_B2_c_210_n 0.0165098f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_135 N_B1_c_128_n N_B2_c_210_n 0.0263437f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B1_c_135_n N_B2_c_210_n 0.00803891f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_137 N_B1_c_130_n N_B2_c_210_n 0.0031808f $X=1.75 $Y=1.445 $X2=0 $Y2=0
cc_138 N_B1_c_131_n N_B2_c_210_n 0.0012824f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_139 N_B1_c_132_n N_B2_c_210_n 0.00409926f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B1_c_126_n B2 7.71575e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B1_c_135_n B2 0.0416942f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_142 N_B1_c_130_n B2 0.00188538f $X=1.75 $Y=1.445 $X2=0 $Y2=0
cc_143 N_B1_c_131_n B2 0.0117655f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_144 N_B1_c_132_n B2 0.0145168f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_145 N_B1_c_129_n N_A_455_21#_c_254_n 0.0262119f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B1_c_128_n N_A_455_21#_c_265_n 0.0091518f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B1_c_128_n N_A_455_21#_c_264_n 0.026706f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B1_c_130_n N_A_455_21#_c_264_n 4.98708e-19 $X=1.75 $Y=1.445 $X2=0 $Y2=0
cc_149 N_B1_c_131_n N_A_455_21#_c_264_n 0.00154647f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_150 N_B1_c_128_n N_A_203_47#_c_530_n 0.00437379f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B1_c_129_n N_A_203_47#_c_530_n 0.0123512f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B1_c_135_n N_A_203_47#_c_530_n 0.00677802f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_153 N_B1_c_131_n N_A_203_47#_c_530_n 0.030608f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_154 N_B1_c_129_n N_A_203_47#_c_549_n 9.08954e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B1_c_128_n N_A_203_47#_c_531_n 7.5473e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_156 N_B1_c_130_n N_A_203_47#_c_531_n 0.00411607f $X=1.75 $Y=1.445 $X2=0 $Y2=0
cc_157 N_B1_c_131_n N_A_203_47#_c_531_n 0.00711829f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_158 N_B1_c_135_n N_A_203_47#_c_543_n 3.01707e-19 $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_159 N_B1_c_130_n N_A_203_47#_c_543_n 8.13951e-19 $X=1.75 $Y=1.445 $X2=0 $Y2=0
cc_160 N_B1_c_132_n N_A_27_297#_M1009_s 0.00284151f $X=0.41 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_161 N_B1_c_135_n N_A_27_297#_M1001_d 0.00187091f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_162 N_B1_c_126_n N_A_27_297#_c_699_n 0.0112216f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_163 N_B1_c_135_n N_A_27_297#_c_699_n 0.02495f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_164 N_B1_c_132_n N_A_27_297#_c_699_n 0.0134161f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B1_c_126_n N_A_27_297#_c_695_n 3.96914e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B1_c_132_n N_A_27_297#_c_695_n 0.0188817f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_167 N_B1_c_128_n N_A_27_297#_c_704_n 0.013306f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_168 N_B1_c_135_n N_A_27_297#_c_704_n 0.0267794f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_169 N_B1_c_131_n N_A_27_297#_c_704_n 0.00448404f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B1_c_128_n N_A_27_297#_c_696_n 0.00441059f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_171 N_B1_c_135_n N_A_27_297#_c_696_n 0.0104943f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_172 N_B1_c_131_n N_A_27_297#_c_696_n 0.00280327f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_173 N_B1_c_135_n N_A_27_297#_c_710_n 0.0143191f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_174 N_B1_c_128_n N_A_27_297#_c_711_n 6.11739e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B1_c_131_n N_A_27_297#_c_711_n 5.83252e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_176 N_B1_c_135_n N_VPWR_M1009_d 0.00187547f $X=1.665 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_177 N_B1_c_135_n N_VPWR_M1023_s 0.00187562f $X=1.665 $Y=1.53 $X2=0 $Y2=0
cc_178 N_B1_c_126_n N_VPWR_c_749_n 0.00300743f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B1_c_128_n N_VPWR_c_751_n 0.00300743f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B1_c_128_n N_VPWR_c_756_n 0.00702461f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_181 N_B1_c_126_n N_VPWR_c_764_n 0.00702461f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B1_c_126_n N_VPWR_c_748_n 0.00787122f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B1_c_128_n N_VPWR_c_748_n 0.006985f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_184 N_B1_c_126_n N_VGND_c_966_n 0.00176179f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B1_c_127_n N_VGND_c_966_n 0.00614111f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_132_n N_VGND_c_966_n 0.0145468f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_187 N_B1_c_129_n N_VGND_c_967_n 0.00268723f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B1_c_127_n N_VGND_c_980_n 0.00463936f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_129_n N_VGND_c_980_n 0.00439206f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B1_c_127_n N_VGND_c_982_n 0.00876414f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_191 N_B1_c_129_n N_VGND_c_982_n 0.00608392f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B1_c_127_n N_A_119_47#_c_1091_n 0.00382935f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_193 N_B1_c_127_n N_A_119_47#_c_1090_n 0.00778436f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_B1_c_135_n N_A_119_47#_c_1090_n 0.00711902f $X=1.665 $Y=1.53 $X2=0
+ $Y2=0
cc_195 N_B1_c_132_n N_A_119_47#_c_1090_n 0.00921104f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_196 N_B2_c_209_n N_A_203_47#_c_530_n 0.0102977f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_197 B2 N_A_203_47#_c_530_n 0.00520428f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_198 N_B2_c_208_n N_A_203_47#_c_532_n 0.00373848f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B2_c_210_n N_A_203_47#_c_532_n 0.00473714f $X=1.435 $Y=1.202 $X2=0
+ $Y2=0
cc_200 B2 N_A_203_47#_c_532_n 0.0287145f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_201 N_B2_c_212_n N_A_27_297#_c_699_n 0.011229f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B2_c_213_n N_A_27_297#_c_704_n 0.011229f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B2_c_212_n N_VPWR_c_749_n 0.00300743f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B2_c_212_n N_VPWR_c_750_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B2_c_213_n N_VPWR_c_750_n 0.00702461f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B2_c_213_n N_VPWR_c_751_n 0.00300743f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B2_c_212_n N_VPWR_c_748_n 0.00695979f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B2_c_213_n N_VPWR_c_748_n 0.00695979f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B2_c_208_n N_VGND_c_980_n 0.00357877f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B2_c_209_n N_VGND_c_980_n 0.00357877f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B2_c_208_n N_VGND_c_982_n 0.005504f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B2_c_209_n N_VGND_c_982_n 0.00562222f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B2_c_208_n N_A_119_47#_c_1095_n 0.0112999f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B2_c_209_n N_A_119_47#_c_1095_n 0.0101752f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_215 B2 N_A_119_47#_c_1095_n 0.00314553f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_216 N_A_455_21#_c_257_n N_A1_N_c_391_n 0.00182734f $X=3.35 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_217 N_A_455_21#_c_258_n N_A1_N_c_391_n 0.0116392f $X=3.35 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_218 N_A_455_21#_c_259_n N_A1_N_c_391_n 0.00437722f $X=3.855 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_219 N_A_455_21#_c_277_p N_A1_N_c_391_n 0.0167894f $X=4.415 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_220 N_A_455_21#_c_262_n N_A1_N_c_391_n 6.99754e-19 $X=3.35 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_221 N_A_455_21#_c_263_n N_A1_N_c_391_n 0.00153445f $X=4.045 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_222 N_A_455_21#_c_264_n N_A1_N_c_391_n 0.010045f $X=2.87 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_223 N_A_455_21#_c_257_n N_A1_N_c_392_n 0.00257611f $X=3.35 $Y=1.075 $X2=0
+ $Y2=0
cc_224 N_A_455_21#_c_259_n N_A1_N_c_392_n 0.00789941f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_225 N_A_455_21#_c_283_p N_A1_N_c_392_n 0.0131824f $X=4.07 $Y=0.39 $X2=0 $Y2=0
cc_226 N_A_455_21#_c_263_n N_A1_N_c_392_n 0.00269099f $X=4.045 $Y=0.815 $X2=0
+ $Y2=0
cc_227 N_A_455_21#_c_261_n N_A1_N_c_393_n 0.00242197f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_228 N_A_455_21#_c_261_n N_A1_N_c_394_n 2.64252e-19 $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_229 N_A_455_21#_M1013_s N_A1_N_c_399_n 0.00187091f $X=4.395 $Y=1.485 $X2=0
+ $Y2=0
cc_230 N_A_455_21#_c_277_p N_A1_N_c_399_n 0.0211921f $X=4.415 $Y=1.875 $X2=0
+ $Y2=0
cc_231 N_A_455_21#_c_261_n N_A1_N_c_399_n 0.00497692f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_232 N_A_455_21#_c_263_n N_A1_N_c_399_n 0.00583827f $X=4.045 $Y=0.815 $X2=0
+ $Y2=0
cc_233 N_A_455_21#_c_291_p N_A1_N_c_399_n 0.012249f $X=4.54 $Y=1.875 $X2=0 $Y2=0
cc_234 N_A_455_21#_c_258_n N_A1_N_c_395_n 0.0218716f $X=3.35 $Y=1.495 $X2=0
+ $Y2=0
cc_235 N_A_455_21#_c_259_n N_A1_N_c_395_n 0.0173881f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_236 N_A_455_21#_c_277_p N_A1_N_c_395_n 0.0139804f $X=4.415 $Y=1.875 $X2=0
+ $Y2=0
cc_237 N_A_455_21#_c_262_n N_A1_N_c_395_n 0.0143867f $X=3.35 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_455_21#_c_263_n N_A1_N_c_395_n 0.012421f $X=4.045 $Y=0.815 $X2=0
+ $Y2=0
cc_239 N_A_455_21#_c_261_n A1_N 0.00754391f $X=4.795 $Y=0.815 $X2=0 $Y2=0
cc_240 N_A_455_21#_c_283_p N_A2_N_c_477_n 0.00693563f $X=4.07 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_241 N_A_455_21#_c_261_n N_A2_N_c_477_n 0.00928566f $X=4.795 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_242 N_A_455_21#_c_300_p N_A2_N_c_477_n 5.69266e-19 $X=5.01 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_243 N_A_455_21#_c_263_n N_A2_N_c_477_n 0.00112628f $X=4.045 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_244 N_A_455_21#_c_277_p N_A2_N_c_481_n 0.0109979f $X=4.415 $Y=1.875 $X2=0
+ $Y2=0
cc_245 N_A_455_21#_c_283_p N_A2_N_c_478_n 5.34196e-19 $X=4.07 $Y=0.39 $X2=0
+ $Y2=0
cc_246 N_A_455_21#_c_261_n N_A2_N_c_478_n 0.00919116f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_247 N_A_455_21#_c_300_p N_A2_N_c_478_n 0.00857123f $X=5.01 $Y=0.39 $X2=0
+ $Y2=0
cc_248 N_A_455_21#_c_261_n N_A2_N_c_479_n 0.0479975f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_249 N_A_455_21#_c_263_n N_A2_N_c_479_n 0.00223111f $X=4.045 $Y=0.815 $X2=0
+ $Y2=0
cc_250 N_A_455_21#_c_261_n N_A2_N_c_480_n 0.00468948f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_251 N_A_455_21#_c_254_n N_A_203_47#_c_530_n 0.0120679f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A_455_21#_c_254_n N_A_203_47#_c_549_n 0.00671955f $X=2.35 $Y=0.995
+ $X2=0 $Y2=0
cc_253 N_A_455_21#_c_254_n N_A_203_47#_c_531_n 0.00229843f $X=2.35 $Y=0.995
+ $X2=0 $Y2=0
cc_254 N_A_455_21#_c_255_n N_A_203_47#_c_531_n 0.00109583f $X=2.87 $Y=0.995
+ $X2=0 $Y2=0
cc_255 N_A_455_21#_c_256_n N_A_203_47#_c_531_n 0.0128172f $X=3.255 $Y=1.16 $X2=0
+ $Y2=0
cc_256 N_A_455_21#_c_257_n N_A_203_47#_c_531_n 0.00533218f $X=3.35 $Y=1.075
+ $X2=0 $Y2=0
cc_257 N_A_455_21#_c_258_n N_A_203_47#_c_531_n 0.00534715f $X=3.35 $Y=1.495
+ $X2=0 $Y2=0
cc_258 N_A_455_21#_c_264_n N_A_203_47#_c_531_n 0.0297448f $X=2.87 $Y=1.202 $X2=0
+ $Y2=0
cc_259 N_A_455_21#_c_254_n N_A_203_47#_c_533_n 0.00221247f $X=2.35 $Y=0.995
+ $X2=0 $Y2=0
cc_260 N_A_455_21#_c_255_n N_A_203_47#_c_533_n 3.09077e-19 $X=2.87 $Y=0.995
+ $X2=0 $Y2=0
cc_261 N_A_455_21#_c_260_n N_A_203_47#_c_533_n 0.00399829f $X=3.445 $Y=0.815
+ $X2=0 $Y2=0
cc_262 N_A_455_21#_c_264_n N_A_203_47#_c_533_n 3.11942e-19 $X=2.87 $Y=1.202
+ $X2=0 $Y2=0
cc_263 N_A_455_21#_c_256_n N_A_203_47#_c_540_n 0.0109126f $X=3.255 $Y=1.16 $X2=0
+ $Y2=0
cc_264 N_A_455_21#_c_258_n N_A_203_47#_c_540_n 0.0326955f $X=3.35 $Y=1.495 $X2=0
+ $Y2=0
cc_265 N_A_455_21#_c_259_n N_A_203_47#_c_540_n 0.00403943f $X=3.855 $Y=0.815
+ $X2=0 $Y2=0
cc_266 N_A_455_21#_c_277_p N_A_203_47#_c_540_n 0.00955488f $X=4.415 $Y=1.875
+ $X2=0 $Y2=0
cc_267 N_A_455_21#_c_261_n N_A_203_47#_c_540_n 0.00186279f $X=4.795 $Y=0.815
+ $X2=0 $Y2=0
cc_268 N_A_455_21#_c_263_n N_A_203_47#_c_540_n 0.00214973f $X=4.045 $Y=0.815
+ $X2=0 $Y2=0
cc_269 N_A_455_21#_c_291_p N_A_203_47#_c_540_n 0.00196365f $X=4.54 $Y=1.875
+ $X2=0 $Y2=0
cc_270 N_A_455_21#_c_264_n N_A_203_47#_c_540_n 0.00651916f $X=2.87 $Y=1.202
+ $X2=0 $Y2=0
cc_271 N_A_455_21#_c_266_n N_A_203_47#_c_541_n 0.0106521f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_272 N_A_455_21#_c_256_n N_A_203_47#_c_541_n 0.00462025f $X=3.255 $Y=1.16
+ $X2=0 $Y2=0
cc_273 N_A_455_21#_c_258_n N_A_203_47#_c_541_n 0.00264115f $X=3.35 $Y=1.495
+ $X2=0 $Y2=0
cc_274 N_A_455_21#_c_264_n N_A_203_47#_c_541_n 0.00127578f $X=2.87 $Y=1.202
+ $X2=0 $Y2=0
cc_275 N_A_455_21#_c_265_n N_A_203_47#_c_543_n 9.19852e-19 $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_276 N_A_455_21#_c_266_n N_A_203_47#_c_543_n 0.0181805f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_277 N_A_455_21#_c_256_n N_A_203_47#_c_543_n 3.03251e-19 $X=3.255 $Y=1.16
+ $X2=0 $Y2=0
cc_278 N_A_455_21#_c_258_n N_A_203_47#_c_543_n 0.016959f $X=3.35 $Y=1.495 $X2=0
+ $Y2=0
cc_279 N_A_455_21#_c_264_n N_A_203_47#_c_543_n 0.00197656f $X=2.87 $Y=1.202
+ $X2=0 $Y2=0
cc_280 N_A_455_21#_c_265_n N_A_27_297#_c_696_n 2.60649e-19 $X=2.375 $Y=1.41
+ $X2=0 $Y2=0
cc_281 N_A_455_21#_c_265_n N_A_27_297#_c_716_n 0.0143148f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_282 N_A_455_21#_c_266_n N_A_27_297#_c_716_n 0.0115264f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_283 N_A_455_21#_c_258_n N_VPWR_M1004_d 0.00804979f $X=3.35 $Y=1.495 $X2=0
+ $Y2=0
cc_284 N_A_455_21#_c_277_p N_VPWR_M1004_d 0.00188124f $X=4.415 $Y=1.875 $X2=0
+ $Y2=0
cc_285 N_A_455_21#_c_266_n N_VPWR_c_752_n 0.00213395f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_286 N_A_455_21#_c_258_n N_VPWR_c_752_n 0.0105983f $X=3.35 $Y=1.495 $X2=0
+ $Y2=0
cc_287 N_A_455_21#_c_277_p N_VPWR_c_752_n 0.00630624f $X=4.415 $Y=1.875 $X2=0
+ $Y2=0
cc_288 N_A_455_21#_c_265_n N_VPWR_c_756_n 0.00429453f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_455_21#_c_266_n N_VPWR_c_756_n 0.00429453f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_290 N_A_455_21#_c_258_n N_VPWR_c_756_n 6.22982e-19 $X=3.35 $Y=1.495 $X2=0
+ $Y2=0
cc_291 N_A_455_21#_c_277_p N_VPWR_c_758_n 0.00256479f $X=4.415 $Y=1.875 $X2=0
+ $Y2=0
cc_292 N_A_455_21#_M1013_s N_VPWR_c_748_n 0.00232092f $X=4.395 $Y=1.485 $X2=0
+ $Y2=0
cc_293 N_A_455_21#_c_265_n N_VPWR_c_748_n 0.00609021f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_294 N_A_455_21#_c_266_n N_VPWR_c_748_n 0.00734734f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_295 N_A_455_21#_c_258_n N_VPWR_c_748_n 0.0016194f $X=3.35 $Y=1.495 $X2=0
+ $Y2=0
cc_296 N_A_455_21#_c_277_p N_VPWR_c_748_n 0.00614279f $X=4.415 $Y=1.875 $X2=0
+ $Y2=0
cc_297 N_A_455_21#_c_277_p N_A_785_297#_M1004_s 0.0035322f $X=4.415 $Y=1.875
+ $X2=-0.19 $Y2=-0.24
cc_298 N_A_455_21#_M1013_s N_A_785_297#_c_867_n 0.00352392f $X=4.395 $Y=1.485
+ $X2=0 $Y2=0
cc_299 N_A_455_21#_c_277_p N_A_785_297#_c_867_n 0.00627679f $X=4.415 $Y=1.875
+ $X2=0 $Y2=0
cc_300 N_A_455_21#_c_291_p N_A_785_297#_c_867_n 0.0127274f $X=4.54 $Y=1.875
+ $X2=0 $Y2=0
cc_301 N_A_455_21#_c_277_p N_A_785_297#_c_870_n 0.0127076f $X=4.415 $Y=1.875
+ $X2=0 $Y2=0
cc_302 N_A_455_21#_c_261_n N_X_c_886_n 3.58584e-19 $X=4.795 $Y=0.815 $X2=0 $Y2=0
cc_303 N_A_455_21#_c_259_n N_VGND_M1022_d 0.00471571f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_304 N_A_455_21#_c_260_n N_VGND_M1022_d 0.0060399f $X=3.445 $Y=0.815 $X2=0
+ $Y2=0
cc_305 N_A_455_21#_c_261_n N_VGND_M1017_s 0.00348805f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_306 N_A_455_21#_c_254_n N_VGND_c_967_n 0.00268723f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_A_455_21#_c_283_p N_VGND_c_968_n 0.0183628f $X=4.07 $Y=0.39 $X2=0 $Y2=0
cc_308 N_A_455_21#_c_261_n N_VGND_c_968_n 0.0131987f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_309 N_A_455_21#_c_300_p N_VGND_c_968_n 0.0223967f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_310 N_A_455_21#_c_261_n N_VGND_c_969_n 6.33233e-19 $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_311 N_A_455_21#_c_259_n N_VGND_c_972_n 0.00199443f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_312 N_A_455_21#_c_283_p N_VGND_c_972_n 0.0222529f $X=4.07 $Y=0.39 $X2=0 $Y2=0
cc_313 N_A_455_21#_c_261_n N_VGND_c_972_n 0.00266636f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_314 N_A_455_21#_c_261_n N_VGND_c_974_n 0.00199443f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_315 N_A_455_21#_c_300_p N_VGND_c_974_n 0.023074f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_316 N_A_455_21#_M1000_d N_VGND_c_982_n 0.00215201f $X=3.935 $Y=0.235 $X2=0
+ $Y2=0
cc_317 N_A_455_21#_M1025_d N_VGND_c_982_n 0.00324782f $X=4.875 $Y=0.235 $X2=0
+ $Y2=0
cc_318 N_A_455_21#_c_254_n N_VGND_c_982_n 0.00600559f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_319 N_A_455_21#_c_255_n N_VGND_c_982_n 0.012103f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_455_21#_c_259_n N_VGND_c_982_n 0.00502905f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_321 N_A_455_21#_c_260_n N_VGND_c_982_n 8.23161e-19 $X=3.445 $Y=0.815 $X2=0
+ $Y2=0
cc_322 N_A_455_21#_c_283_p N_VGND_c_982_n 0.0139016f $X=4.07 $Y=0.39 $X2=0 $Y2=0
cc_323 N_A_455_21#_c_261_n N_VGND_c_982_n 0.0100158f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_324 N_A_455_21#_c_300_p N_VGND_c_982_n 0.0141066f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_325 N_A_455_21#_c_254_n N_VGND_c_984_n 0.00424416f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_326 N_A_455_21#_c_255_n N_VGND_c_984_n 0.00585385f $X=2.87 $Y=0.995 $X2=0
+ $Y2=0
cc_327 N_A_455_21#_c_255_n N_VGND_c_985_n 0.00481673f $X=2.87 $Y=0.995 $X2=0
+ $Y2=0
cc_328 N_A_455_21#_c_256_n N_VGND_c_985_n 0.00843619f $X=3.255 $Y=1.16 $X2=0
+ $Y2=0
cc_329 N_A_455_21#_c_259_n N_VGND_c_985_n 0.0187239f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_330 N_A_455_21#_c_260_n N_VGND_c_985_n 0.0163451f $X=3.445 $Y=0.815 $X2=0
+ $Y2=0
cc_331 N_A_455_21#_c_283_p N_VGND_c_985_n 0.0249664f $X=4.07 $Y=0.39 $X2=0 $Y2=0
cc_332 N_A_455_21#_c_264_n N_VGND_c_985_n 0.0049954f $X=2.87 $Y=1.202 $X2=0
+ $Y2=0
cc_333 N_A1_N_c_392_n N_A2_N_c_477_n 0.0124239f $X=3.86 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_334 N_A1_N_c_391_n N_A2_N_c_481_n 0.0371957f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_335 N_A1_N_c_399_n N_A2_N_c_481_n 0.0118239f $X=5.085 $Y=1.53 $X2=0 $Y2=0
cc_336 N_A1_N_c_395_n N_A2_N_c_481_n 7.38423e-19 $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A1_N_c_393_n N_A2_N_c_482_n 0.0225984f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_338 N_A1_N_c_399_n N_A2_N_c_482_n 0.016887f $X=5.085 $Y=1.53 $X2=0 $Y2=0
cc_339 A1_N N_A2_N_c_482_n 9.66622e-19 $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_340 N_A1_N_c_394_n N_A2_N_c_478_n 0.0103136f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_341 N_A1_N_c_391_n N_A2_N_c_479_n 2.42241e-19 $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_342 N_A1_N_c_393_n N_A2_N_c_479_n 0.00120805f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A1_N_c_399_n N_A2_N_c_479_n 0.0456386f $X=5.085 $Y=1.53 $X2=0 $Y2=0
cc_344 N_A1_N_c_395_n N_A2_N_c_479_n 0.0149938f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_345 A1_N N_A2_N_c_479_n 0.016921f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_346 N_A1_N_c_391_n N_A2_N_c_480_n 0.0264198f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A1_N_c_393_n N_A2_N_c_480_n 0.0260814f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_348 N_A1_N_c_399_n N_A2_N_c_480_n 0.00798993f $X=5.085 $Y=1.53 $X2=0 $Y2=0
cc_349 N_A1_N_c_395_n N_A2_N_c_480_n 0.00372481f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_350 A1_N N_A2_N_c_480_n 0.002584f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_351 N_A1_N_c_394_n N_A_203_47#_c_526_n 0.0122748f $X=5.27 $Y=0.995 $X2=0
+ $Y2=0
cc_352 N_A1_N_c_393_n N_A_203_47#_c_535_n 0.0227843f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_353 A1_N N_A_203_47#_c_535_n 0.00108715f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_354 N_A1_N_c_391_n N_A_203_47#_c_540_n 0.00304243f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_355 N_A1_N_c_399_n N_A_203_47#_c_540_n 0.0493306f $X=5.085 $Y=1.53 $X2=0
+ $Y2=0
cc_356 N_A1_N_c_395_n N_A_203_47#_c_540_n 0.0166195f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_357 A1_N N_A_203_47#_c_540_n 0.030399f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_358 A1_N N_A_203_47#_c_596_n 4.39905e-19 $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_359 N_A1_N_c_393_n N_A_203_47#_c_534_n 0.0265038f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_360 A1_N N_A_203_47#_c_534_n 0.00218276f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_361 N_A1_N_c_393_n N_A_203_47#_c_544_n 6.27534e-19 $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_362 A1_N N_A_203_47#_c_544_n 0.0413009f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_363 A1_N N_VPWR_M1026_d 0.0014745f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_364 N_A1_N_c_391_n N_VPWR_c_752_n 0.0049986f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_365 N_A1_N_c_393_n N_VPWR_c_753_n 0.00314922f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_366 A1_N N_VPWR_c_753_n 0.00550954f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_367 N_A1_N_c_391_n N_VPWR_c_758_n 0.0053025f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_368 N_A1_N_c_393_n N_VPWR_c_758_n 0.00702461f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_369 N_A1_N_c_391_n N_VPWR_c_748_n 0.00821249f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_370 N_A1_N_c_393_n N_VPWR_c_748_n 0.0124596f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_371 N_A1_N_c_399_n N_A_785_297#_M1004_s 0.00161973f $X=5.085 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_372 N_A1_N_c_395_n N_A_785_297#_M1004_s 2.53362e-19 $X=3.78 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_373 N_A1_N_c_399_n N_A_785_297#_M1020_d 0.00176553f $X=5.085 $Y=1.53 $X2=0
+ $Y2=0
cc_374 N_A1_N_c_399_n N_A_785_297#_c_874_n 0.0119288f $X=5.085 $Y=1.53 $X2=0
+ $Y2=0
cc_375 A1_N N_A_785_297#_c_874_n 9.66194e-19 $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_376 N_A1_N_c_393_n N_VGND_c_969_n 2.29798e-19 $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_377 N_A1_N_c_394_n N_VGND_c_969_n 0.00276021f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_378 A1_N N_VGND_c_969_n 0.0057781f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_379 N_A1_N_c_392_n N_VGND_c_972_n 0.00396605f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A1_N_c_394_n N_VGND_c_974_n 0.00585385f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A1_N_c_392_n N_VGND_c_982_n 0.00691418f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_382 N_A1_N_c_394_n N_VGND_c_982_n 0.0107097f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_383 N_A1_N_c_392_n N_VGND_c_985_n 0.00589366f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_384 N_A2_N_c_479_n N_A_203_47#_c_540_n 0.00507142f $X=4.71 $Y=1.16 $X2=0
+ $Y2=0
cc_385 N_A2_N_c_481_n N_VPWR_c_758_n 0.00429453f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_386 N_A2_N_c_482_n N_VPWR_c_758_n 0.00429453f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_387 N_A2_N_c_481_n N_VPWR_c_748_n 0.00609021f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_388 N_A2_N_c_482_n N_VPWR_c_748_n 0.00609021f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_389 N_A2_N_c_481_n N_A_785_297#_c_867_n 0.00995673f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_390 N_A2_N_c_482_n N_A_785_297#_c_867_n 0.0143148f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_391 N_A2_N_c_477_n N_VGND_c_968_n 0.00385467f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_392 N_A2_N_c_478_n N_VGND_c_968_n 0.00365402f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_393 N_A2_N_c_477_n N_VGND_c_972_n 0.00423334f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_394 N_A2_N_c_478_n N_VGND_c_974_n 0.00396605f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_395 N_A2_N_c_477_n N_VGND_c_982_n 0.00610858f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_396 N_A2_N_c_478_n N_VGND_c_982_n 0.00594864f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_397 N_A_203_47#_c_540_n N_A_27_297#_M1011_d 0.00339783f $X=5.67 $Y=1.53 $X2=0
+ $Y2=0
cc_398 N_A_203_47#_c_541_n N_A_27_297#_M1011_d 0.00162011f $X=2.98 $Y=1.53 $X2=0
+ $Y2=0
cc_399 N_A_203_47#_c_530_n N_A_27_297#_c_696_n 0.00630624f $X=2.395 $Y=0.82
+ $X2=0 $Y2=0
cc_400 N_A_203_47#_c_541_n N_A_27_297#_c_696_n 9.93937e-19 $X=2.98 $Y=1.53 $X2=0
+ $Y2=0
cc_401 N_A_203_47#_c_543_n N_A_27_297#_c_696_n 0.00180984f $X=2.61 $Y=1.62 $X2=0
+ $Y2=0
cc_402 N_A_203_47#_M1005_s N_A_27_297#_c_716_n 0.00352392f $X=2.465 $Y=1.485
+ $X2=0 $Y2=0
cc_403 N_A_203_47#_c_543_n N_A_27_297#_c_716_n 0.0177642f $X=2.61 $Y=1.62 $X2=0
+ $Y2=0
cc_404 N_A_203_47#_c_540_n N_A_27_297#_c_725_n 0.00769272f $X=5.67 $Y=1.53 $X2=0
+ $Y2=0
cc_405 N_A_203_47#_c_541_n N_A_27_297#_c_725_n 9.00065e-19 $X=2.98 $Y=1.53 $X2=0
+ $Y2=0
cc_406 N_A_203_47#_c_540_n N_VPWR_M1004_d 0.00112336f $X=5.67 $Y=1.53 $X2=0
+ $Y2=0
cc_407 N_A_203_47#_c_540_n N_VPWR_M1026_d 0.00193338f $X=5.67 $Y=1.53 $X2=0
+ $Y2=0
cc_408 N_A_203_47#_c_540_n N_VPWR_c_752_n 5.37033e-19 $X=5.67 $Y=1.53 $X2=0
+ $Y2=0
cc_409 N_A_203_47#_c_535_n N_VPWR_c_753_n 0.00300743f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_410 N_A_203_47#_c_540_n N_VPWR_c_753_n 0.0080935f $X=5.67 $Y=1.53 $X2=0 $Y2=0
cc_411 N_A_203_47#_c_536_n N_VPWR_c_754_n 0.00300743f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_412 N_A_203_47#_c_537_n N_VPWR_c_754_n 0.00300743f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_413 N_A_203_47#_c_538_n N_VPWR_c_755_n 0.00479105f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_414 N_A_203_47#_c_535_n N_VPWR_c_760_n 0.00702461f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_415 N_A_203_47#_c_536_n N_VPWR_c_760_n 0.00702461f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_416 N_A_203_47#_c_537_n N_VPWR_c_762_n 0.00702461f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_417 N_A_203_47#_c_538_n N_VPWR_c_762_n 0.00702461f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_418 N_A_203_47#_M1005_s N_VPWR_c_748_n 0.00232895f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_419 N_A_203_47#_c_535_n N_VPWR_c_748_n 0.0124344f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_420 N_A_203_47#_c_536_n N_VPWR_c_748_n 0.00693457f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_421 N_A_203_47#_c_537_n N_VPWR_c_748_n 0.00693457f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_422 N_A_203_47#_c_538_n N_VPWR_c_748_n 0.0134606f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_423 N_A_203_47#_c_540_n N_A_785_297#_c_874_n 0.00207051f $X=5.67 $Y=1.53
+ $X2=0 $Y2=0
cc_424 N_A_203_47#_c_596_n N_X_M1003_d 0.00238974f $X=5.815 $Y=1.53 $X2=0 $Y2=0
cc_425 N_A_203_47#_c_544_n N_X_M1003_d 0.00267208f $X=5.822 $Y=1.16 $X2=0 $Y2=0
cc_426 N_A_203_47#_c_526_n N_X_c_897_n 0.00494802f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_427 N_A_203_47#_c_527_n N_X_c_897_n 0.0066581f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_428 N_A_203_47#_c_528_n N_X_c_897_n 5.38967e-19 $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_429 N_A_203_47#_c_536_n N_X_c_900_n 0.0133996f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_430 N_A_203_47#_c_537_n N_X_c_900_n 0.0134427f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_431 N_A_203_47#_c_636_p N_X_c_900_n 0.0164753f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_432 N_A_203_47#_c_534_n N_X_c_900_n 0.00503753f $X=7.125 $Y=1.202 $X2=0 $Y2=0
cc_433 N_A_203_47#_c_636_p N_X_c_904_n 0.0013859f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_434 N_A_203_47#_c_596_n N_X_c_904_n 0.0039661f $X=5.815 $Y=1.53 $X2=0 $Y2=0
cc_435 N_A_203_47#_c_534_n N_X_c_904_n 0.00203852f $X=7.125 $Y=1.202 $X2=0 $Y2=0
cc_436 N_A_203_47#_c_544_n N_X_c_904_n 0.0120687f $X=5.822 $Y=1.16 $X2=0 $Y2=0
cc_437 N_A_203_47#_c_527_n N_X_c_885_n 0.00901745f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_438 N_A_203_47#_c_528_n N_X_c_885_n 0.00901745f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_439 N_A_203_47#_c_636_p N_X_c_885_n 0.0392656f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_440 N_A_203_47#_c_534_n N_X_c_885_n 0.00345541f $X=7.125 $Y=1.202 $X2=0 $Y2=0
cc_441 N_A_203_47#_c_526_n N_X_c_886_n 0.00263405f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_442 N_A_203_47#_c_527_n N_X_c_886_n 0.00116579f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_443 N_A_203_47#_c_636_p N_X_c_886_n 0.00828398f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_444 N_A_203_47#_c_596_n N_X_c_886_n 9.40041e-19 $X=5.815 $Y=1.53 $X2=0 $Y2=0
cc_445 N_A_203_47#_c_534_n N_X_c_886_n 0.00357692f $X=7.125 $Y=1.202 $X2=0 $Y2=0
cc_446 N_A_203_47#_c_544_n N_X_c_886_n 0.0230669f $X=5.822 $Y=1.16 $X2=0 $Y2=0
cc_447 N_A_203_47#_c_527_n N_X_c_918_n 5.19459e-19 $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_448 N_A_203_47#_c_528_n N_X_c_918_n 0.00633209f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_449 N_A_203_47#_c_538_n N_X_c_890_n 0.0215797f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_450 N_A_203_47#_c_636_p N_X_c_890_n 0.00530013f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_451 N_A_203_47#_c_534_n N_X_c_890_n 9.89874e-19 $X=7.125 $Y=1.202 $X2=0 $Y2=0
cc_452 N_A_203_47#_c_529_n N_X_c_887_n 0.0139329f $X=7.15 $Y=0.995 $X2=0 $Y2=0
cc_453 N_A_203_47#_c_636_p N_X_c_887_n 0.00242061f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_454 N_A_203_47#_c_528_n N_X_c_888_n 0.00119508f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_455 N_A_203_47#_c_636_p N_X_c_888_n 0.0303261f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_456 N_A_203_47#_c_534_n N_X_c_888_n 0.00485798f $X=7.125 $Y=1.202 $X2=0 $Y2=0
cc_457 N_A_203_47#_c_537_n N_X_c_891_n 0.00188142f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_458 N_A_203_47#_c_538_n N_X_c_891_n 2.29143e-19 $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_459 N_A_203_47#_c_636_p N_X_c_891_n 0.0200073f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_460 N_A_203_47#_c_534_n N_X_c_891_n 0.00661719f $X=7.125 $Y=1.202 $X2=0 $Y2=0
cc_461 N_A_203_47#_c_529_n X 0.0203559f $X=7.15 $Y=0.995 $X2=0 $Y2=0
cc_462 N_A_203_47#_c_636_p X 0.0116941f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_463 N_A_203_47#_c_530_n N_VGND_M1019_s 0.00165819f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_464 N_A_203_47#_c_530_n N_VGND_c_967_n 0.0116529f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_465 N_A_203_47#_c_526_n N_VGND_c_969_n 0.00275355f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_466 N_A_203_47#_c_540_n N_VGND_c_969_n 0.00390271f $X=5.67 $Y=1.53 $X2=0
+ $Y2=0
cc_467 N_A_203_47#_c_527_n N_VGND_c_970_n 0.00410249f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_468 N_A_203_47#_c_528_n N_VGND_c_970_n 0.00276126f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_469 N_A_203_47#_c_529_n N_VGND_c_971_n 0.00438629f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_470 N_A_203_47#_c_526_n N_VGND_c_976_n 0.00542163f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_471 N_A_203_47#_c_527_n N_VGND_c_976_n 0.00424138f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_203_47#_c_528_n N_VGND_c_978_n 0.00424138f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_473 N_A_203_47#_c_529_n N_VGND_c_978_n 0.00437852f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_203_47#_c_530_n N_VGND_c_980_n 0.00248756f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_475 N_A_203_47#_M1006_d N_VGND_c_982_n 0.00296339f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_476 N_A_203_47#_M1014_s N_VGND_c_982_n 0.00364931f $X=2.425 $Y=0.235 $X2=0
+ $Y2=0
cc_477 N_A_203_47#_c_526_n N_VGND_c_982_n 0.00965669f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_203_47#_c_527_n N_VGND_c_982_n 0.00609398f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_479 N_A_203_47#_c_528_n N_VGND_c_982_n 0.00608656f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_480 N_A_203_47#_c_529_n N_VGND_c_982_n 0.00722755f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_481 N_A_203_47#_c_530_n N_VGND_c_982_n 0.0104586f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_482 N_A_203_47#_c_549_n N_VGND_c_982_n 0.0143448f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_483 N_A_203_47#_c_530_n N_VGND_c_984_n 0.00193763f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_484 N_A_203_47#_c_549_n N_VGND_c_984_n 0.0232294f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_485 N_A_203_47#_c_530_n N_A_119_47#_M1027_s 0.00257722f $X=2.395 $Y=0.82
+ $X2=0 $Y2=0
cc_486 N_A_203_47#_c_532_n N_A_119_47#_c_1090_n 0.0107679f $X=1.2 $Y=0.73 $X2=0
+ $Y2=0
cc_487 N_A_203_47#_M1006_d N_A_119_47#_c_1095_n 0.00507227f $X=1.015 $Y=0.235
+ $X2=0 $Y2=0
cc_488 N_A_203_47#_c_530_n N_A_119_47#_c_1095_n 0.0168825f $X=2.395 $Y=0.82
+ $X2=0 $Y2=0
cc_489 N_A_203_47#_c_532_n N_A_119_47#_c_1095_n 0.0206427f $X=1.2 $Y=0.73 $X2=0
+ $Y2=0
cc_490 N_A_27_297#_c_699_n N_VPWR_M1009_d 0.00370949f $X=1.075 $Y=1.87 $X2=-0.19
+ $Y2=1.305
cc_491 N_A_27_297#_c_704_n N_VPWR_M1023_s 0.00369012f $X=2.015 $Y=1.87 $X2=0
+ $Y2=0
cc_492 N_A_27_297#_c_699_n N_VPWR_c_749_n 0.0139109f $X=1.075 $Y=1.87 $X2=0
+ $Y2=0
cc_493 N_A_27_297#_c_730_p N_VPWR_c_750_n 0.0149311f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_494 N_A_27_297#_c_704_n N_VPWR_c_751_n 0.0139109f $X=2.015 $Y=1.87 $X2=0
+ $Y2=0
cc_495 N_A_27_297#_c_725_n N_VPWR_c_752_n 0.0180653f $X=3.08 $Y=2.3 $X2=0 $Y2=0
cc_496 N_A_27_297#_c_716_n N_VPWR_c_756_n 0.0386815f $X=2.955 $Y=2.38 $X2=0
+ $Y2=0
cc_497 N_A_27_297#_c_734_p N_VPWR_c_756_n 0.015002f $X=2.265 $Y=2.38 $X2=0 $Y2=0
cc_498 N_A_27_297#_c_725_n N_VPWR_c_756_n 0.0154343f $X=3.08 $Y=2.3 $X2=0 $Y2=0
cc_499 N_A_27_297#_c_736_p N_VPWR_c_764_n 0.0161853f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_500 N_A_27_297#_M1009_s N_VPWR_c_748_n 0.00226492f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_501 N_A_27_297#_M1001_d N_VPWR_c_748_n 0.00250817f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_502 N_A_27_297#_M1015_s N_VPWR_c_748_n 0.00241844f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_503 N_A_27_297#_M1011_d N_VPWR_c_748_n 0.00215913f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_504 N_A_27_297#_c_736_p N_VPWR_c_748_n 0.00955092f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_505 N_A_27_297#_c_699_n N_VPWR_c_748_n 0.0141598f $X=1.075 $Y=1.87 $X2=0
+ $Y2=0
cc_506 N_A_27_297#_c_730_p N_VPWR_c_748_n 0.00955092f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_507 N_A_27_297#_c_704_n N_VPWR_c_748_n 0.0141598f $X=2.015 $Y=1.87 $X2=0
+ $Y2=0
cc_508 N_A_27_297#_c_716_n N_VPWR_c_748_n 0.0239184f $X=2.955 $Y=2.38 $X2=0
+ $Y2=0
cc_509 N_A_27_297#_c_734_p N_VPWR_c_748_n 0.00962271f $X=2.265 $Y=2.38 $X2=0
+ $Y2=0
cc_510 N_A_27_297#_c_725_n N_VPWR_c_748_n 0.00938089f $X=3.08 $Y=2.3 $X2=0 $Y2=0
cc_511 N_VPWR_c_748_n N_A_785_297#_M1004_s 0.00241298f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_512 N_VPWR_c_748_n N_A_785_297#_M1020_d 0.00297222f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_758_n N_A_785_297#_c_867_n 0.0536487f $X=5.355 $Y=2.72 $X2=0
+ $Y2=0
cc_514 N_VPWR_c_748_n N_A_785_297#_c_867_n 0.0335411f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_758_n N_A_785_297#_c_870_n 0.0143076f $X=5.355 $Y=2.72 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_748_n N_A_785_297#_c_870_n 0.00938089f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_748_n N_X_M1003_d 0.0031047f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_518 N_VPWR_c_748_n N_X_M1016_d 0.0031047f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_519 N_VPWR_c_760_n N_X_c_936_n 0.0149311f $X=6.295 $Y=2.72 $X2=0 $Y2=0
cc_520 N_VPWR_c_748_n N_X_c_936_n 0.00955092f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_521 N_VPWR_M1012_s N_X_c_900_n 0.0047345f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_522 N_VPWR_c_754_n N_X_c_900_n 0.011587f $X=6.42 $Y=2.33 $X2=0 $Y2=0
cc_523 N_VPWR_c_748_n N_X_c_900_n 0.0142452f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_524 N_VPWR_c_762_n N_X_c_941_n 0.0149311f $X=7.235 $Y=2.72 $X2=0 $Y2=0
cc_525 N_VPWR_c_748_n N_X_c_941_n 0.00955092f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_526 N_VPWR_M1024_s N_X_c_890_n 3.97519e-19 $X=7.215 $Y=1.485 $X2=0 $Y2=0
cc_527 N_VPWR_c_755_n N_X_c_890_n 0.0031267f $X=7.36 $Y=1.99 $X2=0 $Y2=0
cc_528 N_VPWR_M1024_s N_X_c_893_n 0.00277239f $X=7.215 $Y=1.485 $X2=0 $Y2=0
cc_529 N_VPWR_c_755_n N_X_c_893_n 0.0156881f $X=7.36 $Y=1.99 $X2=0 $Y2=0
cc_530 N_X_c_885_n N_VGND_M1007_s 0.00251047f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_531 N_X_c_887_n N_VGND_M1021_s 0.00324195f $X=7.31 $Y=0.815 $X2=0 $Y2=0
cc_532 N_X_c_886_n N_VGND_c_969_n 0.00750114f $X=6.115 $Y=0.815 $X2=0 $Y2=0
cc_533 N_X_c_897_n N_VGND_c_970_n 0.0171386f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_534 N_X_c_885_n N_VGND_c_970_n 0.0127273f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_535 N_X_c_887_n N_VGND_c_971_n 0.013754f $X=7.31 $Y=0.815 $X2=0 $Y2=0
cc_536 N_X_c_897_n N_VGND_c_976_n 0.0198028f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_537 N_X_c_885_n N_VGND_c_976_n 0.00266636f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_538 N_X_c_885_n N_VGND_c_978_n 0.00198695f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_539 N_X_c_918_n N_VGND_c_978_n 0.0205249f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_540 N_X_c_887_n N_VGND_c_978_n 0.00254521f $X=7.31 $Y=0.815 $X2=0 $Y2=0
cc_541 N_X_c_887_n N_VGND_c_981_n 0.00386917f $X=7.31 $Y=0.815 $X2=0 $Y2=0
cc_542 N_X_M1002_d N_VGND_c_982_n 0.00256339f $X=5.765 $Y=0.235 $X2=0 $Y2=0
cc_543 N_X_M1008_d N_VGND_c_982_n 0.00305225f $X=6.705 $Y=0.235 $X2=0 $Y2=0
cc_544 N_X_c_897_n N_VGND_c_982_n 0.0139751f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_545 N_X_c_885_n N_VGND_c_982_n 0.00972452f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_546 N_X_c_918_n N_VGND_c_982_n 0.0141809f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_547 N_X_c_887_n N_VGND_c_982_n 0.0122098f $X=7.31 $Y=0.815 $X2=0 $Y2=0
cc_548 N_VGND_c_982_n N_A_119_47#_M1018_d 0.00215206f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_549 N_VGND_c_982_n N_A_119_47#_M1027_s 0.00265108f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_550 N_VGND_c_966_n N_A_119_47#_c_1091_n 0.0172916f $X=0.26 $Y=0.39 $X2=0
+ $Y2=0
cc_551 N_VGND_c_980_n N_A_119_47#_c_1091_n 0.0186088f $X=2.055 $Y=0 $X2=0 $Y2=0
cc_552 N_VGND_c_982_n N_A_119_47#_c_1091_n 0.0111017f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_c_966_n N_A_119_47#_c_1090_n 0.0307592f $X=0.26 $Y=0.39 $X2=0
+ $Y2=0
cc_554 N_VGND_c_980_n N_A_119_47#_c_1095_n 0.0576174f $X=2.055 $Y=0 $X2=0 $Y2=0
cc_555 N_VGND_c_982_n N_A_119_47#_c_1095_n 0.0366908f $X=7.59 $Y=0 $X2=0 $Y2=0
