* File: sky130_fd_sc_hdll__o22ai_4.pex.spice
* Created: Thu Aug 27 19:21:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 29 34 48 51 55
c121 29 0 1.53825e-20 $X=3.79 $Y=1.16
c122 16 0 2.98607e-20 $X=1.49 $Y=0.995
r123 48 49 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=1.465 $Y=1.202
+ $X2=1.49 $Y2=1.202
r124 46 48 14.8606 $w=3.73e-07 $l=1.15e-07 $layer=POLY_cond $X=1.35 $Y=1.202
+ $X2=1.465 $Y2=1.202
r125 44 46 42.6434 $w=3.73e-07 $l=3.3e-07 $layer=POLY_cond $X=1.02 $Y=1.202
+ $X2=1.35 $Y2=1.202
r126 43 44 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.995 $Y=1.202
+ $X2=1.02 $Y2=1.202
r127 42 55 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=0.96 $Y=1.175
+ $X2=1.15 $Y2=1.175
r128 41 43 4.52279 $w=3.73e-07 $l=3.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.995 $Y2=1.202
r129 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.96
+ $Y=1.16 $X2=0.96 $Y2=1.16
r130 39 41 52.9812 $w=3.73e-07 $l=4.1e-07 $layer=POLY_cond $X=0.55 $Y=1.202
+ $X2=0.96 $Y2=1.202
r131 38 39 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.525 $Y=1.202
+ $X2=0.55 $Y2=1.202
r132 34 51 4.44006 $w=2e-07 $l=1.57e-07 $layer=LI1_cond $X=1.407 $Y=1.175
+ $X2=1.25 $Y2=1.175
r133 34 51 2.38455 $w=1.98e-07 $l=4.3e-08 $layer=LI1_cond $X=1.207 $Y=1.175
+ $X2=1.25 $Y2=1.175
r134 34 55 3.16091 $w=1.98e-07 $l=5.7e-08 $layer=LI1_cond $X=1.207 $Y=1.175
+ $X2=1.15 $Y2=1.175
r135 34 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.35
+ $Y=1.16 $X2=1.35 $Y2=1.16
r136 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.79
+ $Y=1.16 $X2=3.79 $Y2=1.16
r137 27 34 5.45027 $w=3.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.407 $Y=1.445
+ $X2=1.407 $Y2=1.275
r138 26 27 7.64049 $w=1.7e-07 $l=1.95944e-07 $layer=LI1_cond $X=1.565 $Y=1.53
+ $X2=1.407 $Y2=1.445
r139 25 29 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.827 $Y=1.53
+ $X2=3.827 $Y2=1.16
r140 25 26 134.396 $w=1.68e-07 $l=2.06e-06 $layer=LI1_cond $X=3.625 $Y=1.53
+ $X2=1.565 $Y2=1.53
r141 22 30 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.84 $Y=0.995
+ $X2=3.815 $Y2=1.16
r142 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.84 $Y=0.995
+ $X2=3.84 $Y2=0.56
r143 19 30 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.815 $Y=1.41
+ $X2=3.815 $Y2=1.16
r144 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.815 $Y=1.41
+ $X2=3.815 $Y2=1.985
r145 16 49 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.49 $Y=0.995
+ $X2=1.49 $Y2=1.202
r146 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.49 $Y=0.995
+ $X2=1.49 $Y2=0.56
r147 13 48 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.465 $Y=1.41
+ $X2=1.465 $Y2=1.202
r148 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.465 $Y=1.41
+ $X2=1.465 $Y2=1.985
r149 10 44 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.02 $Y=0.995
+ $X2=1.02 $Y2=1.202
r150 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.02 $Y=0.995
+ $X2=1.02 $Y2=0.56
r151 7 43 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.995 $Y=1.41
+ $X2=0.995 $Y2=1.202
r152 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.995 $Y=1.41
+ $X2=0.995 $Y2=1.985
r153 4 39 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.55 $Y=0.995
+ $X2=0.55 $Y2=1.202
r154 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.55 $Y=0.995
+ $X2=0.55 $Y2=0.56
r155 1 38 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.525 $Y=1.41
+ $X2=0.525 $Y2=1.202
r156 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.525 $Y=1.41
+ $X2=0.525 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 44
r81 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.345 $Y=1.202
+ $X2=3.37 $Y2=1.202
r82 37 39 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=3.23 $Y=1.202
+ $X2=3.345 $Y2=1.202
r83 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.23
+ $Y=1.16 $X2=3.23 $Y2=1.16
r84 35 37 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=2.875 $Y=1.202
+ $X2=3.23 $Y2=1.202
r85 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.85 $Y=1.202
+ $X2=2.875 $Y2=1.202
r86 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.405 $Y=1.202
+ $X2=2.85 $Y2=1.202
r87 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.38 $Y=1.202
+ $X2=2.405 $Y2=1.202
r88 31 44 26.0636 $w=1.98e-07 $l=4.7e-07 $layer=LI1_cond $X=2.06 $Y=1.175
+ $X2=2.53 $Y2=1.175
r89 30 32 41.4624 $w=3.72e-07 $l=3.2e-07 $layer=POLY_cond $X=2.06 $Y=1.202
+ $X2=2.38 $Y2=1.202
r90 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.06
+ $Y=1.16 $X2=2.06 $Y2=1.16
r91 28 30 16.1962 $w=3.72e-07 $l=1.25e-07 $layer=POLY_cond $X=1.935 $Y=1.202
+ $X2=2.06 $Y2=1.202
r92 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.91 $Y=1.202
+ $X2=1.935 $Y2=1.202
r93 25 38 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=2.78 $Y=1.175
+ $X2=3.23 $Y2=1.175
r94 25 44 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=2.78 $Y=1.175
+ $X2=2.53 $Y2=1.175
r95 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.37 $Y=0.995
+ $X2=3.37 $Y2=1.202
r96 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.37 $Y=0.995
+ $X2=3.37 $Y2=0.56
r97 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.345 $Y=1.41
+ $X2=3.345 $Y2=1.202
r98 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.345 $Y=1.41
+ $X2=3.345 $Y2=1.985
r99 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.875 $Y=1.41
+ $X2=2.875 $Y2=1.202
r100 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.875 $Y=1.41
+ $X2=2.875 $Y2=1.985
r101 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.85 $Y=0.995
+ $X2=2.85 $Y2=1.202
r102 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.85 $Y=0.995
+ $X2=2.85 $Y2=0.56
r103 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.405 $Y=1.41
+ $X2=2.405 $Y2=1.202
r104 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.405 $Y=1.41
+ $X2=2.405 $Y2=1.985
r105 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.38 $Y=0.995
+ $X2=2.38 $Y2=1.202
r106 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.38 $Y=0.995
+ $X2=2.38 $Y2=0.56
r107 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.935 $Y=1.41
+ $X2=1.935 $Y2=1.202
r108 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.935 $Y=1.41
+ $X2=1.935 $Y2=1.985
r109 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.91 $Y=0.995
+ $X2=1.91 $Y2=1.202
r110 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.91 $Y=0.995
+ $X2=1.91 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 29 32 41 45 50
c108 10 0 1.63013e-19 $X=4.805 $Y=1.41
c109 1 0 1.69878e-19 $X=4.31 $Y=0.995
r110 41 42 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.275 $Y=1.202
+ $X2=5.3 $Y2=1.202
r111 40 45 7.52372 $w=6.18e-07 $l=3.9e-07 $layer=LI1_cond $X=5.22 $Y=1.305
+ $X2=4.83 $Y2=1.305
r112 39 41 7.12634 $w=3.72e-07 $l=5.5e-08 $layer=POLY_cond $X=5.22 $Y=1.202
+ $X2=5.275 $Y2=1.202
r113 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.22
+ $Y=1.16 $X2=5.22 $Y2=1.16
r114 37 39 53.7715 $w=3.72e-07 $l=4.15e-07 $layer=POLY_cond $X=4.805 $Y=1.202
+ $X2=5.22 $Y2=1.202
r115 36 37 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.78 $Y=1.202
+ $X2=4.805 $Y2=1.202
r116 35 36 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.335 $Y=1.202
+ $X2=4.78 $Y2=1.202
r117 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.31 $Y=1.202
+ $X2=4.335 $Y2=1.202
r118 32 50 10.19 $w=6.18e-07 $l=1.6e-07 $layer=LI1_cond $X=5.33 $Y=1.305
+ $X2=5.49 $Y2=1.305
r119 32 40 2.12207 $w=6.18e-07 $l=1.1e-07 $layer=LI1_cond $X=5.33 $Y=1.305
+ $X2=5.22 $Y2=1.305
r120 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.6
+ $Y=1.16 $X2=7.6 $Y2=1.16
r121 27 29 12.1647 $w=2.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.6 $Y=1.445
+ $X2=7.6 $Y2=1.16
r122 25 27 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.465 $Y=1.53
+ $X2=7.6 $Y2=1.445
r123 25 50 128.85 $w=1.68e-07 $l=1.975e-06 $layer=LI1_cond $X=7.465 $Y=1.53
+ $X2=5.49 $Y2=1.53
r124 22 30 38.5462 $w=3.19e-07 $l=1.69926e-07 $layer=POLY_cond $X=7.65 $Y=0.995
+ $X2=7.64 $Y2=1.16
r125 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.65 $Y=0.995
+ $X2=7.65 $Y2=0.56
r126 19 30 46.8511 $w=3.19e-07 $l=2.57391e-07 $layer=POLY_cond $X=7.625 $Y=1.41
+ $X2=7.64 $Y2=1.16
r127 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.625 $Y=1.41
+ $X2=7.625 $Y2=1.985
r128 16 42 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.3 $Y=0.995
+ $X2=5.3 $Y2=1.202
r129 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.3 $Y=0.995
+ $X2=5.3 $Y2=0.56
r130 13 41 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.275 $Y=1.41
+ $X2=5.275 $Y2=1.202
r131 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.275 $Y=1.41
+ $X2=5.275 $Y2=1.985
r132 10 37 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.805 $Y=1.41
+ $X2=4.805 $Y2=1.202
r133 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.805 $Y=1.41
+ $X2=4.805 $Y2=1.985
r134 7 36 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.78 $Y=0.995
+ $X2=4.78 $Y2=1.202
r135 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.78 $Y=0.995
+ $X2=4.78 $Y2=0.56
r136 4 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.335 $Y=1.41
+ $X2=4.335 $Y2=1.202
r137 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.335 $Y=1.41
+ $X2=4.335 $Y2=1.985
r138 1 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.31 $Y=0.995
+ $X2=4.31 $Y2=1.202
r139 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.31 $Y=0.995
+ $X2=4.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%B2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 39 44
r63 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.155 $Y=1.202
+ $X2=7.18 $Y2=1.202
r64 37 39 20.7312 $w=3.72e-07 $l=1.6e-07 $layer=POLY_cond $X=6.995 $Y=1.202
+ $X2=7.155 $Y2=1.202
r65 35 37 40.1667 $w=3.72e-07 $l=3.1e-07 $layer=POLY_cond $X=6.685 $Y=1.202
+ $X2=6.995 $Y2=1.202
r66 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.66 $Y=1.202
+ $X2=6.685 $Y2=1.202
r67 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=6.215 $Y=1.202
+ $X2=6.66 $Y2=1.202
r68 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.19 $Y=1.202
+ $X2=6.215 $Y2=1.202
r69 31 44 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=5.825 $Y=1.175
+ $X2=6.21 $Y2=1.175
r70 30 32 47.293 $w=3.72e-07 $l=3.65e-07 $layer=POLY_cond $X=5.825 $Y=1.202
+ $X2=6.19 $Y2=1.202
r71 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.825
+ $Y=1.16 $X2=5.825 $Y2=1.16
r72 28 30 10.3656 $w=3.72e-07 $l=8e-08 $layer=POLY_cond $X=5.745 $Y=1.202
+ $X2=5.825 $Y2=1.202
r73 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.72 $Y=1.202
+ $X2=5.745 $Y2=1.202
r74 25 44 38.8182 $w=1.98e-07 $l=7e-07 $layer=LI1_cond $X=6.91 $Y=1.175 $X2=6.21
+ $Y2=1.175
r75 25 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.995
+ $Y=1.16 $X2=6.995 $Y2=1.16
r76 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.18 $Y=0.995
+ $X2=7.18 $Y2=1.202
r77 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.18 $Y=0.995
+ $X2=7.18 $Y2=0.56
r78 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.155 $Y=1.41
+ $X2=7.155 $Y2=1.202
r79 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.155 $Y=1.41
+ $X2=7.155 $Y2=1.985
r80 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.685 $Y=1.41
+ $X2=6.685 $Y2=1.202
r81 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.685 $Y=1.41
+ $X2=6.685 $Y2=1.985
r82 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.66 $Y=0.995
+ $X2=6.66 $Y2=1.202
r83 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.66 $Y=0.995
+ $X2=6.66 $Y2=0.56
r84 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.215 $Y=1.41
+ $X2=6.215 $Y2=1.202
r85 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.215 $Y=1.41
+ $X2=6.215 $Y2=1.985
r86 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.19 $Y=0.995
+ $X2=6.19 $Y2=1.202
r87 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.19 $Y=0.995 $X2=6.19
+ $Y2=0.56
r88 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.745 $Y=1.41
+ $X2=5.745 $Y2=1.202
r89 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.745 $Y=1.41
+ $X2=5.745 $Y2=1.985
r90 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.72 $Y=0.995
+ $X2=5.72 $Y2=1.202
r91 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.72 $Y=0.995 $X2=5.72
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%VPWR 1 2 3 4 5 16 18 22 26 30 34 36 38 41
+ 42 44 45 46 58 69 73
r116 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r117 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 64 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r119 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r120 61 64 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=7.59 $Y2=2.72
r121 60 63 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=7.59 $Y2=2.72
r122 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r123 58 72 4.09394 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=7.735 $Y=2.72
+ $X2=8.007 $Y2=2.72
r124 58 63 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.735 $Y=2.72
+ $X2=7.59 $Y2=2.72
r125 57 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r126 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r127 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r128 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r129 51 54 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r130 51 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r131 50 53 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r132 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r133 48 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.23 $Y2=2.72
r134 48 50 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.61 $Y2=2.72
r135 46 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r136 46 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r137 44 56 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.925 $Y=2.72
+ $X2=4.83 $Y2=2.72
r138 44 45 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.925 $Y=2.72
+ $X2=5.045 $Y2=2.72
r139 43 60 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.165 $Y=2.72
+ $X2=5.29 $Y2=2.72
r140 43 45 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.165 $Y=2.72
+ $X2=5.045 $Y2=2.72
r141 41 53 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.965 $Y=2.72
+ $X2=3.91 $Y2=2.72
r142 41 42 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.965 $Y=2.72
+ $X2=4.075 $Y2=2.72
r143 40 56 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.83 $Y2=2.72
r144 40 42 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.075 $Y2=2.72
r145 36 72 3.26612 $w=2.8e-07 $l=1.69245e-07 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=8.007 $Y2=2.72
r146 36 38 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=7.875 $Y2=2.3
r147 32 45 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=2.635
+ $X2=5.045 $Y2=2.72
r148 32 34 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=5.045 $Y=2.635
+ $X2=5.045 $Y2=2.3
r149 28 42 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=2.635
+ $X2=4.075 $Y2=2.72
r150 28 30 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=4.075 $Y=2.635
+ $X2=4.075 $Y2=2.3
r151 24 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.72
r152 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.3
r153 23 66 3.95154 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=2.72
+ $X2=0.207 $Y2=2.72
r154 22 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.105 $Y=2.72
+ $X2=1.23 $Y2=2.72
r155 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.105 $Y=2.72
+ $X2=0.415 $Y2=2.72
r156 18 21 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.29 $Y=1.62
+ $X2=0.29 $Y2=2.3
r157 16 66 3.19163 $w=2.5e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.29 $Y=2.635
+ $X2=0.207 $Y2=2.72
r158 16 21 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.29 $Y=2.635
+ $X2=0.29 $Y2=2.3
r159 5 38 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.715
+ $Y=1.485 $X2=7.86 $Y2=2.3
r160 4 34 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.485 $X2=5.04 $Y2=2.3
r161 3 30 600 $w=1.7e-07 $l=9.02773e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.485 $X2=4.09 $Y2=2.3
r162 2 26 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.485 $X2=1.23 $Y2=2.3
r163 1 21 400 $w=1.7e-07 $l=8.89129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.29 $Y2=2.3
r164 1 18 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.29 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%A_123_297# 1 2 3 4 15 19 21 26 27 28 29 33
+ 38
r55 38 40 3.17915 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=3.6 $Y=2.3 $X2=3.6
+ $Y2=2.38
r56 33 35 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.64 $Y=2.3 $X2=2.64
+ $Y2=2.38
r57 30 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.765 $Y=2.38
+ $X2=2.64 $Y2=2.38
r58 29 40 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.455 $Y=2.38
+ $X2=3.6 $Y2=2.38
r59 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.455 $Y=2.38
+ $X2=2.765 $Y2=2.38
r60 27 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.515 $Y=2.38
+ $X2=2.64 $Y2=2.38
r61 27 28 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.515 $Y=2.38
+ $X2=1.785 $Y2=2.38
r62 24 28 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.68 $Y=2.295
+ $X2=1.785 $Y2=2.38
r63 24 26 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=1.68 $Y=2.295
+ $X2=1.68 $Y2=1.96
r64 23 26 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=1.68 $Y=1.955
+ $X2=1.68 $Y2=1.96
r65 22 31 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.885 $Y=1.87
+ $X2=0.76 $Y2=1.87
r66 21 23 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.575 $Y=1.87
+ $X2=1.68 $Y2=1.955
r67 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.575 $Y=1.87
+ $X2=0.885 $Y2=1.87
r68 17 31 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=1.955
+ $X2=0.76 $Y2=1.87
r69 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.76 $Y=1.955
+ $X2=0.76 $Y2=1.96
r70 13 31 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=1.785
+ $X2=0.76 $Y2=1.87
r71 13 15 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=1.785
+ $X2=0.76 $Y2=1.62
r72 4 38 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.485 $X2=3.58 $Y2=2.3
r73 3 33 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.485 $X2=2.64 $Y2=2.3
r74 2 26 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.555
+ $Y=1.485 $X2=1.7 $Y2=1.96
r75 1 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.615
+ $Y=1.485 $X2=0.76 $Y2=1.96
r76 1 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.485 $X2=0.76 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%Y 1 2 3 4 5 6 7 8 25 28 29 30 31 39 41 44
+ 45 54 57 62 67 72
c120 54 0 1.47631e-19 $X=4.2 $Y=1.87
r121 70 72 1.50053 $w=1.68e-07 $l=2.3e-08 $layer=LI1_cond $X=3.235 $Y=1.87
+ $X2=3.258 $Y2=1.87
r122 67 77 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.11 $Y=1.87 $X2=3.11
+ $Y2=1.96
r123 67 70 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.11 $Y=1.87
+ $X2=3.235 $Y2=1.87
r124 67 72 3.06631 $w=1.68e-07 $l=4.7e-08 $layer=LI1_cond $X=3.305 $Y=1.87
+ $X2=3.258 $Y2=1.87
r125 62 65 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=6.92 $Y=1.87 $X2=6.92
+ $Y2=1.96
r126 57 60 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.98 $Y=1.87 $X2=5.98
+ $Y2=1.96
r127 54 67 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=4.2 $Y=1.87
+ $X2=3.305 $Y2=1.87
r128 45 48 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=2.125 $Y=1.87
+ $X2=2.125 $Y2=1.96
r129 43 44 41.9663 $w=2.63e-07 $l=9.65e-07 $layer=LI1_cond $X=8.037 $Y=0.82
+ $X2=8.037 $Y2=1.785
r130 42 62 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.045 $Y=1.87
+ $X2=6.92 $Y2=1.87
r131 41 44 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=7.905 $Y=1.87
+ $X2=8.037 $Y2=1.785
r132 41 42 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=7.905 $Y=1.87
+ $X2=7.045 $Y2=1.87
r133 40 57 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.105 $Y=1.87
+ $X2=5.98 $Y2=1.87
r134 39 62 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.795 $Y=1.87
+ $X2=6.92 $Y2=1.87
r135 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.795 $Y=1.87
+ $X2=6.105 $Y2=1.87
r136 36 38 59.574 $w=1.73e-07 $l=9.4e-07 $layer=LI1_cond $X=6.45 $Y=0.732
+ $X2=7.39 $Y2=0.732
r137 34 36 59.574 $w=1.73e-07 $l=9.4e-07 $layer=LI1_cond $X=5.51 $Y=0.732
+ $X2=6.45 $Y2=0.732
r138 32 56 3.85122 $w=1.75e-07 $l=1.1e-07 $layer=LI1_cond $X=4.575 $Y=0.732
+ $X2=4.465 $Y2=0.732
r139 32 34 59.2571 $w=1.73e-07 $l=9.35e-07 $layer=LI1_cond $X=4.575 $Y=0.732
+ $X2=5.51 $Y2=0.732
r140 31 43 7.19411 $w=1.75e-07 $l=1.70411e-07 $layer=LI1_cond $X=7.905 $Y=0.732
+ $X2=8.037 $Y2=0.82
r141 31 38 32.639 $w=1.73e-07 $l=5.15e-07 $layer=LI1_cond $X=7.905 $Y=0.732
+ $X2=7.39 $Y2=0.732
r142 30 50 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.465 $Y=1.53
+ $X2=4.285 $Y2=1.53
r143 29 56 3.08098 $w=2.2e-07 $l=8.8e-08 $layer=LI1_cond $X=4.465 $Y=0.82
+ $X2=4.465 $Y2=0.732
r144 29 30 32.7399 $w=2.18e-07 $l=6.25e-07 $layer=LI1_cond $X=4.465 $Y=0.82
+ $X2=4.465 $Y2=1.445
r145 28 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.285 $Y=1.785
+ $X2=4.2 $Y2=1.87
r146 27 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.285 $Y=1.615
+ $X2=4.285 $Y2=1.53
r147 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.285 $Y=1.615
+ $X2=4.285 $Y2=1.785
r148 26 45 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.295 $Y=1.87
+ $X2=2.125 $Y2=1.87
r149 25 67 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.985 $Y=1.87
+ $X2=3.11 $Y2=1.87
r150 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.985 $Y=1.87
+ $X2=2.295 $Y2=1.87
r151 8 65 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=6.775
+ $Y=1.485 $X2=6.92 $Y2=1.96
r152 7 60 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=1.485 $X2=5.98 $Y2=1.96
r153 6 77 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.965
+ $Y=1.485 $X2=3.11 $Y2=1.96
r154 5 48 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.025
+ $Y=1.485 $X2=2.17 $Y2=1.96
r155 4 38 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=7.255
+ $Y=0.235 $X2=7.39 $Y2=0.73
r156 3 36 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=6.265
+ $Y=0.235 $X2=6.45 $Y2=0.73
r157 2 34 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.375
+ $Y=0.235 $X2=5.51 $Y2=0.73
r158 1 56 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.235 $X2=4.57 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%A_885_297# 1 2 3 4 15 16 21 22 23 26 27 30
+ 35
r52 35 37 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=7.39 $Y=2.3 $X2=7.39
+ $Y2=2.38
r53 30 32 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=6.45 $Y=2.3 $X2=6.45
+ $Y2=2.38
r54 26 27 8.82369 $w=3.53e-07 $l=1.75e-07 $layer=LI1_cond $X=4.532 $Y=2.3
+ $X2=4.532 $Y2=2.125
r55 24 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.575 $Y=2.38
+ $X2=6.45 $Y2=2.38
r56 23 37 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.265 $Y=2.38
+ $X2=7.39 $Y2=2.38
r57 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.265 $Y=2.38
+ $X2=6.575 $Y2=2.38
r58 21 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.325 $Y=2.38
+ $X2=6.45 $Y2=2.38
r59 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.325 $Y=2.38
+ $X2=5.635 $Y2=2.38
r60 18 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.51 $Y=2.295
+ $X2=5.635 $Y2=2.38
r61 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.51 $Y=2.295
+ $X2=5.51 $Y2=1.96
r62 17 20 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.51 $Y=1.955
+ $X2=5.51 $Y2=1.96
r63 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.385 $Y=1.87
+ $X2=5.51 $Y2=1.955
r64 15 16 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.385 $Y=1.87
+ $X2=4.71 $Y2=1.87
r65 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.625 $Y=1.955
+ $X2=4.71 $Y2=1.87
r66 13 27 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.625 $Y=1.955
+ $X2=4.625 $Y2=2.125
r67 4 35 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.485 $X2=7.39 $Y2=2.3
r68 3 30 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=1.485 $X2=6.45 $Y2=2.3
r69 2 20 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.365
+ $Y=1.485 $X2=5.51 $Y2=1.96
r70 1 26 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.57 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%A_33_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 52 55 64 66 67 68
c119 67 0 2.98607e-20 $X=2.145 $Y=0.815
c120 50 0 1.69878e-19 $X=3.835 $Y=0.82
r121 62 64 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=6.92 $Y=0.365
+ $X2=7.86 $Y2=0.365
r122 60 62 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=5.98 $Y=0.365
+ $X2=6.92 $Y2=0.365
r123 58 60 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=5.04 $Y=0.365
+ $X2=5.98 $Y2=0.365
r124 56 70 4.47512 $w=2.2e-07 $l=1.75e-07 $layer=LI1_cond $X=4.185 $Y=0.365
+ $X2=4.01 $Y2=0.365
r125 56 58 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=4.185 $Y=0.365
+ $X2=5.04 $Y2=0.365
r126 53 55 0.164635 $w=3.48e-07 $l=5e-09 $layer=LI1_cond $X=4.01 $Y=0.735
+ $X2=4.01 $Y2=0.73
r127 52 70 2.81293 $w=3.5e-07 $l=1.1e-07 $layer=LI1_cond $X=4.01 $Y=0.475
+ $X2=4.01 $Y2=0.365
r128 52 55 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.01 $Y=0.475
+ $X2=4.01 $Y2=0.73
r129 51 68 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=3.275 $Y=0.82
+ $X2=3.085 $Y2=0.815
r130 50 53 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=3.835 $Y=0.82
+ $X2=4.01 $Y2=0.735
r131 50 51 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.835 $Y=0.82
+ $X2=3.275 $Y2=0.82
r132 46 68 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.085 $Y=0.725
+ $X2=3.085 $Y2=0.815
r133 46 48 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.085 $Y=0.725
+ $X2=3.085 $Y2=0.39
r134 45 67 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=2.335 $Y=0.815
+ $X2=2.145 $Y2=0.815
r135 44 68 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=2.895 $Y=0.815
+ $X2=3.085 $Y2=0.815
r136 44 45 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.895 $Y=0.815
+ $X2=2.335 $Y2=0.815
r137 40 67 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=2.145 $Y=0.725
+ $X2=2.145 $Y2=0.815
r138 40 42 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.145 $Y=0.725
+ $X2=2.145 $Y2=0.39
r139 39 66 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=1.395 $Y=0.82
+ $X2=1.205 $Y2=0.815
r140 38 67 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=1.955 $Y=0.82
+ $X2=2.145 $Y2=0.815
r141 38 39 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.955 $Y=0.82
+ $X2=1.395 $Y2=0.82
r142 34 66 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.205 $Y=0.725
+ $X2=1.205 $Y2=0.815
r143 34 36 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.205 $Y=0.725
+ $X2=1.205 $Y2=0.39
r144 32 66 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=1.015 $Y=0.815
+ $X2=1.205 $Y2=0.815
r145 32 33 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.015 $Y=0.815
+ $X2=0.455 $Y2=0.815
r146 28 33 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.29 $Y=0.725
+ $X2=0.455 $Y2=0.815
r147 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.29 $Y=0.725
+ $X2=0.29 $Y2=0.39
r148 9 64 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.725
+ $Y=0.235 $X2=7.86 $Y2=0.39
r149 8 62 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.735
+ $Y=0.235 $X2=6.92 $Y2=0.39
r150 7 60 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.235 $X2=5.98 $Y2=0.39
r151 6 58 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.855
+ $Y=0.235 $X2=5.04 $Y2=0.39
r152 5 70 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.235 $X2=4.05 $Y2=0.39
r153 5 55 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.235 $X2=4.05 $Y2=0.73
r154 4 48 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.925
+ $Y=0.235 $X2=3.11 $Y2=0.39
r155 3 42 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.985
+ $Y=0.235 $X2=2.17 $Y2=0.39
r156 2 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.095
+ $Y=0.235 $X2=1.23 $Y2=0.39
r157 1 30 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_4%VGND 1 2 3 4 17 21 25 29 32 33 35 36 38 39
+ 40 56 57 60
r104 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r105 56 57 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r106 54 57 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=3.91 $Y=0 $X2=8.05
+ $Y2=0
r107 53 56 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=8.05
+ $Y2=0
r108 53 54 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r109 51 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r110 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r111 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r112 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r113 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r114 45 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r115 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r116 42 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.76
+ $Y2=0
r117 42 44 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r118 40 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r119 38 50 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.45
+ $Y2=0
r120 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.58
+ $Y2=0
r121 37 53 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.91
+ $Y2=0
r122 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.58
+ $Y2=0
r123 35 47 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.555 $Y=0 $X2=2.53
+ $Y2=0
r124 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=0 $X2=2.64
+ $Y2=0
r125 34 50 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=3.45 $Y2=0
r126 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.64
+ $Y2=0
r127 32 44 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.61
+ $Y2=0
r128 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.7
+ $Y2=0
r129 31 47 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.53 $Y2=0
r130 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.7
+ $Y2=0
r131 27 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.58 $Y2=0
r132 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.58 $Y2=0.39
r133 23 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0
r134 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0.39
r135 19 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r136 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.7 $Y=0.085
+ $X2=1.7 $Y2=0.39
r137 15 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0
r138 15 17 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.39
r139 4 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.235 $X2=3.58 $Y2=0.39
r140 3 25 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.455
+ $Y=0.235 $X2=2.64 $Y2=0.39
r141 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.235 $X2=1.7 $Y2=0.39
r142 1 17 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.235 $X2=0.76 $Y2=0.39
.ends

