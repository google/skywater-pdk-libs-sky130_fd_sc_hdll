* File: sky130_fd_sc_hdll__o22ai_2.pxi.spice
* Created: Wed Sep  2 08:45:44 2020
* 
x_PM_SKY130_FD_SC_HDLL__O22AI_2%B1 N_B1_c_66_n N_B1_M1006_g N_B1_c_70_n
+ N_B1_M1001_g N_B1_c_71_n N_B1_M1011_g N_B1_c_67_n N_B1_M1013_g B1 N_B1_c_68_n
+ N_B1_c_69_n B1 PM_SKY130_FD_SC_HDLL__O22AI_2%B1
x_PM_SKY130_FD_SC_HDLL__O22AI_2%B2 N_B2_c_104_n N_B2_M1007_g N_B2_c_108_n
+ N_B2_M1003_g N_B2_c_109_n N_B2_M1005_g N_B2_c_105_n N_B2_M1012_g B2
+ N_B2_c_106_n N_B2_c_107_n B2 PM_SKY130_FD_SC_HDLL__O22AI_2%B2
x_PM_SKY130_FD_SC_HDLL__O22AI_2%A2 N_A2_c_145_n N_A2_M1002_g N_A2_c_149_n
+ N_A2_M1000_g N_A2_c_150_n N_A2_M1015_g N_A2_c_146_n N_A2_M1009_g A2
+ N_A2_c_147_n N_A2_c_148_n A2 PM_SKY130_FD_SC_HDLL__O22AI_2%A2
x_PM_SKY130_FD_SC_HDLL__O22AI_2%A1 N_A1_c_196_n N_A1_M1004_g N_A1_c_200_n
+ N_A1_M1008_g N_A1_c_201_n N_A1_M1010_g N_A1_c_197_n N_A1_M1014_g A1
+ N_A1_c_199_n A1 PM_SKY130_FD_SC_HDLL__O22AI_2%A1
x_PM_SKY130_FD_SC_HDLL__O22AI_2%A_27_297# N_A_27_297#_M1001_s
+ N_A_27_297#_M1011_s N_A_27_297#_M1005_d N_A_27_297#_c_237_n
+ N_A_27_297#_c_257_p N_A_27_297#_c_238_n N_A_27_297#_c_239_n
+ N_A_27_297#_c_252_p N_A_27_297#_c_248_n N_A_27_297#_c_267_p
+ PM_SKY130_FD_SC_HDLL__O22AI_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__O22AI_2%VPWR N_VPWR_M1001_d N_VPWR_M1008_s
+ N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n VPWR
+ N_VPWR_c_276_n N_VPWR_c_271_n N_VPWR_c_278_n
+ PM_SKY130_FD_SC_HDLL__O22AI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O22AI_2%Y N_Y_M1006_d N_Y_M1007_s N_Y_M1003_s
+ N_Y_M1000_d N_Y_c_325_n N_Y_c_326_n N_Y_c_328_n N_Y_c_329_n N_Y_c_330_n
+ N_Y_c_331_n N_Y_c_332_n Y PM_SKY130_FD_SC_HDLL__O22AI_2%Y
x_PM_SKY130_FD_SC_HDLL__O22AI_2%A_515_297# N_A_515_297#_M1000_s
+ N_A_515_297#_M1015_s N_A_515_297#_M1010_d N_A_515_297#_c_402_n
+ N_A_515_297#_c_392_n N_A_515_297#_c_403_n N_A_515_297#_c_389_n
+ N_A_515_297#_c_411_n N_A_515_297#_c_390_n N_A_515_297#_c_391_n
+ N_A_515_297#_c_415_n PM_SKY130_FD_SC_HDLL__O22AI_2%A_515_297#
x_PM_SKY130_FD_SC_HDLL__O22AI_2%A_27_47# N_A_27_47#_M1006_s N_A_27_47#_M1013_s
+ N_A_27_47#_M1012_d N_A_27_47#_M1009_d N_A_27_47#_M1014_s N_A_27_47#_c_427_n
+ N_A_27_47#_c_428_n N_A_27_47#_c_436_n N_A_27_47#_c_442_n N_A_27_47#_c_429_n
+ N_A_27_47#_c_430_n N_A_27_47#_c_450_n N_A_27_47#_c_431_n N_A_27_47#_c_432_n
+ N_A_27_47#_c_433_n PM_SKY130_FD_SC_HDLL__O22AI_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O22AI_2%VGND N_VGND_M1002_s N_VGND_M1004_d
+ N_VGND_c_502_n N_VGND_c_503_n N_VGND_c_504_n N_VGND_c_505_n N_VGND_c_506_n
+ N_VGND_c_507_n VGND N_VGND_c_508_n N_VGND_c_509_n
+ PM_SKY130_FD_SC_HDLL__O22AI_2%VGND
cc_1 VNB N_B1_c_66_n 0.02229f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_B1_c_67_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_3 VNB N_B1_c_68_n 0.0150426f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_4 VNB N_B1_c_69_n 0.0426817f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_5 VNB N_B2_c_104_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B2_c_105_n 0.0204783f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_7 VNB N_B2_c_106_n 0.00625032f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_8 VNB N_B2_c_107_n 0.0402394f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_9 VNB N_A2_c_145_n 0.0202392f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_10 VNB N_A2_c_146_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_11 VNB N_A2_c_147_n 0.00446114f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_12 VNB N_A2_c_148_n 0.0398469f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_13 VNB N_A1_c_196_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_14 VNB N_A1_c_197_n 0.0223965f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_15 VNB A1 0.0123277f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_16 VNB N_A1_c_199_n 0.0426817f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_17 VNB N_VPWR_c_271_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_325_n 0.014401f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_19 VNB N_Y_c_326_n 0.0108356f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.18
cc_20 VNB N_A_27_47#_c_427_n 0.0075557f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_21 VNB N_A_27_47#_c_428_n 0.0212442f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_22 VNB N_A_27_47#_c_429_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_430_n 6.74925e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_431_n 0.0153158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_432_n 0.0187437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_433_n 0.00384559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_502_n 0.00464797f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_28 VNB N_VGND_c_503_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_29 VNB N_VGND_c_504_n 0.077256f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_30 VNB N_VGND_c_505_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.202
cc_31 VNB N_VGND_c_506_n 0.0180705f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_32 VNB N_VGND_c_507_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_33 VNB N_VGND_c_508_n 0.024694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_509_n 0.266034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VPB N_B1_c_70_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_36 VPB N_B1_c_71_n 0.0161059f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_37 VPB N_B1_c_69_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_38 VPB N_B2_c_108_n 0.0164196f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_39 VPB N_B2_c_109_n 0.0193324f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_40 VPB N_B2_c_107_n 0.0212133f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_41 VPB N_A2_c_149_n 0.0192267f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_42 VPB N_A2_c_150_n 0.0164192f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_43 VPB N_A2_c_148_n 0.0208791f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_44 VPB N_A1_c_200_n 0.0161059f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_45 VPB N_A1_c_201_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_46 VPB N_A1_c_199_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_47 VPB N_A_27_297#_c_237_n 0.00403131f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_48 VPB N_A_27_297#_c_238_n 0.00199216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_297#_c_239_n 0.00394856f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_50 VPB N_VPWR_c_272_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_51 VPB N_VPWR_c_273_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_52 VPB N_VPWR_c_274_n 0.0765778f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_53 VPB N_VPWR_c_275_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_54 VPB N_VPWR_c_276_n 0.0253799f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_271_n 0.0660401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_278_n 0.0244347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_Y_c_326_n 0.00432817f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.18
cc_58 VPB N_Y_c_328_n 0.00655386f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_59 VPB N_Y_c_329_n 0.00188018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_Y_c_330_n 0.00901475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_Y_c_331_n 0.00811829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_Y_c_332_n 0.00188018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_515_297#_c_389_n 0.00394549f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_64 VPB N_A_515_297#_c_390_n 0.00199216f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_65 VPB N_A_515_297#_c_391_n 0.0047508f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_66 N_B1_c_67_n N_B2_c_104_n 0.0247747f $X=1.01 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_67 N_B1_c_71_n N_B2_c_108_n 0.00966468f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_68 N_B1_c_68_n N_B2_c_106_n 0.0159646f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_69 N_B1_c_69_n N_B2_c_106_n 7.75592e-19 $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_70 N_B1_c_68_n N_B2_c_107_n 0.00103982f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_71 N_B1_c_69_n N_B2_c_107_n 0.0247747f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_72 N_B1_c_68_n N_A_27_297#_c_237_n 0.0175673f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_73 N_B1_c_70_n N_A_27_297#_c_238_n 0.0158351f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_74 N_B1_c_71_n N_A_27_297#_c_238_n 0.0155666f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_75 N_B1_c_68_n N_A_27_297#_c_238_n 0.0487774f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B1_c_69_n N_A_27_297#_c_238_n 0.00789593f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_77 N_B1_c_68_n N_A_27_297#_c_239_n 0.00171388f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B1_c_70_n N_VPWR_c_272_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_79 N_B1_c_71_n N_VPWR_c_272_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_80 N_B1_c_71_n N_VPWR_c_274_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_81 N_B1_c_70_n N_VPWR_c_271_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B1_c_71_n N_VPWR_c_271_n 0.0124344f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B1_c_70_n N_VPWR_c_278_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B1_c_66_n N_Y_c_325_n 0.0039356f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B1_c_67_n N_Y_c_325_n 0.0109542f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_86 N_B1_c_68_n N_Y_c_325_n 0.0429922f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B1_c_69_n N_Y_c_325_n 0.0047334f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_88 N_B1_c_66_n N_A_27_47#_c_428_n 4.6346e-19 $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B1_c_68_n N_A_27_47#_c_428_n 0.0139112f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B1_c_66_n N_A_27_47#_c_436_n 0.0101308f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B1_c_67_n N_A_27_47#_c_436_n 0.00851183f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_92 N_B1_c_68_n N_A_27_47#_c_436_n 0.00371054f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B1_c_66_n N_VGND_c_504_n 0.00368123f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B1_c_67_n N_VGND_c_504_n 0.00368123f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B1_c_66_n N_VGND_c_509_n 0.00647085f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B1_c_67_n N_VGND_c_509_n 0.00552518f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B2_c_108_n N_A_27_297#_c_239_n 2.98195e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B2_c_106_n N_A_27_297#_c_239_n 0.00164027f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B2_c_108_n N_A_27_297#_c_248_n 0.0143578f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B2_c_109_n N_A_27_297#_c_248_n 0.01161f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B2_c_108_n N_VPWR_c_274_n 0.00429453f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B2_c_109_n N_VPWR_c_274_n 0.00429453f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B2_c_108_n N_VPWR_c_271_n 0.00609021f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B2_c_109_n N_VPWR_c_271_n 0.00734734f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B2_c_104_n N_Y_c_325_n 0.0109542f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B2_c_105_n N_Y_c_325_n 0.0140712f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B2_c_106_n N_Y_c_325_n 0.0592259f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_108 N_B2_c_107_n N_Y_c_325_n 0.0047334f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_109 N_B2_c_109_n N_Y_c_326_n 9.79927e-19 $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_110 N_B2_c_105_n N_Y_c_326_n 0.00529891f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B2_c_106_n N_Y_c_326_n 0.0120878f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B2_c_107_n N_Y_c_326_n 0.00529466f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_113 N_B2_c_108_n N_Y_c_329_n 6.32035e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B2_c_106_n N_Y_c_329_n 0.020385f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_115 N_B2_c_107_n N_Y_c_329_n 0.00642616f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_116 N_B2_c_109_n N_Y_c_330_n 0.0153517f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_117 N_B2_c_106_n N_Y_c_330_n 0.0222091f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_118 N_B2_c_107_n N_Y_c_330_n 8.96166e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_119 N_B2_c_104_n N_A_27_47#_c_436_n 0.00851183f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B2_c_105_n N_A_27_47#_c_436_n 0.00851183f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B2_c_104_n N_VGND_c_504_n 0.00368123f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B2_c_105_n N_VGND_c_504_n 0.00368123f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B2_c_104_n N_VGND_c_509_n 0.00552518f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B2_c_105_n N_VGND_c_509_n 0.00682404f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A2_c_146_n N_A1_c_196_n 0.0175389f $X=3.45 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_126 N_A2_c_150_n N_A1_c_200_n 0.00966468f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A2_c_147_n A1 0.0160335f $X=3.39 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A2_c_148_n A1 0.00103982f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_129 N_A2_c_147_n N_A1_c_199_n 7.75592e-19 $X=3.39 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A2_c_148_n N_A1_c_199_n 0.0175389f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_131 N_A2_c_149_n N_VPWR_c_274_n 0.00429453f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A2_c_150_n N_VPWR_c_274_n 0.00429453f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A2_c_149_n N_VPWR_c_271_n 0.00734734f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A2_c_150_n N_VPWR_c_271_n 0.00609021f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A2_c_145_n N_Y_c_325_n 0.0018815f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A2_c_145_n N_Y_c_326_n 0.00634182f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A2_c_149_n N_Y_c_326_n 0.0011724f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A2_c_147_n N_Y_c_326_n 0.0159001f $X=3.39 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A2_c_148_n N_Y_c_326_n 0.00638916f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_140 N_A2_c_149_n N_Y_c_328_n 0.0153517f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A2_c_147_n N_Y_c_328_n 0.0160833f $X=3.39 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A2_c_148_n N_Y_c_328_n 8.96166e-19 $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_143 N_A2_c_150_n N_Y_c_332_n 6.32035e-19 $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A2_c_147_n N_Y_c_332_n 0.020385f $X=3.39 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A2_c_148_n N_Y_c_332_n 0.00642616f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_146 N_A2_c_149_n N_A_515_297#_c_392_n 0.01161f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A2_c_150_n N_A_515_297#_c_392_n 0.0143578f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A2_c_150_n N_A_515_297#_c_389_n 2.98195e-19 $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_149 N_A2_c_147_n N_A_515_297#_c_389_n 0.00164027f $X=3.39 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_c_145_n N_A_27_47#_c_436_n 0.00431104f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A2_c_145_n N_A_27_47#_c_442_n 0.00753478f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A2_c_146_n N_A_27_47#_c_442_n 5.58349e-19 $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A2_c_145_n N_A_27_47#_c_429_n 0.00370881f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A2_c_146_n N_A_27_47#_c_429_n 0.00922411f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A2_c_147_n N_A_27_47#_c_429_n 0.0364875f $X=3.39 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A2_c_148_n N_A_27_47#_c_429_n 0.00468948f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_157 N_A2_c_145_n N_A_27_47#_c_430_n 0.00673692f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A2_c_147_n N_A_27_47#_c_430_n 0.0116023f $X=3.39 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_c_145_n N_A_27_47#_c_450_n 5.79895e-19 $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_c_146_n N_A_27_47#_c_450_n 0.00643512f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A2_c_146_n N_A_27_47#_c_433_n 0.00112787f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_c_147_n N_A_27_47#_c_433_n 0.00485548f $X=3.39 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A2_c_145_n N_VGND_c_502_n 0.00550862f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_146_n N_VGND_c_502_n 0.00283206f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A2_c_145_n N_VGND_c_504_n 0.00377246f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A2_c_146_n N_VGND_c_506_n 0.00423334f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A2_c_145_n N_VGND_c_509_n 0.00693186f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A2_c_146_n N_VGND_c_509_n 0.00598581f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A1_c_200_n N_VPWR_c_273_n 0.00300743f $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A1_c_201_n N_VPWR_c_273_n 0.00300743f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A1_c_200_n N_VPWR_c_274_n 0.00702461f $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A1_c_201_n N_VPWR_c_276_n 0.00702461f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A1_c_200_n N_VPWR_c_271_n 0.0124344f $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A1_c_201_n N_VPWR_c_271_n 0.0134606f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_175 A1 N_A_515_297#_c_389_n 0.00171388f $X=4.2 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A1_c_200_n N_A_515_297#_c_390_n 0.0155666f $X=3.895 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A1_c_201_n N_A_515_297#_c_390_n 0.0158351f $X=4.365 $Y=1.41 $X2=0 $Y2=0
cc_178 A1 N_A_515_297#_c_390_n 0.0487774f $X=4.2 $Y=1.105 $X2=0 $Y2=0
cc_179 N_A1_c_199_n N_A_515_297#_c_390_n 0.00789593f $X=4.365 $Y=1.202 $X2=0
+ $Y2=0
cc_180 A1 N_A_515_297#_c_391_n 0.00771248f $X=4.2 $Y=1.105 $X2=0 $Y2=0
cc_181 N_A1_c_196_n N_A_27_47#_c_450_n 0.00693563f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_c_197_n N_A_27_47#_c_450_n 5.34901e-19 $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A1_c_196_n N_A_27_47#_c_431_n 0.00929182f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A1_c_197_n N_A_27_47#_c_431_n 0.00936658f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_185 A1 N_A_27_47#_c_431_n 0.05478f $X=4.2 $Y=1.105 $X2=0 $Y2=0
cc_186 N_A1_c_199_n N_A_27_47#_c_431_n 0.00468948f $X=4.365 $Y=1.202 $X2=0 $Y2=0
cc_187 N_A1_c_196_n N_A_27_47#_c_432_n 5.69266e-19 $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_197_n N_A_27_47#_c_432_n 0.00857123f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_196_n N_A_27_47#_c_433_n 0.00112787f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_190 A1 N_A_27_47#_c_433_n 0.00487201f $X=4.2 $Y=1.105 $X2=0 $Y2=0
cc_191 N_A1_c_196_n N_VGND_c_503_n 0.00385467f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A1_c_197_n N_VGND_c_503_n 0.00365402f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A1_c_196_n N_VGND_c_506_n 0.00423334f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A1_c_197_n N_VGND_c_508_n 0.00396605f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A1_c_196_n N_VGND_c_509_n 0.00610858f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_197_n N_VGND_c_509_n 0.00690174f $X=4.39 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_27_297#_c_238_n N_VPWR_M1001_d 0.00187091f $X=1.095 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_198 N_A_27_297#_c_238_n N_VPWR_c_272_n 0.0143191f $X=1.095 $Y=1.54 $X2=0
+ $Y2=0
cc_199 N_A_27_297#_c_252_p N_VPWR_c_274_n 0.015002f $X=1.22 $Y=2.295 $X2=0 $Y2=0
cc_200 N_A_27_297#_c_248_n N_VPWR_c_274_n 0.0549564f $X=2.035 $Y=2.38 $X2=0
+ $Y2=0
cc_201 N_A_27_297#_M1001_s N_VPWR_c_271_n 0.00358889f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_202 N_A_27_297#_M1011_s N_VPWR_c_271_n 0.00297222f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_203 N_A_27_297#_M1005_d N_VPWR_c_271_n 0.00303346f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_204 N_A_27_297#_c_257_p N_VPWR_c_271_n 0.00974347f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_205 N_A_27_297#_c_252_p N_VPWR_c_271_n 0.00962794f $X=1.22 $Y=2.295 $X2=0
+ $Y2=0
cc_206 N_A_27_297#_c_248_n N_VPWR_c_271_n 0.0335386f $X=2.035 $Y=2.38 $X2=0
+ $Y2=0
cc_207 N_A_27_297#_c_257_p N_VPWR_c_278_n 0.0165369f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_208 N_A_27_297#_c_248_n N_Y_M1003_s 0.00352392f $X=2.035 $Y=2.38 $X2=0 $Y2=0
cc_209 N_A_27_297#_c_239_n N_Y_c_325_n 0.00806986f $X=1.22 $Y=1.625 $X2=0 $Y2=0
cc_210 N_A_27_297#_c_239_n N_Y_c_329_n 0.00226124f $X=1.22 $Y=1.625 $X2=0 $Y2=0
cc_211 N_A_27_297#_c_248_n N_Y_c_329_n 0.0134104f $X=2.035 $Y=2.38 $X2=0 $Y2=0
cc_212 N_A_27_297#_M1005_d N_Y_c_330_n 0.00391072f $X=2.015 $Y=1.485 $X2=0 $Y2=0
cc_213 N_A_27_297#_c_248_n N_Y_c_330_n 0.00387236f $X=2.035 $Y=2.38 $X2=0 $Y2=0
cc_214 N_A_27_297#_c_267_p N_Y_c_330_n 0.0172937f $X=2.16 $Y=1.96 $X2=0 $Y2=0
cc_215 N_A_27_297#_c_267_p N_A_515_297#_c_402_n 0.0246907f $X=2.16 $Y=1.96 $X2=0
+ $Y2=0
cc_216 N_A_27_297#_c_248_n N_A_515_297#_c_403_n 0.00981548f $X=2.035 $Y=2.38
+ $X2=0 $Y2=0
cc_217 N_A_27_297#_c_237_n N_A_27_47#_c_428_n 0.00204459f $X=0.277 $Y=1.625
+ $X2=0 $Y2=0
cc_218 N_VPWR_c_271_n N_Y_M1003_s 0.00232895f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_c_271_n N_Y_M1000_d 0.00232895f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_c_271_n N_A_515_297#_M1000_s 0.00303346f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_221 N_VPWR_c_271_n N_A_515_297#_M1015_s 0.00297222f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_271_n N_A_515_297#_M1010_d 0.00358889f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_274_n N_A_515_297#_c_392_n 0.0386815f $X=4.005 $Y=2.72 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_271_n N_A_515_297#_c_392_n 0.0239144f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_274_n N_A_515_297#_c_403_n 0.0162749f $X=4.005 $Y=2.72 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_271_n N_A_515_297#_c_403_n 0.00962421f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_274_n N_A_515_297#_c_411_n 0.015002f $X=4.005 $Y=2.72 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_271_n N_A_515_297#_c_411_n 0.00962794f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_229 N_VPWR_M1008_s N_A_515_297#_c_390_n 0.00187091f $X=3.985 $Y=1.485 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_273_n N_A_515_297#_c_390_n 0.0143191f $X=4.13 $Y=1.96 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_276_n N_A_515_297#_c_415_n 0.0165369f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_271_n N_A_515_297#_c_415_n 0.00974347f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_233 N_Y_c_328_n N_A_515_297#_M1000_s 0.00202519f $X=3.065 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_234 N_Y_c_331_n N_A_515_297#_M1000_s 0.002032f $X=2.525 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_235 N_Y_c_328_n N_A_515_297#_c_402_n 0.0132598f $X=3.065 $Y=1.535 $X2=0 $Y2=0
cc_236 N_Y_c_331_n N_A_515_297#_c_402_n 0.00441308f $X=2.525 $Y=1.535 $X2=0
+ $Y2=0
cc_237 N_Y_M1000_d N_A_515_297#_c_392_n 0.00352392f $X=3.045 $Y=1.485 $X2=0
+ $Y2=0
cc_238 N_Y_c_328_n N_A_515_297#_c_392_n 0.00387236f $X=3.065 $Y=1.535 $X2=0
+ $Y2=0
cc_239 N_Y_c_332_n N_A_515_297#_c_392_n 0.0134104f $X=3.19 $Y=1.62 $X2=0 $Y2=0
cc_240 N_Y_c_332_n N_A_515_297#_c_389_n 0.00226124f $X=3.19 $Y=1.62 $X2=0 $Y2=0
cc_241 N_Y_c_325_n N_A_27_47#_M1013_s 0.00162317f $X=2.405 $Y=0.775 $X2=0 $Y2=0
cc_242 N_Y_c_325_n N_A_27_47#_M1012_d 0.0138543f $X=2.405 $Y=0.775 $X2=0 $Y2=0
cc_243 N_Y_c_325_n N_A_27_47#_c_428_n 0.0115996f $X=2.405 $Y=0.775 $X2=0 $Y2=0
cc_244 N_Y_M1006_d N_A_27_47#_c_436_n 0.00527949f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_245 N_Y_M1007_s N_A_27_47#_c_436_n 0.00527949f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_246 N_Y_c_325_n N_A_27_47#_c_436_n 0.120686f $X=2.405 $Y=0.775 $X2=0 $Y2=0
cc_247 N_Y_c_325_n N_A_27_47#_c_430_n 0.00903954f $X=2.405 $Y=0.775 $X2=0 $Y2=0
cc_248 N_Y_c_328_n N_A_27_47#_c_430_n 7.51328e-19 $X=3.065 $Y=1.535 $X2=0 $Y2=0
cc_249 N_Y_M1006_d N_VGND_c_509_n 0.00301822f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_250 N_Y_M1007_s N_VGND_c_509_n 0.00301822f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_251 N_A_515_297#_c_391_n N_A_27_47#_c_431_n 0.0067876f $X=4.602 $Y=1.625
+ $X2=0 $Y2=0
cc_252 N_A_515_297#_c_389_n N_A_27_47#_c_433_n 0.00863876f $X=3.66 $Y=1.625
+ $X2=0 $Y2=0
cc_253 N_A_27_47#_c_429_n N_VGND_M1002_s 0.00356038f $X=3.495 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_254 N_A_27_47#_c_431_n N_VGND_M1004_d 0.00348805f $X=4.385 $Y=0.815 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_436_n N_VGND_c_502_n 0.0133618f $X=2.815 $Y=0.39 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_442_n N_VGND_c_502_n 0.00558251f $X=2.9 $Y=0.725 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_429_n N_VGND_c_502_n 0.0127273f $X=3.495 $Y=0.815 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_450_n N_VGND_c_503_n 0.0181628f $X=3.66 $Y=0.39 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_431_n N_VGND_c_503_n 0.0131987f $X=4.385 $Y=0.815 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_432_n N_VGND_c_503_n 0.0223967f $X=4.6 $Y=0.39 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_427_n N_VGND_c_504_n 0.0143679f $X=0.227 $Y=0.475 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_436_n N_VGND_c_504_n 0.114807f $X=2.815 $Y=0.39 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_429_n N_VGND_c_504_n 0.00204938f $X=3.495 $Y=0.815 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_429_n N_VGND_c_506_n 0.00198695f $X=3.495 $Y=0.815 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_450_n N_VGND_c_506_n 0.0188551f $X=3.66 $Y=0.39 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_431_n N_VGND_c_506_n 0.00266636f $X=4.385 $Y=0.815 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_431_n N_VGND_c_508_n 0.00199443f $X=4.385 $Y=0.815 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_432_n N_VGND_c_508_n 0.024373f $X=4.6 $Y=0.39 $X2=0 $Y2=0
cc_269 N_A_27_47#_M1006_s N_VGND_c_509_n 0.00229179f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_M1013_s N_VGND_c_509_n 0.00218617f $X=1.085 $Y=0.235 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1012_d N_VGND_c_509_n 0.00683313f $X=2.025 $Y=0.235 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1009_d N_VGND_c_509_n 0.00215201f $X=3.525 $Y=0.235 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1014_s N_VGND_c_509_n 0.00209319f $X=4.465 $Y=0.235 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_427_n N_VGND_c_509_n 0.0102867f $X=0.227 $Y=0.475 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_436_n N_VGND_c_509_n 0.0910547f $X=2.815 $Y=0.39 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_429_n N_VGND_c_509_n 0.00893695f $X=3.495 $Y=0.815 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_450_n N_VGND_c_509_n 0.0122069f $X=3.66 $Y=0.39 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_431_n N_VGND_c_509_n 0.0100158f $X=4.385 $Y=0.815 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_432_n N_VGND_c_509_n 0.0141066f $X=4.6 $Y=0.39 $X2=0 $Y2=0
