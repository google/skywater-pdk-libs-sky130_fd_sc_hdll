* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand4_4 A B C D VGND VNB VPB VPWR Y
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_485_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_883_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_485_47# B a_883_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_883_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_485_47# B a_883_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_27_47# C a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_27_47# C a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_883_47# B a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 Y A a_883_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 a_883_47# B a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 Y A a_883_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 a_485_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
