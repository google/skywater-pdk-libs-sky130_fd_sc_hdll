* File: sky130_fd_sc_hdll__and3_1.pex.spice
* Created: Wed Sep  2 08:22:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND3_1%A 1 3 4 6 7
r26 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=0.93 $X2=0.26 $Y2=0.93
r27 4 10 43.8307 $w=4.03e-07 $l=2.68328e-07 $layer=POLY_cond $X=0.52 $Y=0.73
+ $X2=0.36 $Y2=0.93
r28 4 6 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r29 1 10 74.1653 $w=4.03e-07 $l=5.58435e-07 $layer=POLY_cond $X=0.495 $Y=1.425
+ $X2=0.36 $Y2=0.93
r30 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.425
+ $X2=0.495 $Y2=1.71
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_1%B 2 4 7 10 11 20
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=2.295
+ $X2=1 $Y2=2.295
r36 11 20 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=1.145 $Y=2.295
+ $X2=1.15 $Y2=2.295
r37 11 15 4.91483 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=1.145 $Y=2.295
+ $X2=1 $Y2=2.295
r38 9 10 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.97 $Y=1.275
+ $X2=0.97 $Y2=1.425
r39 7 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=0.99 $Y=0.445 $X2=0.99
+ $Y2=1.275
r40 4 10 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.965 $Y=1.71
+ $X2=0.965 $Y2=1.425
r41 2 14 47.2445 $w=2.96e-07 $l=2.73359e-07 $layer=POLY_cond $X=0.965 $Y=2.05
+ $X2=1.025 $Y2=2.295
r42 2 4 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.965 $Y=2.05
+ $X2=0.965 $Y2=1.71
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_1%C 1 3 6 8
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.575
+ $Y=1.115 $X2=1.575 $Y2=1.115
r32 8 12 8.25398 $w=3.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.575 $Y=0.85
+ $X2=1.575 $Y2=1.115
r33 4 11 42.1211 $w=2.82e-07 $l=2.21416e-07 $layer=POLY_cond $X=1.675 $Y=0.93
+ $X2=1.595 $Y2=1.115
r34 4 6 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.675 $Y=0.93
+ $X2=1.675 $Y2=0.445
r35 1 11 59.2695 $w=2.82e-07 $l=3.36378e-07 $layer=POLY_cond $X=1.65 $Y=1.425
+ $X2=1.595 $Y2=1.115
r36 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.65 $Y=1.425
+ $X2=1.65 $Y2=1.71
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_1%A_27_47# 1 2 3 10 12 13 15 16 22 24 25 27
+ 28 29 32
r73 35 37 8.87273 $w=3.85e-07 $l=2.8e-07 $layer=LI1_cond $X=0.965 $Y=1.537
+ $X2=1.245 $Y2=1.537
r74 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.185
+ $Y=1.16 $X2=2.185 $Y2=1.16
r75 30 32 10.5223 $w=2.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.155 $Y=1.37
+ $X2=2.155 $Y2=1.16
r76 29 37 4.87876 $w=5.15e-07 $l=2.12283e-07 $layer=LI1_cond $X=1.417 $Y=1.627
+ $X2=1.245 $Y2=1.537
r77 28 30 4.96033 $w=6.15e-07 $l=3.09199e-07 $layer=LI1_cond $X=2.04 $Y=1.627
+ $X2=2.155 $Y2=1.37
r78 28 29 14.4691 $w=5.13e-07 $l=6.23e-07 $layer=LI1_cond $X=2.04 $Y=1.627
+ $X2=1.417 $Y2=1.627
r79 27 35 4.01183 $w=2.2e-07 $l=3.47e-07 $layer=LI1_cond $X=0.965 $Y=1.19
+ $X2=0.965 $Y2=1.537
r80 26 27 37.9782 $w=2.18e-07 $l=7.25e-07 $layer=LI1_cond $X=0.965 $Y=0.465
+ $X2=0.965 $Y2=1.19
r81 24 35 7.34957 $w=3.85e-07 $l=3.12192e-07 $layer=LI1_cond $X=0.855 $Y=1.275
+ $X2=0.965 $Y2=1.537
r82 24 25 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.855 $Y=1.275
+ $X2=0.345 $Y2=1.275
r83 20 25 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=1.36
+ $X2=0.345 $Y2=1.275
r84 20 22 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=0.215 $Y=1.36
+ $X2=0.215 $Y2=1.645
r85 16 26 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.855 $Y=0.38
+ $X2=0.965 $Y2=0.465
r86 16 18 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.855 $Y=0.38
+ $X2=0.26 $Y2=0.38
r87 13 33 38.7444 $w=2.79e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.2 $Y2=1.16
r88 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.275 $Y2=0.56
r89 10 33 49.2447 $w=2.79e-07 $l=2.73861e-07 $layer=POLY_cond $X=2.25 $Y=1.41
+ $X2=2.2 $Y2=1.16
r90 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.25 $Y=1.41
+ $X2=2.25 $Y2=1.985
r91 3 37 600 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.5 $X2=1.245 $Y2=1.7
r92 2 22 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.5 $X2=0.26 $Y2=1.645
r93 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_1%VPWR 1 2 9 11 13 20 21 26 31
r31 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 26 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r33 24 26 18.9028 $w=5.97e-07 $l=1.05707e-06 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.447 $Y2=2.72
r34 21 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r35 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 18 31 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.037 $Y2=2.72
r37 18 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.53 $Y2=2.72
r38 17 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r39 17 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 16 26 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=0.74 $Y2=2.72
r41 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r42 13 31 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.91 $Y=2.72
+ $X2=2.037 $Y2=2.72
r43 13 16 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.91 $Y=2.72 $X2=1.61
+ $Y2=2.72
r44 11 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 11 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r46 7 31 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.037 $Y=2.635
+ $X2=2.037 $Y2=2.72
r47 7 9 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=2.037 $Y=2.635
+ $X2=2.037 $Y2=2.34
r48 2 9 600 $w=1.7e-07 $l=9.67781e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.5 $X2=2.015 $Y2=2.34
r49 1 24 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.5 $X2=0.73 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_1%X 1 2 9 10 12 13 14 22
r16 14 22 11.734 $w=2.73e-07 $l=2.8e-07 $layer=LI1_cond $X=2.522 $Y=2.21
+ $X2=2.522 $Y2=1.93
r17 11 13 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=2.53 $Y=0.605
+ $X2=2.53 $Y2=0.51
r18 11 12 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.53 $Y=0.605
+ $X2=2.53 $Y2=0.735
r19 10 12 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.575 $Y=1.765
+ $X2=2.575 $Y2=0.735
r20 9 22 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=2.522 $Y=1.902
+ $X2=2.522 $Y2=1.93
r21 9 10 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.522 $Y=1.902
+ $X2=2.522 $Y2=1.765
r22 2 22 300 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_PDIFF $count=2 $X=2.34
+ $Y=1.485 $X2=2.485 $Y2=1.93
r23 1 13 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.235 $X2=2.485 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_1%VGND 1 6 9 10 11 21 22
r27 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r28 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r29 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r30 14 18 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r31 11 19 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r32 11 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r33 9 18 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.61
+ $Y2=0
r34 9 10 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.015
+ $Y2=0
r35 8 21 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=2.53
+ $Y2=0
r36 8 10 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=0 $X2=2.015
+ $Y2=0
r37 4 10 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0
r38 4 6 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0.46
r39 1 6 182 $w=1.7e-07 $l=3.60347e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.235 $X2=2.015 $Y2=0.46
.ends

