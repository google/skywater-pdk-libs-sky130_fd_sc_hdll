* File: sky130_fd_sc_hdll__and4bb_1.pxi.spice
* Created: Wed Sep  2 08:23:34 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%A_N N_A_N_M1008_g N_A_N_c_99_n N_A_N_M1011_g
+ A_N N_A_N_c_100_n PM_SKY130_FD_SC_HDLL__AND4BB_1%A_N
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%B_N N_B_N_c_128_n N_B_N_c_134_n N_B_N_M1004_g
+ N_B_N_M1007_g N_B_N_c_130_n N_B_N_c_131_n B_N
+ PM_SKY130_FD_SC_HDLL__AND4BB_1%B_N
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1011_s
+ N_A_27_47#_c_176_n N_A_27_47#_M1012_g N_A_27_47#_M1000_g N_A_27_47#_c_178_n
+ N_A_27_47#_c_179_n N_A_27_47#_c_171_n N_A_27_47#_c_180_n N_A_27_47#_c_172_n
+ N_A_27_47#_c_182_n N_A_27_47#_c_173_n N_A_27_47#_c_174_n N_A_27_47#_c_184_n
+ N_A_27_47#_c_175_n PM_SKY130_FD_SC_HDLL__AND4BB_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%A_225_413# N_A_225_413#_M1007_d
+ N_A_225_413#_M1004_d N_A_225_413#_M1003_g N_A_225_413#_c_263_n
+ N_A_225_413#_c_264_n N_A_225_413#_M1005_g N_A_225_413#_c_283_n
+ N_A_225_413#_c_265_n N_A_225_413#_c_266_n N_A_225_413#_c_255_n
+ N_A_225_413#_c_256_n N_A_225_413#_c_257_n N_A_225_413#_c_258_n
+ N_A_225_413#_c_269_n N_A_225_413#_c_259_n N_A_225_413#_c_260_n
+ N_A_225_413#_c_261_n N_A_225_413#_c_262_n
+ PM_SKY130_FD_SC_HDLL__AND4BB_1%A_225_413#
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%C N_C_M1001_g N_C_c_359_n N_C_c_360_n
+ N_C_M1002_g C C C C N_C_c_357_n N_C_c_358_n PM_SKY130_FD_SC_HDLL__AND4BB_1%C
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%D N_D_c_402_n N_D_c_403_n N_D_M1006_g
+ N_D_M1009_g D D D D N_D_c_400_n N_D_c_401_n PM_SKY130_FD_SC_HDLL__AND4BB_1%D
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%A_339_93# N_A_339_93#_M1000_s
+ N_A_339_93#_M1012_d N_A_339_93#_M1002_d N_A_339_93#_c_443_n
+ N_A_339_93#_M1010_g N_A_339_93#_c_444_n N_A_339_93#_M1013_g
+ N_A_339_93#_c_445_n N_A_339_93#_c_446_n N_A_339_93#_c_459_n
+ N_A_339_93#_c_450_n N_A_339_93#_c_481_n N_A_339_93#_c_451_n
+ N_A_339_93#_c_452_n N_A_339_93#_c_453_n N_A_339_93#_c_454_n
+ N_A_339_93#_c_447_n PM_SKY130_FD_SC_HDLL__AND4BB_1%A_339_93#
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%VPWR N_VPWR_M1011_d N_VPWR_M1012_s
+ N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n
+ N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n VPWR N_VPWR_c_539_n
+ N_VPWR_c_540_n N_VPWR_c_541_n N_VPWR_c_532_n N_VPWR_c_543_n N_VPWR_c_544_n
+ PM_SKY130_FD_SC_HDLL__AND4BB_1%VPWR
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%X N_X_M1013_d N_X_M1010_d X X X X X N_X_c_612_n
+ X X PM_SKY130_FD_SC_HDLL__AND4BB_1%X
x_PM_SKY130_FD_SC_HDLL__AND4BB_1%VGND N_VGND_M1008_d N_VGND_M1009_d
+ N_VGND_c_630_n N_VGND_c_631_n N_VGND_c_632_n VGND N_VGND_c_633_n
+ N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n
+ PM_SKY130_FD_SC_HDLL__AND4BB_1%VGND
cc_1 VNB N_A_N_M1008_g 0.0497384f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.445
cc_2 VNB N_B_N_c_128_n 0.00725872f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.445
cc_3 VNB N_B_N_M1007_g 0.0266123f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.76
cc_4 VNB N_B_N_c_130_n 0.0053045f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.745
cc_5 VNB N_B_N_c_131_n 0.0290221f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.745
cc_6 VNB B_N 0.00537982f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.845
cc_7 VNB N_A_27_47#_M1000_g 0.0527313f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.745
cc_8 VNB N_A_27_47#_c_171_n 0.0333864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_172_n 0.00963418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_173_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_174_n 9.40304e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_175_n 0.00201385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_225_413#_c_255_n 0.0117941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_225_413#_c_256_n 0.0217164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_225_413#_c_257_n 0.00892306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_225_413#_c_258_n 0.00117256f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_225_413#_c_259_n 0.001001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_225_413#_c_260_n 0.0270053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_225_413#_c_261_n 0.0181419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_225_413#_c_262_n 0.0277242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB C 0.00561886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_C_c_357_n 0.0210286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_C_c_358_n 0.0313368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB D 0.00458461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_D_c_400_n 0.0205545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_D_c_401_n 0.03233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_339_93#_c_443_n 0.0272592f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.745
cc_28 VNB N_A_339_93#_c_444_n 0.0203302f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.745
cc_29 VNB N_A_339_93#_c_445_n 0.00371172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_339_93#_c_446_n 0.00655544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_339_93#_c_447_n 0.0028761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_532_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB X 0.0233241f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.745
cc_34 VNB N_X_c_612_n 0.0170421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB X 0.00494099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_630_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_631_n 0.0725815f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.745
cc_38 VNB N_VGND_c_632_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.745
cc_39 VNB N_VGND_c_633_n 0.0169726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_634_n 0.0194457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_635_n 0.266255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_636_n 0.00916597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VPB N_A_N_M1008_g 0.0163349f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.445
cc_44 VPB N_A_N_c_99_n 0.0519782f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.99
cc_45 VPB N_A_N_c_100_n 0.00916721f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.745
cc_46 VPB N_B_N_c_128_n 0.0337516f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.445
cc_47 VPB N_B_N_c_134_n 0.0263129f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.445
cc_48 VPB N_A_27_47#_c_176_n 0.0190089f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=2.275
cc_49 VPB N_A_27_47#_M1000_g 0.0119488f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.745
cc_50 VPB N_A_27_47#_c_178_n 0.0547027f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_179_n 0.0269023f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.845
cc_52 VPB N_A_27_47#_c_180_n 0.032116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_172_n 0.0118901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_182_n 0.00509725f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_174_n 0.00705228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_184_n 0.0129899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_175_n 0.00522225f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_225_413#_c_263_n 0.0342985f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.745
cc_59 VPB N_A_225_413#_c_264_n 0.021613f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.745
cc_60 VPB N_A_225_413#_c_265_n 0.00791382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_225_413#_c_266_n 0.00439727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_225_413#_c_257_n 0.00184366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_225_413#_c_258_n 0.00224508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_225_413#_c_269_n 0.00243664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_225_413#_c_259_n 9.58049e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_225_413#_c_260_n 0.00471825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_C_c_359_n 0.0323379f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.99
cc_68 VPB N_C_c_360_n 0.0227211f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=2.275
cc_69 VPB C 0.00630188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_C_c_357_n 0.00317326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_D_c_402_n 0.0342198f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.445
cc_72 VPB N_D_c_403_n 0.0228233f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.445
cc_73 VPB D 0.00351196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_D_c_400_n 0.00309074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_339_93#_c_443_n 0.0310548f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.745
cc_76 VPB N_A_339_93#_c_446_n 0.0118067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_339_93#_c_450_n 0.0103802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_339_93#_c_451_n 0.00346224f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_339_93#_c_452_n 0.00226073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_339_93#_c_453_n 0.00236125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_339_93#_c_454_n 0.00573096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_339_93#_c_447_n 3.24692e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_533_n 0.00481032f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.845
cc_84 VPB N_VPWR_c_534_n 0.00285982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_535_n 0.0171603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_536_n 0.00513086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_537_n 0.0088967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_538_n 0.0140593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_539_n 0.0169726f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_540_n 0.0202037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_541_n 0.0168079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_532_n 0.0466503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_543_n 0.00548208f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_544_n 0.00513086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB X 0.0400932f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.76
cc_96 VPB X 0.00700168f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.745
cc_97 N_A_N_M1008_g N_B_N_c_128_n 0.0142989f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_N_c_99_n N_B_N_c_128_n 0.0198667f $X=0.555 $Y=1.99 $X2=0 $Y2=0
cc_99 N_A_N_c_100_n N_B_N_c_128_n 0.00543863f $X=0.59 $Y=1.745 $X2=0 $Y2=0
cc_100 N_A_N_c_99_n N_B_N_c_134_n 0.0151811f $X=0.555 $Y=1.99 $X2=0 $Y2=0
cc_101 N_A_N_M1008_g N_B_N_M1007_g 0.0133634f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A_N_M1008_g N_B_N_c_131_n 0.0163781f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_103 N_A_N_M1008_g B_N 0.0117317f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_N_M1008_g N_A_27_47#_c_171_n 0.0179224f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_N_M1008_g N_A_27_47#_c_180_n 0.00570754f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_N_c_99_n N_A_27_47#_c_180_n 0.0081859f $X=0.555 $Y=1.99 $X2=0 $Y2=0
cc_107 N_A_N_c_100_n N_A_27_47#_c_180_n 0.0265113f $X=0.59 $Y=1.745 $X2=0 $Y2=0
cc_108 N_A_N_M1008_g N_A_27_47#_c_172_n 0.0144243f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_N_c_99_n N_A_27_47#_c_172_n 0.00301157f $X=0.555 $Y=1.99 $X2=0 $Y2=0
cc_110 N_A_N_c_100_n N_A_27_47#_c_172_n 0.02923f $X=0.59 $Y=1.745 $X2=0 $Y2=0
cc_111 N_A_N_c_99_n N_A_27_47#_c_184_n 0.00925204f $X=0.555 $Y=1.99 $X2=0 $Y2=0
cc_112 N_A_N_M1008_g N_A_27_47#_c_175_n 7.40684e-19 $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_N_c_99_n N_A_27_47#_c_175_n 3.76438e-19 $X=0.555 $Y=1.99 $X2=0 $Y2=0
cc_114 N_A_N_c_100_n N_A_27_47#_c_175_n 0.00828295f $X=0.59 $Y=1.745 $X2=0 $Y2=0
cc_115 N_A_N_c_100_n N_A_225_413#_c_266_n 0.00216044f $X=0.59 $Y=1.745 $X2=0
+ $Y2=0
cc_116 N_A_N_c_99_n N_VPWR_c_539_n 0.00449985f $X=0.555 $Y=1.99 $X2=0 $Y2=0
cc_117 N_A_N_c_99_n N_VPWR_c_532_n 0.00526272f $X=0.555 $Y=1.99 $X2=0 $Y2=0
cc_118 N_A_N_c_100_n N_VPWR_c_532_n 0.00613174f $X=0.59 $Y=1.745 $X2=0 $Y2=0
cc_119 N_A_N_c_99_n N_VPWR_c_543_n 0.012042f $X=0.555 $Y=1.99 $X2=0 $Y2=0
cc_120 N_A_N_c_100_n N_VPWR_c_543_n 0.0100255f $X=0.59 $Y=1.745 $X2=0 $Y2=0
cc_121 N_A_N_M1008_g N_VGND_c_633_n 0.00468308f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_N_M1008_g N_VGND_c_635_n 0.00736021f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_123 N_A_N_M1008_g N_VGND_c_636_n 0.00907591f $X=0.53 $Y=0.445 $X2=0 $Y2=0
cc_124 N_B_N_c_128_n N_A_27_47#_c_178_n 0.0219544f $X=1.035 $Y=1.89 $X2=0 $Y2=0
cc_125 B_N N_A_27_47#_c_171_n 0.0182918f $X=0.525 $Y=0.765 $X2=0 $Y2=0
cc_126 N_B_N_c_128_n N_A_27_47#_c_172_n 0.00865462f $X=1.035 $Y=1.89 $X2=0 $Y2=0
cc_127 N_B_N_c_130_n N_A_27_47#_c_172_n 0.0164527f $X=1 $Y=1.03 $X2=0 $Y2=0
cc_128 N_B_N_c_131_n N_A_27_47#_c_172_n 0.0017253f $X=1 $Y=1.03 $X2=0 $Y2=0
cc_129 B_N N_A_27_47#_c_172_n 0.0200226f $X=0.525 $Y=0.765 $X2=0 $Y2=0
cc_130 N_B_N_c_128_n N_A_27_47#_c_175_n 0.0210969f $X=1.035 $Y=1.89 $X2=0 $Y2=0
cc_131 N_B_N_c_130_n N_A_27_47#_c_175_n 0.0112293f $X=1 $Y=1.03 $X2=0 $Y2=0
cc_132 N_B_N_c_134_n N_A_225_413#_c_266_n 0.00684819f $X=1.035 $Y=1.99 $X2=0
+ $Y2=0
cc_133 N_B_N_M1007_g N_A_225_413#_c_255_n 0.00417602f $X=1.06 $Y=0.445 $X2=0
+ $Y2=0
cc_134 N_B_N_c_130_n N_A_225_413#_c_255_n 0.0103273f $X=1 $Y=1.03 $X2=0 $Y2=0
cc_135 N_B_N_c_131_n N_A_225_413#_c_255_n 0.00488012f $X=1 $Y=1.03 $X2=0 $Y2=0
cc_136 B_N N_A_225_413#_c_255_n 0.00561822f $X=0.525 $Y=0.765 $X2=0 $Y2=0
cc_137 N_B_N_c_128_n N_A_225_413#_c_258_n 0.00255105f $X=1.035 $Y=1.89 $X2=0
+ $Y2=0
cc_138 N_B_N_c_128_n N_A_225_413#_c_269_n 0.00256293f $X=1.035 $Y=1.89 $X2=0
+ $Y2=0
cc_139 N_B_N_M1007_g N_A_225_413#_c_261_n 0.00507874f $X=1.06 $Y=0.445 $X2=0
+ $Y2=0
cc_140 N_B_N_c_134_n N_VPWR_c_533_n 0.00185679f $X=1.035 $Y=1.99 $X2=0 $Y2=0
cc_141 N_B_N_c_134_n N_VPWR_c_535_n 0.00684138f $X=1.035 $Y=1.99 $X2=0 $Y2=0
cc_142 N_B_N_c_134_n N_VPWR_c_532_n 0.0125562f $X=1.035 $Y=1.99 $X2=0 $Y2=0
cc_143 N_B_N_c_134_n N_VPWR_c_543_n 0.00685265f $X=1.035 $Y=1.99 $X2=0 $Y2=0
cc_144 N_B_N_M1007_g N_VGND_c_631_n 0.00585385f $X=1.06 $Y=0.445 $X2=0 $Y2=0
cc_145 N_B_N_M1007_g N_VGND_c_635_n 0.0120869f $X=1.06 $Y=0.445 $X2=0 $Y2=0
cc_146 N_B_N_c_131_n N_VGND_c_635_n 7.41941e-19 $X=1 $Y=1.03 $X2=0 $Y2=0
cc_147 B_N N_VGND_c_635_n 0.00262068f $X=0.525 $Y=0.765 $X2=0 $Y2=0
cc_148 N_B_N_M1007_g N_VGND_c_636_n 0.0032017f $X=1.06 $Y=0.445 $X2=0 $Y2=0
cc_149 N_B_N_c_130_n N_VGND_c_636_n 0.00564865f $X=1 $Y=1.03 $X2=0 $Y2=0
cc_150 N_B_N_c_131_n N_VGND_c_636_n 0.00177008f $X=1 $Y=1.03 $X2=0 $Y2=0
cc_151 B_N N_VGND_c_636_n 0.00881422f $X=0.525 $Y=0.765 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_179_n N_A_225_413#_c_263_n 0.0382486f $X=2.025 $Y=1.742
+ $X2=0 $Y2=0
cc_153 N_A_27_47#_c_176_n N_A_225_413#_c_264_n 0.0102171f $X=2.025 $Y=1.99 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_c_176_n N_A_225_413#_c_283_n 0.00275289f $X=2.025 $Y=1.99
+ $X2=0 $Y2=0
cc_155 N_A_27_47#_c_176_n N_A_225_413#_c_265_n 0.00442205f $X=2.025 $Y=1.99
+ $X2=0 $Y2=0
cc_156 N_A_27_47#_c_178_n N_A_225_413#_c_265_n 0.0115347f $X=1.925 $Y=1.66 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_179_n N_A_225_413#_c_265_n 0.00301619f $X=2.025 $Y=1.742
+ $X2=0 $Y2=0
cc_158 N_A_27_47#_c_182_n N_A_225_413#_c_265_n 0.0192719f $X=1.48 $Y=1.66 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_178_n N_A_225_413#_c_266_n 7.6408e-19 $X=1.925 $Y=1.66 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_182_n N_A_225_413#_c_266_n 0.0115073f $X=1.48 $Y=1.66 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_175_n N_A_225_413#_c_266_n 0.00618061f $X=1.125 $Y=1.37
+ $X2=0 $Y2=0
cc_162 N_A_27_47#_M1000_g N_A_225_413#_c_255_n 0.00548918f $X=2.05 $Y=0.675
+ $X2=0 $Y2=0
cc_163 N_A_27_47#_M1000_g N_A_225_413#_c_256_n 0.0112684f $X=2.05 $Y=0.675 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_M1000_g N_A_225_413#_c_257_n 0.00567735f $X=2.05 $Y=0.675
+ $X2=0 $Y2=0
cc_165 N_A_27_47#_c_178_n N_A_225_413#_c_257_n 0.00635877f $X=1.925 $Y=1.66
+ $X2=0 $Y2=0
cc_166 N_A_27_47#_c_182_n N_A_225_413#_c_257_n 0.00425338f $X=1.48 $Y=1.66 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_178_n N_A_225_413#_c_258_n 0.0043649f $X=1.925 $Y=1.66 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_182_n N_A_225_413#_c_258_n 0.0137147f $X=1.48 $Y=1.66 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_175_n N_A_225_413#_c_258_n 0.00976481f $X=1.125 $Y=1.37
+ $X2=0 $Y2=0
cc_170 N_A_27_47#_M1000_g N_A_225_413#_c_269_n 0.0023513f $X=2.05 $Y=0.675 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_178_n N_A_225_413#_c_269_n 0.0132593f $X=1.925 $Y=1.66 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_179_n N_A_225_413#_c_269_n 0.00825107f $X=2.025 $Y=1.742
+ $X2=0 $Y2=0
cc_173 N_A_27_47#_c_182_n N_A_225_413#_c_269_n 0.012273f $X=1.48 $Y=1.66 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_175_n N_A_225_413#_c_269_n 0.00529234f $X=1.125 $Y=1.37
+ $X2=0 $Y2=0
cc_175 N_A_27_47#_M1000_g N_A_225_413#_c_259_n 0.00129037f $X=2.05 $Y=0.675
+ $X2=0 $Y2=0
cc_176 N_A_27_47#_M1000_g N_A_225_413#_c_261_n 0.00587557f $X=2.05 $Y=0.675
+ $X2=0 $Y2=0
cc_177 N_A_27_47#_c_175_n N_A_225_413#_c_261_n 0.00193045f $X=1.125 $Y=1.37
+ $X2=0 $Y2=0
cc_178 N_A_27_47#_M1000_g N_A_225_413#_c_262_n 0.0382486f $X=2.05 $Y=0.675 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1000_g N_A_339_93#_c_445_n 0.0170762f $X=2.05 $Y=0.675 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_178_n N_A_339_93#_c_445_n 8.04243e-19 $X=1.925 $Y=1.66 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1000_g N_A_339_93#_c_446_n 0.00956499f $X=2.05 $Y=0.675 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_176_n N_A_339_93#_c_459_n 0.00410146f $X=2.025 $Y=1.99 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_176_n N_A_339_93#_c_453_n 7.4621e-19 $X=2.025 $Y=1.99 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_179_n N_A_339_93#_c_453_n 6.59561e-19 $X=2.025 $Y=1.742
+ $X2=0 $Y2=0
cc_185 N_A_27_47#_c_176_n N_VPWR_c_533_n 0.00794629f $X=2.025 $Y=1.99 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_178_n N_VPWR_c_533_n 7.38178e-19 $X=1.925 $Y=1.66 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_176_n N_VPWR_c_537_n 5.17995e-19 $X=2.025 $Y=1.99 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_176_n N_VPWR_c_538_n 0.00591615f $X=2.025 $Y=1.99 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_179_n N_VPWR_c_538_n 2.07025e-19 $X=2.025 $Y=1.742 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_184_n N_VPWR_c_539_n 0.0173041f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_191 N_A_27_47#_M1011_s N_VPWR_c_532_n 0.00570386f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_176_n N_VPWR_c_532_n 0.00942972f $X=2.025 $Y=1.99 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_179_n N_VPWR_c_532_n 2.58415e-19 $X=2.025 $Y=1.742 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_184_n N_VPWR_c_532_n 0.00982816f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_184_n N_VPWR_c_543_n 0.0128131f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_196 N_A_27_47#_M1000_g N_VGND_c_631_n 0.00357877f $X=2.05 $Y=0.675 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_173_n N_VGND_c_633_n 0.0173041f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_198 N_A_27_47#_M1008_s N_VGND_c_635_n 0.00636928f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_M1000_g N_VGND_c_635_n 0.00669482f $X=2.05 $Y=0.675 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_173_n N_VGND_c_635_n 0.00982816f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_173_n N_VGND_c_636_n 0.0128131f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_202 N_A_225_413#_c_263_n N_C_c_359_n 0.0128797f $X=2.505 $Y=1.89 $X2=0 $Y2=0
cc_203 N_A_225_413#_c_264_n N_C_c_360_n 0.023211f $X=2.505 $Y=1.99 $X2=0 $Y2=0
cc_204 N_A_225_413#_c_263_n C 0.00282404f $X=2.505 $Y=1.89 $X2=0 $Y2=0
cc_205 N_A_225_413#_c_256_n C 7.56833e-19 $X=2.495 $Y=0.34 $X2=0 $Y2=0
cc_206 N_A_225_413#_c_259_n C 0.0442317f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_225_413#_c_260_n C 0.00204344f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_225_413#_c_262_n C 7.91571e-19 $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_225_413#_c_259_n N_C_c_357_n 3.5305e-19 $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_225_413#_c_260_n N_C_c_357_n 0.0204839f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_225_413#_c_256_n N_C_c_358_n 0.00413197f $X=2.495 $Y=0.34 $X2=0 $Y2=0
cc_212 N_A_225_413#_c_259_n N_C_c_358_n 0.00178229f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_225_413#_c_262_n N_C_c_358_n 0.0280081f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_225_413#_c_256_n N_A_339_93#_c_445_n 0.0373229f $X=2.495 $Y=0.34
+ $X2=0 $Y2=0
cc_215 N_A_225_413#_c_257_n N_A_339_93#_c_445_n 0.0129212f $X=1.815 $Y=1.32
+ $X2=0 $Y2=0
cc_216 N_A_225_413#_c_259_n N_A_339_93#_c_445_n 0.0257339f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_217 N_A_225_413#_c_261_n N_A_339_93#_c_445_n 0.0276024f $X=1.385 $Y=0.34
+ $X2=0 $Y2=0
cc_218 N_A_225_413#_c_262_n N_A_339_93#_c_445_n 0.00246803f $X=2.56 $Y=0.995
+ $X2=0 $Y2=0
cc_219 N_A_225_413#_c_255_n N_A_339_93#_c_446_n 0.00995712f $X=1.5 $Y=1.235
+ $X2=0 $Y2=0
cc_220 N_A_225_413#_c_257_n N_A_339_93#_c_446_n 0.0133941f $X=1.815 $Y=1.32
+ $X2=0 $Y2=0
cc_221 N_A_225_413#_c_269_n N_A_339_93#_c_446_n 0.0363324f $X=1.9 $Y=1.915 $X2=0
+ $Y2=0
cc_222 N_A_225_413#_c_259_n N_A_339_93#_c_446_n 0.0285349f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_223 N_A_225_413#_c_262_n N_A_339_93#_c_446_n 0.0129756f $X=2.56 $Y=0.995
+ $X2=0 $Y2=0
cc_224 N_A_225_413#_c_264_n N_A_339_93#_c_459_n 0.00405026f $X=2.505 $Y=1.99
+ $X2=0 $Y2=0
cc_225 N_A_225_413#_c_264_n N_A_339_93#_c_450_n 0.0178382f $X=2.505 $Y=1.99
+ $X2=0 $Y2=0
cc_226 N_A_225_413#_c_259_n N_A_339_93#_c_450_n 0.00478459f $X=2.58 $Y=1.16
+ $X2=0 $Y2=0
cc_227 N_A_225_413#_c_260_n N_A_339_93#_c_450_n 0.00153955f $X=2.58 $Y=1.16
+ $X2=0 $Y2=0
cc_228 N_A_225_413#_c_265_n N_A_339_93#_c_453_n 0.0141285f $X=1.815 $Y=2 $X2=0
+ $Y2=0
cc_229 N_A_225_413#_c_265_n N_VPWR_M1012_s 0.0022786f $X=1.815 $Y=2 $X2=0 $Y2=0
cc_230 N_A_225_413#_c_264_n N_VPWR_c_533_n 4.94036e-19 $X=2.505 $Y=1.99 $X2=0
+ $Y2=0
cc_231 N_A_225_413#_c_283_n N_VPWR_c_533_n 0.0126073f $X=1.27 $Y=2.3 $X2=0 $Y2=0
cc_232 N_A_225_413#_c_265_n N_VPWR_c_533_n 0.021271f $X=1.815 $Y=2 $X2=0 $Y2=0
cc_233 N_A_225_413#_c_283_n N_VPWR_c_535_n 0.013862f $X=1.27 $Y=2.3 $X2=0 $Y2=0
cc_234 N_A_225_413#_c_265_n N_VPWR_c_535_n 0.00453603f $X=1.815 $Y=2 $X2=0 $Y2=0
cc_235 N_A_225_413#_c_264_n N_VPWR_c_537_n 0.00819146f $X=2.505 $Y=1.99 $X2=0
+ $Y2=0
cc_236 N_A_225_413#_c_264_n N_VPWR_c_538_n 0.00385862f $X=2.505 $Y=1.99 $X2=0
+ $Y2=0
cc_237 N_A_225_413#_c_265_n N_VPWR_c_538_n 5.29119e-19 $X=1.815 $Y=2 $X2=0 $Y2=0
cc_238 N_A_225_413#_M1004_d N_VPWR_c_532_n 0.00341979f $X=1.125 $Y=2.065 $X2=0
+ $Y2=0
cc_239 N_A_225_413#_c_264_n N_VPWR_c_532_n 0.00447322f $X=2.505 $Y=1.99 $X2=0
+ $Y2=0
cc_240 N_A_225_413#_c_283_n N_VPWR_c_532_n 0.0079665f $X=1.27 $Y=2.3 $X2=0 $Y2=0
cc_241 N_A_225_413#_c_265_n N_VPWR_c_532_n 0.00943611f $X=1.815 $Y=2 $X2=0 $Y2=0
cc_242 N_A_225_413#_c_256_n N_VGND_c_631_n 0.0698796f $X=2.495 $Y=0.34 $X2=0
+ $Y2=0
cc_243 N_A_225_413#_c_261_n N_VGND_c_631_n 0.0276904f $X=1.385 $Y=0.34 $X2=0
+ $Y2=0
cc_244 N_A_225_413#_c_262_n N_VGND_c_631_n 0.00357794f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_225_413#_M1007_d N_VGND_c_635_n 0.00382897f $X=1.135 $Y=0.235 $X2=0
+ $Y2=0
cc_246 N_A_225_413#_c_256_n N_VGND_c_635_n 0.0390712f $X=2.495 $Y=0.34 $X2=0
+ $Y2=0
cc_247 N_A_225_413#_c_261_n N_VGND_c_635_n 0.0152582f $X=1.385 $Y=0.34 $X2=0
+ $Y2=0
cc_248 N_A_225_413#_c_262_n N_VGND_c_635_n 0.0055808f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_A_225_413#_c_259_n A_511_93# 0.00394853f $X=2.58 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_250 N_C_c_359_n N_D_c_402_n 0.0119822f $X=3.025 $Y=1.89 $X2=0 $Y2=0
cc_251 C N_D_c_402_n 8.33079e-19 $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_252 N_C_c_360_n N_D_c_403_n 0.0201971f $X=3.025 $Y=1.99 $X2=0 $Y2=0
cc_253 N_C_c_359_n D 0.00100057f $X=3.025 $Y=1.89 $X2=0 $Y2=0
cc_254 C D 0.0969853f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_255 N_C_c_357_n D 0.00186563f $X=3.06 $Y=1.16 $X2=0 $Y2=0
cc_256 N_C_c_358_n D 0.00176743f $X=3.06 $Y=0.995 $X2=0 $Y2=0
cc_257 C N_D_c_400_n 3.54745e-19 $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_258 N_C_c_357_n N_D_c_400_n 0.0202531f $X=3.06 $Y=1.16 $X2=0 $Y2=0
cc_259 C N_D_c_401_n 0.00152811f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_260 N_C_c_358_n N_D_c_401_n 0.0229874f $X=3.06 $Y=0.995 $X2=0 $Y2=0
cc_261 C N_A_339_93#_c_446_n 0.0107074f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_262 N_C_c_360_n N_A_339_93#_c_450_n 0.0156108f $X=3.025 $Y=1.99 $X2=0 $Y2=0
cc_263 C N_A_339_93#_c_450_n 0.0160489f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_264 N_C_c_357_n N_A_339_93#_c_450_n 6.85542e-19 $X=3.06 $Y=1.16 $X2=0 $Y2=0
cc_265 N_C_c_360_n N_A_339_93#_c_481_n 0.00412322f $X=3.025 $Y=1.99 $X2=0 $Y2=0
cc_266 N_C_c_360_n N_VPWR_c_537_n 0.00331435f $X=3.025 $Y=1.99 $X2=0 $Y2=0
cc_267 N_C_c_360_n N_VPWR_c_540_n 0.00515029f $X=3.025 $Y=1.99 $X2=0 $Y2=0
cc_268 N_C_c_360_n N_VPWR_c_532_n 0.0068585f $X=3.025 $Y=1.99 $X2=0 $Y2=0
cc_269 C N_VGND_c_631_n 0.0101411f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_270 N_C_c_358_n N_VGND_c_631_n 0.00388886f $X=3.06 $Y=0.995 $X2=0 $Y2=0
cc_271 C N_VGND_c_635_n 0.00972827f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_272 N_C_c_358_n N_VGND_c_635_n 0.00609803f $X=3.06 $Y=0.995 $X2=0 $Y2=0
cc_273 C A_615_93# 0.00383554f $X=2.9 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_274 N_D_c_402_n N_A_339_93#_c_443_n 0.0190571f $X=3.575 $Y=1.89 $X2=0 $Y2=0
cc_275 N_D_c_403_n N_A_339_93#_c_443_n 0.0147349f $X=3.575 $Y=1.99 $X2=0 $Y2=0
cc_276 D N_A_339_93#_c_443_n 3.32786e-19 $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_277 N_D_c_400_n N_A_339_93#_c_443_n 0.0202459f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_278 D N_A_339_93#_c_444_n 0.00159999f $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_279 N_D_c_401_n N_A_339_93#_c_444_n 0.0207554f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_280 N_D_c_403_n N_A_339_93#_c_481_n 0.00417168f $X=3.575 $Y=1.99 $X2=0 $Y2=0
cc_281 N_D_c_403_n N_A_339_93#_c_451_n 0.0163111f $X=3.575 $Y=1.99 $X2=0 $Y2=0
cc_282 D N_A_339_93#_c_451_n 0.0140063f $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_283 N_D_c_400_n N_A_339_93#_c_451_n 2.50922e-19 $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_284 N_D_c_402_n N_A_339_93#_c_452_n 0.00837562f $X=3.575 $Y=1.89 $X2=0 $Y2=0
cc_285 D N_A_339_93#_c_452_n 0.0228651f $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_286 D N_A_339_93#_c_454_n 0.0022108f $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_287 D N_A_339_93#_c_447_n 0.0257124f $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_288 N_D_c_400_n N_A_339_93#_c_447_n 0.00191833f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_289 N_D_c_403_n N_VPWR_c_534_n 0.00434612f $X=3.575 $Y=1.99 $X2=0 $Y2=0
cc_290 N_D_c_403_n N_VPWR_c_540_n 0.00516667f $X=3.575 $Y=1.99 $X2=0 $Y2=0
cc_291 N_D_c_403_n N_VPWR_c_532_n 0.00699514f $X=3.575 $Y=1.99 $X2=0 $Y2=0
cc_292 D X 0.00459138f $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_293 D N_VGND_c_630_n 0.00914978f $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_294 N_D_c_401_n N_VGND_c_630_n 0.00735865f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_295 D N_VGND_c_631_n 0.00990013f $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_296 N_D_c_401_n N_VGND_c_631_n 0.00436733f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_297 D N_VGND_c_635_n 0.00969574f $X=3.39 $Y=0.425 $X2=0 $Y2=0
cc_298 N_D_c_401_n N_VGND_c_635_n 0.00741063f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_299 D A_615_93# 0.00371251f $X=3.39 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_300 N_A_339_93#_c_450_n N_VPWR_M1005_d 0.00231127f $X=3.21 $Y=2 $X2=0 $Y2=0
cc_301 N_A_339_93#_c_451_n N_VPWR_M1006_d 0.00552046f $X=3.81 $Y=2 $X2=0 $Y2=0
cc_302 N_A_339_93#_c_452_n N_VPWR_M1006_d 0.00709531f $X=3.895 $Y=1.915 $X2=0
+ $Y2=0
cc_303 N_A_339_93#_c_459_n N_VPWR_c_533_n 0.0122881f $X=2.27 $Y=2.3 $X2=0 $Y2=0
cc_304 N_A_339_93#_c_443_n N_VPWR_c_534_n 0.00896655f $X=4.1 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A_339_93#_c_451_n N_VPWR_c_534_n 0.0186919f $X=3.81 $Y=2 $X2=0 $Y2=0
cc_306 N_A_339_93#_c_459_n N_VPWR_c_537_n 0.0141017f $X=2.27 $Y=2.3 $X2=0 $Y2=0
cc_307 N_A_339_93#_c_450_n N_VPWR_c_537_n 0.0203444f $X=3.21 $Y=2 $X2=0 $Y2=0
cc_308 N_A_339_93#_c_459_n N_VPWR_c_538_n 0.0117826f $X=2.27 $Y=2.3 $X2=0 $Y2=0
cc_309 N_A_339_93#_c_450_n N_VPWR_c_538_n 0.00279618f $X=3.21 $Y=2 $X2=0 $Y2=0
cc_310 N_A_339_93#_c_453_n N_VPWR_c_538_n 4.17989e-19 $X=2.255 $Y=2 $X2=0 $Y2=0
cc_311 N_A_339_93#_c_450_n N_VPWR_c_540_n 0.00420952f $X=3.21 $Y=2 $X2=0 $Y2=0
cc_312 N_A_339_93#_c_481_n N_VPWR_c_540_n 0.0116326f $X=3.295 $Y=2.3 $X2=0 $Y2=0
cc_313 N_A_339_93#_c_451_n N_VPWR_c_540_n 0.00466831f $X=3.81 $Y=2 $X2=0 $Y2=0
cc_314 N_A_339_93#_c_443_n N_VPWR_c_541_n 0.00622633f $X=4.1 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A_339_93#_M1012_d N_VPWR_c_532_n 0.00384607f $X=2.115 $Y=2.065 $X2=0
+ $Y2=0
cc_316 N_A_339_93#_M1002_d N_VPWR_c_532_n 0.00366129f $X=3.115 $Y=2.065 $X2=0
+ $Y2=0
cc_317 N_A_339_93#_c_443_n N_VPWR_c_532_n 0.0113172f $X=4.1 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_339_93#_c_459_n N_VPWR_c_532_n 0.00646385f $X=2.27 $Y=2.3 $X2=0 $Y2=0
cc_319 N_A_339_93#_c_450_n N_VPWR_c_532_n 0.0134292f $X=3.21 $Y=2 $X2=0 $Y2=0
cc_320 N_A_339_93#_c_481_n N_VPWR_c_532_n 0.00643448f $X=3.295 $Y=2.3 $X2=0
+ $Y2=0
cc_321 N_A_339_93#_c_451_n N_VPWR_c_532_n 0.00944974f $X=3.81 $Y=2 $X2=0 $Y2=0
cc_322 N_A_339_93#_c_453_n N_VPWR_c_532_n 9.02646e-19 $X=2.255 $Y=2 $X2=0 $Y2=0
cc_323 N_A_339_93#_c_443_n X 0.0137578f $X=4.1 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A_339_93#_c_452_n X 0.0140305f $X=3.895 $Y=1.915 $X2=0 $Y2=0
cc_325 N_A_339_93#_c_443_n X 8.0628e-19 $X=4.1 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A_339_93#_c_444_n X 0.0148436f $X=4.125 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_339_93#_c_452_n X 0.00611378f $X=3.895 $Y=1.915 $X2=0 $Y2=0
cc_328 N_A_339_93#_c_447_n X 0.0251619f $X=4.02 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_339_93#_c_443_n N_VGND_c_630_n 0.00181646f $X=4.1 $Y=1.41 $X2=0 $Y2=0
cc_330 N_A_339_93#_c_444_n N_VGND_c_630_n 0.00425225f $X=4.125 $Y=0.995 $X2=0
+ $Y2=0
cc_331 N_A_339_93#_c_447_n N_VGND_c_630_n 0.00680524f $X=4.02 $Y=1.16 $X2=0
+ $Y2=0
cc_332 N_A_339_93#_c_444_n N_VGND_c_634_n 0.00585385f $X=4.125 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_A_339_93#_c_444_n N_VGND_c_635_n 0.0118099f $X=4.125 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_339_93#_c_445_n A_425_93# 0.00412933f $X=2.155 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_335 N_VPWR_c_532_n N_X_M1010_d 0.00425811f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_336 N_VPWR_c_534_n X 0.0131278f $X=3.865 $Y=2.34 $X2=0 $Y2=0
cc_337 N_VPWR_c_541_n X 0.0182101f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_338 N_VPWR_c_532_n X 0.00993603f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_339 N_X_c_612_n N_VGND_c_634_n 0.0179758f $X=4.335 $Y=0.42 $X2=0 $Y2=0
cc_340 N_X_M1013_d N_VGND_c_635_n 0.00382897f $X=4.2 $Y=0.235 $X2=0 $Y2=0
cc_341 N_X_c_612_n N_VGND_c_635_n 0.00993004f $X=4.335 $Y=0.42 $X2=0 $Y2=0
