* File: sky130_fd_sc_hdll__bufinv_16.pex.spice
* Created: Wed Sep  2 08:24:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUFINV_16%A 3 5 7 10 12 14 15 17 20 22 30 31
c69 30 0 1.39726e-19 $X=1.07 $Y=1.16
c70 20 0 1.25206e-19 $X=1.46 $Y=0.56
c71 15 0 1.26528e-19 $X=1.435 $Y=1.41
r72 31 32 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.217
+ $X2=1.46 $Y2=1.217
r73 29 31 53.3121 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=1.07 $Y=1.217
+ $X2=1.435 $Y2=1.217
r74 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.07
+ $Y=1.16 $X2=1.07 $Y2=1.16
r75 27 29 15.3364 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.965 $Y=1.217
+ $X2=1.07 $Y2=1.217
r76 26 27 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.217
+ $X2=0.965 $Y2=1.217
r77 25 26 64.997 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.217
+ $X2=0.94 $Y2=1.217
r78 24 25 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.217
+ $X2=0.495 $Y2=1.217
r79 22 30 46.3045 $w=1.98e-07 $l=8.35e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=1.07 $Y2=1.175
r80 18 32 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.217
r81 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r82 15 31 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.217
r83 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r84 12 27 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.217
r85 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r86 8 26 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=1.217
r87 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=0.56
r88 5 25 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.217
r89 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r90 1 24 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.217
r91 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_16%A_27_47# 1 2 3 4 15 17 19 22 24 26 29 31
+ 33 36 38 40 43 45 47 48 50 53 57 61 65 66 67 68 71 75 79 81 84 86 92 95 96 97
+ 110
c208 110 0 1.39726e-19 $X=4.255 $Y=1.217
c209 92 0 1.34672e-19 $X=3.91 $Y=1.16
c210 53 0 1.25206e-19 $X=4.28 $Y=0.56
c211 48 0 1.26528e-19 $X=4.255 $Y=1.41
r212 110 111 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=4.255 $Y=1.217
+ $X2=4.28 $Y2=1.217
r213 107 108 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.217
+ $X2=3.785 $Y2=1.217
r214 106 107 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=3.315 $Y=1.217
+ $X2=3.76 $Y2=1.217
r215 105 106 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.217
+ $X2=3.315 $Y2=1.217
r216 104 105 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=3.29 $Y2=1.217
r217 103 104 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.217
+ $X2=2.845 $Y2=1.217
r218 102 103 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.82 $Y2=1.217
r219 101 102 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r220 98 99 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.217
+ $X2=1.905 $Y2=1.217
r221 93 110 51.3241 $w=3.24e-07 $l=3.45e-07 $layer=POLY_cond $X=3.91 $Y=1.217
+ $X2=4.255 $Y2=1.217
r222 93 108 18.5957 $w=3.24e-07 $l=1.25e-07 $layer=POLY_cond $X=3.91 $Y=1.217
+ $X2=3.785 $Y2=1.217
r223 92 93 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.91
+ $Y=1.16 $X2=3.91 $Y2=1.16
r224 90 101 50.5802 $w=3.24e-07 $l=3.4e-07 $layer=POLY_cond $X=2.01 $Y=1.217
+ $X2=2.35 $Y2=1.217
r225 90 99 15.6204 $w=3.24e-07 $l=1.05e-07 $layer=POLY_cond $X=2.01 $Y=1.217
+ $X2=1.905 $Y2=1.217
r226 89 92 105.364 $w=1.98e-07 $l=1.9e-06 $layer=LI1_cond $X=2.01 $Y=1.175
+ $X2=3.91 $Y2=1.175
r227 89 90 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.01
+ $Y=1.16 $X2=2.01 $Y2=1.16
r228 87 97 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=1.175
+ $X2=1.67 $Y2=1.175
r229 87 89 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=1.755 $Y=1.175
+ $X2=2.01 $Y2=1.175
r230 85 97 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.67 $Y=1.275 $X2=1.67
+ $Y2=1.175
r231 85 86 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.67 $Y=1.275
+ $X2=1.67 $Y2=1.445
r232 84 97 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.67 $Y=1.075 $X2=1.67
+ $Y2=1.175
r233 83 84 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.67 $Y=0.905
+ $X2=1.67 $Y2=1.075
r234 82 96 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=1.53
+ $X2=1.175 $Y2=1.53
r235 81 86 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.585 $Y=1.53
+ $X2=1.67 $Y2=1.445
r236 81 82 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.585 $Y=1.53
+ $X2=1.365 $Y2=1.53
r237 80 95 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0.82
+ $X2=1.175 $Y2=0.82
r238 79 83 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.585 $Y=0.82
+ $X2=1.67 $Y2=0.905
r239 79 80 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.585 $Y=0.82
+ $X2=1.365 $Y2=0.82
r240 75 77 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.175 $Y=1.63
+ $X2=1.175 $Y2=2.31
r241 73 96 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=1.615
+ $X2=1.175 $Y2=1.53
r242 73 75 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.175 $Y=1.615
+ $X2=1.175 $Y2=1.63
r243 69 95 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=0.735
+ $X2=1.175 $Y2=0.82
r244 69 71 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.175 $Y=0.735
+ $X2=1.175 $Y2=0.4
r245 67 96 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=1.53
+ $X2=1.175 $Y2=1.53
r246 67 68 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=1.53
+ $X2=0.425 $Y2=1.53
r247 65 95 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0.82
+ $X2=1.175 $Y2=0.82
r248 65 66 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.82
+ $X2=0.425 $Y2=0.82
r249 61 63 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r250 59 68 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.425 $Y2=1.53
r251 59 61 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.63
r252 55 66 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.425 $Y2=0.82
r253 55 57 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.4
r254 51 111 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.28 $Y=1.025
+ $X2=4.28 $Y2=1.217
r255 51 53 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.28 $Y=1.025
+ $X2=4.28 $Y2=0.56
r256 48 110 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.217
r257 48 50 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r258 45 108 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.217
r259 45 47 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r260 41 107 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.76 $Y=1.025
+ $X2=3.76 $Y2=1.217
r261 41 43 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.76 $Y=1.025
+ $X2=3.76 $Y2=0.56
r262 38 106 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r263 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r264 34 105 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r265 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r266 31 104 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r267 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r268 27 103 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=1.217
r269 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=0.56
r270 24 102 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r271 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r272 20 101 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r273 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
r274 17 99 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r275 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r276 13 98 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=1.217
r277 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=0.56
r278 4 77 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.31
r279 4 75 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.63
r280 3 63 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r281 3 61 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r282 2 71 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.4
r283 1 57 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_16%A_391_47# 1 2 3 4 5 6 21 23 25 28 30 32
+ 35 37 39 42 44 46 49 51 53 56 58 60 63 65 67 70 72 74 77 79 81 84 86 88 91 93
+ 95 98 100 102 105 107 109 112 114 116 119 121 123 124 126 129 133 137 141 142
+ 143 144 147 151 155 157 161 165 169 171 174 176 182 185 186 187 188 189 222
c462 222 0 1.34672e-19 $X=11.775 $Y=1.217
c463 144 0 1.26528e-19 $X=2.305 $Y=1.53
c464 142 0 1.25206e-19 $X=2.305 $Y=0.82
r465 222 223 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=11.775 $Y=1.217
+ $X2=11.8 $Y2=1.217
r466 221 222 70.7937 $w=3.2e-07 $l=4.7e-07 $layer=POLY_cond $X=11.305 $Y=1.217
+ $X2=11.775 $Y2=1.217
r467 218 219 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=10.835 $Y=1.217
+ $X2=11.28 $Y2=1.217
r468 217 218 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=10.81 $Y=1.217
+ $X2=10.835 $Y2=1.217
r469 216 217 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=10.365 $Y=1.217
+ $X2=10.81 $Y2=1.217
r470 215 216 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=10.34 $Y=1.217
+ $X2=10.365 $Y2=1.217
r471 214 215 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=9.895 $Y=1.217
+ $X2=10.34 $Y2=1.217
r472 213 214 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=9.87 $Y=1.217
+ $X2=9.895 $Y2=1.217
r473 212 213 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=9.425 $Y=1.217
+ $X2=9.87 $Y2=1.217
r474 211 212 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=9.4 $Y=1.217
+ $X2=9.425 $Y2=1.217
r475 210 211 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=8.955 $Y=1.217
+ $X2=9.4 $Y2=1.217
r476 209 210 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=8.93 $Y=1.217
+ $X2=8.955 $Y2=1.217
r477 208 209 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=8.485 $Y=1.217
+ $X2=8.93 $Y2=1.217
r478 207 208 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=8.46 $Y=1.217
+ $X2=8.485 $Y2=1.217
r479 206 207 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=8.015 $Y=1.217
+ $X2=8.46 $Y2=1.217
r480 205 206 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=7.99 $Y=1.217
+ $X2=8.015 $Y2=1.217
r481 204 205 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=7.545 $Y=1.217
+ $X2=7.99 $Y2=1.217
r482 203 204 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=7.52 $Y=1.217
+ $X2=7.545 $Y2=1.217
r483 202 203 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=7.075 $Y=1.217
+ $X2=7.52 $Y2=1.217
r484 201 202 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=7.05 $Y=1.217
+ $X2=7.075 $Y2=1.217
r485 200 201 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=6.605 $Y=1.217
+ $X2=7.05 $Y2=1.217
r486 199 200 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=6.58 $Y=1.217
+ $X2=6.605 $Y2=1.217
r487 198 199 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=6.135 $Y=1.217
+ $X2=6.58 $Y2=1.217
r488 197 198 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=6.11 $Y=1.217
+ $X2=6.135 $Y2=1.217
r489 196 197 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=5.665 $Y=1.217
+ $X2=6.11 $Y2=1.217
r490 195 196 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=5.64 $Y=1.217
+ $X2=5.665 $Y2=1.217
r491 194 195 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=5.195 $Y=1.217
+ $X2=5.64 $Y2=1.217
r492 193 194 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.217
+ $X2=5.195 $Y2=1.217
r493 190 191 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.217
+ $X2=4.725 $Y2=1.217
r494 183 221 2.25938 $w=3.2e-07 $l=1.5e-08 $layer=POLY_cond $X=11.29 $Y=1.217
+ $X2=11.305 $Y2=1.217
r495 183 219 1.50625 $w=3.2e-07 $l=1e-08 $layer=POLY_cond $X=11.29 $Y=1.217
+ $X2=11.28 $Y2=1.217
r496 182 183 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=11.29
+ $Y=1.16 $X2=11.29 $Y2=1.16
r497 180 193 54.225 $w=3.2e-07 $l=3.6e-07 $layer=POLY_cond $X=4.81 $Y=1.217
+ $X2=5.17 $Y2=1.217
r498 180 191 12.8031 $w=3.2e-07 $l=8.5e-08 $layer=POLY_cond $X=4.81 $Y=1.217
+ $X2=4.725 $Y2=1.217
r499 179 182 359.345 $w=1.98e-07 $l=6.48e-06 $layer=LI1_cond $X=4.81 $Y=1.175
+ $X2=11.29 $Y2=1.175
r500 179 180 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=4.81
+ $Y=1.16 $X2=4.81 $Y2=1.16
r501 177 189 0.866423 $w=2e-07 $l=8.8e-08 $layer=LI1_cond $X=4.575 $Y=1.175
+ $X2=4.487 $Y2=1.175
r502 177 179 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=4.575 $Y=1.175
+ $X2=4.81 $Y2=1.175
r503 175 189 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=4.487 $Y=1.275
+ $X2=4.487 $Y2=1.175
r504 175 176 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=4.487 $Y=1.275
+ $X2=4.487 $Y2=1.445
r505 174 189 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=4.487 $Y=1.075
+ $X2=4.487 $Y2=1.175
r506 173 174 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=4.487 $Y=0.905
+ $X2=4.487 $Y2=1.075
r507 172 188 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.185 $Y=1.53
+ $X2=3.995 $Y2=1.53
r508 171 176 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=4.4 $Y=1.53
+ $X2=4.487 $Y2=1.445
r509 171 172 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.4 $Y=1.53
+ $X2=4.185 $Y2=1.53
r510 170 187 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.185 $Y=0.82
+ $X2=3.995 $Y2=0.82
r511 169 173 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=4.4 $Y=0.82
+ $X2=4.487 $Y2=0.905
r512 169 170 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.4 $Y=0.82
+ $X2=4.185 $Y2=0.82
r513 165 167 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.995 $Y=1.63
+ $X2=3.995 $Y2=2.31
r514 163 188 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=1.615
+ $X2=3.995 $Y2=1.53
r515 163 165 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.995 $Y=1.615
+ $X2=3.995 $Y2=1.63
r516 159 187 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=0.735
+ $X2=3.995 $Y2=0.82
r517 159 161 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.995 $Y=0.735
+ $X2=3.995 $Y2=0.4
r518 158 186 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.245 $Y=1.53
+ $X2=3.055 $Y2=1.53
r519 157 188 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=1.53
+ $X2=3.995 $Y2=1.53
r520 157 158 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.805 $Y=1.53
+ $X2=3.245 $Y2=1.53
r521 156 185 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.245 $Y=0.82
+ $X2=3.055 $Y2=0.82
r522 155 187 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=0.82
+ $X2=3.995 $Y2=0.82
r523 155 156 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.805 $Y=0.82
+ $X2=3.245 $Y2=0.82
r524 151 153 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.055 $Y=1.63
+ $X2=3.055 $Y2=2.31
r525 149 186 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=1.615
+ $X2=3.055 $Y2=1.53
r526 149 151 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.055 $Y=1.615
+ $X2=3.055 $Y2=1.63
r527 145 185 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.735
+ $X2=3.055 $Y2=0.82
r528 145 147 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.055 $Y=0.735
+ $X2=3.055 $Y2=0.4
r529 143 186 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=1.53
+ $X2=3.055 $Y2=1.53
r530 143 144 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.865 $Y=1.53
+ $X2=2.305 $Y2=1.53
r531 141 185 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=0.82
+ $X2=3.055 $Y2=0.82
r532 141 142 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.865 $Y=0.82
+ $X2=2.305 $Y2=0.82
r533 137 139 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.115 $Y=1.63
+ $X2=2.115 $Y2=2.31
r534 135 144 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.115 $Y=1.615
+ $X2=2.305 $Y2=1.53
r535 135 137 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.115 $Y=1.615
+ $X2=2.115 $Y2=1.63
r536 131 142 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.115 $Y=0.735
+ $X2=2.305 $Y2=0.82
r537 131 133 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.115 $Y=0.735
+ $X2=2.115 $Y2=0.4
r538 127 223 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=11.8 $Y=1.025
+ $X2=11.8 $Y2=1.217
r539 127 129 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.8 $Y=1.025
+ $X2=11.8 $Y2=0.56
r540 124 222 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=11.775 $Y=1.41
+ $X2=11.775 $Y2=1.217
r541 124 126 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.775 $Y=1.41
+ $X2=11.775 $Y2=1.985
r542 121 221 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=11.305 $Y=1.41
+ $X2=11.305 $Y2=1.217
r543 121 123 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.305 $Y=1.41
+ $X2=11.305 $Y2=1.985
r544 117 219 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=11.28 $Y=1.025
+ $X2=11.28 $Y2=1.217
r545 117 119 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.28 $Y=1.025
+ $X2=11.28 $Y2=0.56
r546 114 218 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.835 $Y=1.41
+ $X2=10.835 $Y2=1.217
r547 114 116 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.835 $Y=1.41
+ $X2=10.835 $Y2=1.985
r548 110 217 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10.81 $Y=1.025
+ $X2=10.81 $Y2=1.217
r549 110 112 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.81 $Y=1.025
+ $X2=10.81 $Y2=0.56
r550 107 216 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.365 $Y=1.41
+ $X2=10.365 $Y2=1.217
r551 107 109 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.365 $Y=1.41
+ $X2=10.365 $Y2=1.985
r552 103 215 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10.34 $Y=1.025
+ $X2=10.34 $Y2=1.217
r553 103 105 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.34 $Y=1.025
+ $X2=10.34 $Y2=0.56
r554 100 214 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.895 $Y=1.41
+ $X2=9.895 $Y2=1.217
r555 100 102 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.895 $Y=1.41
+ $X2=9.895 $Y2=1.985
r556 96 213 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.87 $Y=1.025
+ $X2=9.87 $Y2=1.217
r557 96 98 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.87 $Y=1.025
+ $X2=9.87 $Y2=0.56
r558 93 212 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.425 $Y=1.41
+ $X2=9.425 $Y2=1.217
r559 93 95 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.425 $Y=1.41
+ $X2=9.425 $Y2=1.985
r560 89 211 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.4 $Y=1.025
+ $X2=9.4 $Y2=1.217
r561 89 91 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.4 $Y=1.025
+ $X2=9.4 $Y2=0.56
r562 86 210 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.955 $Y=1.41
+ $X2=8.955 $Y2=1.217
r563 86 88 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.955 $Y=1.41
+ $X2=8.955 $Y2=1.985
r564 82 209 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.93 $Y=1.025
+ $X2=8.93 $Y2=1.217
r565 82 84 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.93 $Y=1.025
+ $X2=8.93 $Y2=0.56
r566 79 208 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.217
r567 79 81 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.985
r568 75 207 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.46 $Y=1.025
+ $X2=8.46 $Y2=1.217
r569 75 77 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.46 $Y=1.025
+ $X2=8.46 $Y2=0.56
r570 72 206 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.217
r571 72 74 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.985
r572 68 205 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.99 $Y=1.025
+ $X2=7.99 $Y2=1.217
r573 68 70 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.99 $Y=1.025
+ $X2=7.99 $Y2=0.56
r574 65 204 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.217
r575 65 67 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.985
r576 61 203 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.52 $Y=1.025
+ $X2=7.52 $Y2=1.217
r577 61 63 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.52 $Y=1.025
+ $X2=7.52 $Y2=0.56
r578 58 202 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.217
r579 58 60 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.985
r580 54 201 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.05 $Y=1.025
+ $X2=7.05 $Y2=1.217
r581 54 56 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.05 $Y=1.025
+ $X2=7.05 $Y2=0.56
r582 51 200 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.217
r583 51 53 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.985
r584 47 199 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.58 $Y=1.025
+ $X2=6.58 $Y2=1.217
r585 47 49 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.58 $Y=1.025
+ $X2=6.58 $Y2=0.56
r586 44 198 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.217
r587 44 46 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.985
r588 40 197 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.11 $Y=1.025
+ $X2=6.11 $Y2=1.217
r589 40 42 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.11 $Y=1.025
+ $X2=6.11 $Y2=0.56
r590 37 196 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.217
r591 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r592 33 195 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.64 $Y=1.025
+ $X2=5.64 $Y2=1.217
r593 33 35 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.64 $Y=1.025
+ $X2=5.64 $Y2=0.56
r594 30 194 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.217
r595 30 32 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r596 26 193 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=1.217
r597 26 28 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=0.56
r598 23 191 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.217
r599 23 25 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r600 19 190 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=1.217
r601 19 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=0.56
r602 6 167 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2.31
r603 6 165 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.63
r604 5 153 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2.31
r605 5 151 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.63
r606 4 139 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.31
r607 4 137 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.63
r608 3 161 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.4
r609 2 147 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.4
r610 1 133 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 44 46
+ 50 52 56 60 64 68 72 76 80 84 88 92 96 99 100 102 103 105 106 108 109 111 112
+ 114 115 117 118 120 121 123 124 126 127 128 162 163 166 169 172 175
r207 172 173 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r208 170 173 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r209 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r210 167 170 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r211 166 167 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r212 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r213 160 163 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r214 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r215 157 160 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.73 $Y2=2.72
r216 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r217 154 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r218 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r219 151 154 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r220 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r221 148 151 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r222 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r223 145 148 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r224 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r225 142 145 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r226 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r227 139 142 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r228 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r229 136 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r230 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r231 133 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r232 133 173 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r233 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r234 130 172 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.61 $Y2=2.72
r235 130 132 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=3.45 $Y2=2.72
r236 128 167 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r237 128 175 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r238 126 159 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=11.925 $Y=2.72
+ $X2=11.73 $Y2=2.72
r239 126 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.925 $Y=2.72
+ $X2=12.01 $Y2=2.72
r240 125 162 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=12.095 $Y=2.72
+ $X2=12.19 $Y2=2.72
r241 125 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.095 $Y=2.72
+ $X2=12.01 $Y2=2.72
r242 123 156 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.985 $Y=2.72
+ $X2=10.81 $Y2=2.72
r243 123 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.985 $Y=2.72
+ $X2=11.07 $Y2=2.72
r244 122 159 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=11.155 $Y=2.72
+ $X2=11.73 $Y2=2.72
r245 122 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.155 $Y=2.72
+ $X2=11.07 $Y2=2.72
r246 120 153 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.045 $Y=2.72
+ $X2=9.89 $Y2=2.72
r247 120 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.045 $Y=2.72
+ $X2=10.13 $Y2=2.72
r248 119 156 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=10.215 $Y=2.72
+ $X2=10.81 $Y2=2.72
r249 119 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.215 $Y=2.72
+ $X2=10.13 $Y2=2.72
r250 117 150 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=9.105 $Y=2.72
+ $X2=8.97 $Y2=2.72
r251 117 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.105 $Y=2.72
+ $X2=9.19 $Y2=2.72
r252 116 153 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=9.275 $Y=2.72
+ $X2=9.89 $Y2=2.72
r253 116 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.275 $Y=2.72
+ $X2=9.19 $Y2=2.72
r254 114 147 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.165 $Y=2.72
+ $X2=8.05 $Y2=2.72
r255 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.165 $Y=2.72
+ $X2=8.25 $Y2=2.72
r256 113 150 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.335 $Y=2.72
+ $X2=8.97 $Y2=2.72
r257 113 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=2.72
+ $X2=8.25 $Y2=2.72
r258 111 144 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.225 $Y=2.72
+ $X2=7.13 $Y2=2.72
r259 111 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.225 $Y=2.72
+ $X2=7.31 $Y2=2.72
r260 110 147 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=7.395 $Y=2.72
+ $X2=8.05 $Y2=2.72
r261 110 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=2.72
+ $X2=7.31 $Y2=2.72
r262 108 141 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.285 $Y=2.72
+ $X2=6.21 $Y2=2.72
r263 108 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.285 $Y=2.72
+ $X2=6.37 $Y2=2.72
r264 107 144 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.455 $Y=2.72
+ $X2=7.13 $Y2=2.72
r265 107 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=2.72
+ $X2=6.37 $Y2=2.72
r266 105 138 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.29 $Y2=2.72
r267 105 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.43 $Y2=2.72
r268 104 141 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.515 $Y=2.72
+ $X2=6.21 $Y2=2.72
r269 104 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.515 $Y=2.72
+ $X2=5.43 $Y2=2.72
r270 102 135 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.405 $Y=2.72
+ $X2=4.37 $Y2=2.72
r271 102 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=2.72
+ $X2=4.49 $Y2=2.72
r272 101 138 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=4.575 $Y=2.72
+ $X2=5.29 $Y2=2.72
r273 101 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=2.72
+ $X2=4.49 $Y2=2.72
r274 99 132 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.45 $Y2=2.72
r275 99 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.55 $Y2=2.72
r276 98 135 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=4.37 $Y2=2.72
r277 98 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=3.55 $Y2=2.72
r278 94 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.01 $Y=2.635
+ $X2=12.01 $Y2=2.72
r279 94 96 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=12.01 $Y=2.635
+ $X2=12.01 $Y2=2
r280 90 124 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.07 $Y=2.635
+ $X2=11.07 $Y2=2.72
r281 90 92 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.07 $Y=2.635
+ $X2=11.07 $Y2=2
r282 86 121 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.13 $Y=2.635
+ $X2=10.13 $Y2=2.72
r283 86 88 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.13 $Y=2.635
+ $X2=10.13 $Y2=2
r284 82 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.19 $Y=2.635
+ $X2=9.19 $Y2=2.72
r285 82 84 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.19 $Y=2.635
+ $X2=9.19 $Y2=2
r286 78 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.25 $Y=2.635
+ $X2=8.25 $Y2=2.72
r287 78 80 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.25 $Y=2.635
+ $X2=8.25 $Y2=2
r288 74 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=2.635
+ $X2=7.31 $Y2=2.72
r289 74 76 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.31 $Y=2.635
+ $X2=7.31 $Y2=2
r290 70 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=2.635
+ $X2=6.37 $Y2=2.72
r291 70 72 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.37 $Y=2.635
+ $X2=6.37 $Y2=2
r292 66 106 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=2.635
+ $X2=5.43 $Y2=2.72
r293 66 68 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.43 $Y=2.635
+ $X2=5.43 $Y2=2
r294 62 103 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=2.635
+ $X2=4.49 $Y2=2.72
r295 62 64 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.49 $Y=2.635
+ $X2=4.49 $Y2=2
r296 58 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2.72
r297 58 60 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2
r298 54 172 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=2.72
r299 54 56 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=2
r300 53 169 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=2.72
+ $X2=1.67 $Y2=2.72
r301 52 172 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.61 $Y2=2.72
r302 52 53 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=1.755 $Y2=2.72
r303 48 169 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r304 48 50 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2
r305 47 166 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.73 $Y2=2.72
r306 46 169 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=1.67 $Y2=2.72
r307 46 47 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=0.815 $Y2=2.72
r308 42 166 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r309 42 44 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2
r310 13 96 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=11.865
+ $Y=1.485 $X2=12.01 $Y2=2
r311 12 92 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=10.925
+ $Y=1.485 $X2=11.07 $Y2=2
r312 11 88 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.985
+ $Y=1.485 $X2=10.13 $Y2=2
r313 10 84 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.045
+ $Y=1.485 $X2=9.19 $Y2=2
r314 9 80 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.105
+ $Y=1.485 $X2=8.25 $Y2=2
r315 8 76 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=2
r316 7 72 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=2
r317 6 68 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2
r318 5 64 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2
r319 4 60 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2
r320 3 56 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2
r321 2 50 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2
r322 1 44 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 49 50 53 57 58 59 60 61 62 65 69 71 73 74 77 81 83 87 91 95 97 101 105 109 111
+ 115 119 123 125 129 133 137 139 143 147 151 153 159 160 163 164 165 166 167
+ 168 169 170 171 172 173 174 176 177
c363 60 0 1.26528e-19 $X=5.125 $Y=1.53
c364 58 0 1.25206e-19 $X=5.125 $Y=0.82
r365 176 177 8.27522 $w=4.43e-07 $l=2.55e-07 $layer=LI1_cond $X=12.067 $Y=1.19
+ $X2=12.067 $Y2=1.445
r366 175 176 11.9435 $w=2.73e-07 $l=2.85e-07 $layer=LI1_cond $X=12.067 $Y=0.905
+ $X2=12.067 $Y2=1.19
r367 154 174 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.705 $Y=1.53
+ $X2=11.515 $Y2=1.53
r368 153 177 4.51856 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=11.93 $Y=1.53
+ $X2=12.067 $Y2=1.53
r369 153 154 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.93 $Y=1.53
+ $X2=11.705 $Y2=1.53
r370 152 173 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.705 $Y=0.82
+ $X2=11.515 $Y2=0.82
r371 151 175 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=11.93 $Y=0.82
+ $X2=12.067 $Y2=0.905
r372 151 152 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.93 $Y=0.82
+ $X2=11.705 $Y2=0.82
r373 147 149 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=11.515 $Y=1.63
+ $X2=11.515 $Y2=2.31
r374 145 174 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.515 $Y=1.615
+ $X2=11.515 $Y2=1.53
r375 145 147 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=11.515 $Y=1.615
+ $X2=11.515 $Y2=1.63
r376 141 173 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.515 $Y=0.735
+ $X2=11.515 $Y2=0.82
r377 141 143 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=11.515 $Y=0.735
+ $X2=11.515 $Y2=0.4
r378 140 172 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.765 $Y=1.53
+ $X2=10.575 $Y2=1.53
r379 139 174 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.325 $Y=1.53
+ $X2=11.515 $Y2=1.53
r380 139 140 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=11.325 $Y=1.53
+ $X2=10.765 $Y2=1.53
r381 138 171 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.765 $Y=0.82
+ $X2=10.575 $Y2=0.82
r382 137 173 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.325 $Y=0.82
+ $X2=11.515 $Y2=0.82
r383 137 138 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=11.325 $Y=0.82
+ $X2=10.765 $Y2=0.82
r384 133 135 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=10.575 $Y=1.63
+ $X2=10.575 $Y2=2.31
r385 131 172 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.575 $Y=1.615
+ $X2=10.575 $Y2=1.53
r386 131 133 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=10.575 $Y=1.615
+ $X2=10.575 $Y2=1.63
r387 127 171 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.575 $Y=0.735
+ $X2=10.575 $Y2=0.82
r388 127 129 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=10.575 $Y=0.735
+ $X2=10.575 $Y2=0.4
r389 126 170 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.825 $Y=1.53
+ $X2=9.635 $Y2=1.53
r390 125 172 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.385 $Y=1.53
+ $X2=10.575 $Y2=1.53
r391 125 126 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=10.385 $Y=1.53
+ $X2=9.825 $Y2=1.53
r392 124 169 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.825 $Y=0.82
+ $X2=9.635 $Y2=0.82
r393 123 171 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.385 $Y=0.82
+ $X2=10.575 $Y2=0.82
r394 123 124 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=10.385 $Y=0.82
+ $X2=9.825 $Y2=0.82
r395 119 121 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=9.635 $Y=1.63
+ $X2=9.635 $Y2=2.31
r396 117 170 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.635 $Y=1.615
+ $X2=9.635 $Y2=1.53
r397 117 119 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=9.635 $Y=1.615
+ $X2=9.635 $Y2=1.63
r398 113 169 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.635 $Y=0.735
+ $X2=9.635 $Y2=0.82
r399 113 115 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.635 $Y=0.735
+ $X2=9.635 $Y2=0.4
r400 112 168 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.885 $Y=1.53
+ $X2=8.695 $Y2=1.53
r401 111 170 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.445 $Y=1.53
+ $X2=9.635 $Y2=1.53
r402 111 112 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=9.445 $Y=1.53
+ $X2=8.885 $Y2=1.53
r403 110 167 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.885 $Y=0.82
+ $X2=8.695 $Y2=0.82
r404 109 169 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.445 $Y=0.82
+ $X2=9.635 $Y2=0.82
r405 109 110 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=9.445 $Y=0.82
+ $X2=8.885 $Y2=0.82
r406 105 107 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=8.695 $Y=1.63
+ $X2=8.695 $Y2=2.31
r407 103 168 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.695 $Y=1.615
+ $X2=8.695 $Y2=1.53
r408 103 105 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=8.695 $Y=1.615
+ $X2=8.695 $Y2=1.63
r409 99 167 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.695 $Y=0.735
+ $X2=8.695 $Y2=0.82
r410 99 101 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.695 $Y=0.735
+ $X2=8.695 $Y2=0.4
r411 98 166 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.945 $Y=1.53
+ $X2=7.755 $Y2=1.53
r412 97 168 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.505 $Y=1.53
+ $X2=8.695 $Y2=1.53
r413 97 98 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.505 $Y=1.53
+ $X2=7.945 $Y2=1.53
r414 96 165 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.945 $Y=0.82
+ $X2=7.755 $Y2=0.82
r415 95 167 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.505 $Y=0.82
+ $X2=8.695 $Y2=0.82
r416 95 96 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.505 $Y=0.82
+ $X2=7.945 $Y2=0.82
r417 91 93 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=7.755 $Y=1.63
+ $X2=7.755 $Y2=2.31
r418 89 166 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.755 $Y=1.615
+ $X2=7.755 $Y2=1.53
r419 89 91 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=7.755 $Y=1.615
+ $X2=7.755 $Y2=1.63
r420 85 165 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.755 $Y=0.735
+ $X2=7.755 $Y2=0.82
r421 85 87 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.755 $Y=0.735
+ $X2=7.755 $Y2=0.4
r422 84 164 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.005 $Y=1.53
+ $X2=6.815 $Y2=1.53
r423 83 166 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.565 $Y=1.53
+ $X2=7.755 $Y2=1.53
r424 83 84 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.565 $Y=1.53
+ $X2=7.005 $Y2=1.53
r425 82 163 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.005 $Y=0.82
+ $X2=6.815 $Y2=0.82
r426 81 165 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.565 $Y=0.82
+ $X2=7.755 $Y2=0.82
r427 81 82 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.565 $Y=0.82
+ $X2=7.005 $Y2=0.82
r428 77 79 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.815 $Y=1.63
+ $X2=6.815 $Y2=2.31
r429 75 164 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=1.615
+ $X2=6.815 $Y2=1.53
r430 75 77 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=6.815 $Y=1.615
+ $X2=6.815 $Y2=1.63
r431 74 163 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=0.735
+ $X2=6.815 $Y2=0.82
r432 73 162 1.60526 $w=3.8e-07 $l=5e-08 $layer=LI1_cond $X=6.815 $Y=0.45
+ $X2=6.815 $Y2=0.4
r433 73 74 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=6.815 $Y=0.45
+ $X2=6.815 $Y2=0.735
r434 72 160 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.065 $Y=1.53
+ $X2=5.875 $Y2=1.53
r435 71 164 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.625 $Y=1.53
+ $X2=6.815 $Y2=1.53
r436 71 72 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.625 $Y=1.53
+ $X2=6.065 $Y2=1.53
r437 70 159 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.065 $Y=0.82
+ $X2=5.875 $Y2=0.82
r438 69 163 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.625 $Y=0.82
+ $X2=6.815 $Y2=0.82
r439 69 70 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.625 $Y=0.82
+ $X2=6.065 $Y2=0.82
r440 65 67 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=5.875 $Y=1.63
+ $X2=5.875 $Y2=2.31
r441 63 160 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=1.615
+ $X2=5.875 $Y2=1.53
r442 63 65 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=5.875 $Y=1.615
+ $X2=5.875 $Y2=1.63
r443 62 159 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=0.735
+ $X2=5.875 $Y2=0.82
r444 61 158 1.60526 $w=3.8e-07 $l=5e-08 $layer=LI1_cond $X=5.875 $Y=0.45
+ $X2=5.875 $Y2=0.4
r445 61 62 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=5.875 $Y=0.45
+ $X2=5.875 $Y2=0.735
r446 59 160 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.685 $Y=1.53
+ $X2=5.875 $Y2=1.53
r447 59 60 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.685 $Y=1.53
+ $X2=5.125 $Y2=1.53
r448 57 159 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.685 $Y=0.82
+ $X2=5.875 $Y2=0.82
r449 57 58 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.685 $Y=0.82
+ $X2=5.125 $Y2=0.82
r450 53 55 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=4.935 $Y=1.63
+ $X2=4.935 $Y2=2.31
r451 51 60 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=4.935 $Y=1.615
+ $X2=5.125 $Y2=1.53
r452 51 53 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=4.935 $Y=1.615
+ $X2=4.935 $Y2=1.63
r453 50 58 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=4.935 $Y=0.735
+ $X2=5.125 $Y2=0.82
r454 49 156 1.60526 $w=3.8e-07 $l=5e-08 $layer=LI1_cond $X=4.935 $Y=0.45
+ $X2=4.935 $Y2=0.4
r455 49 50 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=4.935 $Y=0.45
+ $X2=4.935 $Y2=0.735
r456 16 149 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=11.395
+ $Y=1.485 $X2=11.54 $Y2=2.31
r457 16 147 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.395
+ $Y=1.485 $X2=11.54 $Y2=1.63
r458 15 135 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.455
+ $Y=1.485 $X2=10.6 $Y2=2.31
r459 15 133 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.455
+ $Y=1.485 $X2=10.6 $Y2=1.63
r460 14 121 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=9.515
+ $Y=1.485 $X2=9.66 $Y2=2.31
r461 14 119 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.515
+ $Y=1.485 $X2=9.66 $Y2=1.63
r462 13 107 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.485 $X2=8.72 $Y2=2.31
r463 13 105 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.485 $X2=8.72 $Y2=1.63
r464 12 93 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=2.31
r465 12 91 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=1.63
r466 11 79 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=2.31
r467 11 77 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=1.63
r468 10 67 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=2.31
r469 10 65 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=1.63
r470 9 55 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=2.31
r471 9 53 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.63
r472 8 143 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=11.355
+ $Y=0.235 $X2=11.54 $Y2=0.4
r473 7 129 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=10.415
+ $Y=0.235 $X2=10.6 $Y2=0.4
r474 6 115 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=9.475
+ $Y=0.235 $X2=9.66 $Y2=0.4
r475 5 101 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=8.535
+ $Y=0.235 $X2=8.72 $Y2=0.4
r476 4 87 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=7.595
+ $Y=0.235 $X2=7.78 $Y2=0.4
r477 3 162 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=6.655
+ $Y=0.235 $X2=6.84 $Y2=0.4
r478 2 158 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=5.715
+ $Y=0.235 $X2=5.9 $Y2=0.4
r479 1 156 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFINV_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 44 46
+ 50 52 56 60 64 68 72 76 80 84 88 92 96 99 100 102 103 105 106 108 109 111 112
+ 114 115 117 118 120 121 123 124 126 127 128 162 163 166 169 172 175
r230 172 173 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r231 170 173 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r232 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r233 167 170 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r234 166 167 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r235 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r236 160 163 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r237 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r238 157 160 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.73 $Y2=0
r239 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r240 154 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r241 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r242 151 154 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r243 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r244 148 151 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r245 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r246 145 148 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r247 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r248 142 145 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r249 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r250 139 142 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r251 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r252 136 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r253 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r254 133 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r255 133 173 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.53 $Y2=0
r256 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r257 130 172 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0
+ $X2=2.61 $Y2=0
r258 130 132 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.695 $Y=0
+ $X2=3.45 $Y2=0
r259 128 167 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r260 128 175 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r261 126 159 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=11.925 $Y=0
+ $X2=11.73 $Y2=0
r262 126 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.925 $Y=0
+ $X2=12.01 $Y2=0
r263 125 162 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=12.095 $Y=0
+ $X2=12.19 $Y2=0
r264 125 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.095 $Y=0
+ $X2=12.01 $Y2=0
r265 123 156 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.985 $Y=0
+ $X2=10.81 $Y2=0
r266 123 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.985 $Y=0
+ $X2=11.07 $Y2=0
r267 122 159 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=11.155 $Y=0
+ $X2=11.73 $Y2=0
r268 122 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.155 $Y=0
+ $X2=11.07 $Y2=0
r269 120 153 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.045 $Y=0
+ $X2=9.89 $Y2=0
r270 120 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.045 $Y=0
+ $X2=10.13 $Y2=0
r271 119 156 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=10.215 $Y=0
+ $X2=10.81 $Y2=0
r272 119 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.215 $Y=0
+ $X2=10.13 $Y2=0
r273 117 150 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=9.105 $Y=0
+ $X2=8.97 $Y2=0
r274 117 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.105 $Y=0
+ $X2=9.19 $Y2=0
r275 116 153 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=9.275 $Y=0
+ $X2=9.89 $Y2=0
r276 116 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.275 $Y=0
+ $X2=9.19 $Y2=0
r277 114 147 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.165 $Y=0
+ $X2=8.05 $Y2=0
r278 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.165 $Y=0
+ $X2=8.25 $Y2=0
r279 113 150 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.335 $Y=0
+ $X2=8.97 $Y2=0
r280 113 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=0
+ $X2=8.25 $Y2=0
r281 111 144 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.225 $Y=0
+ $X2=7.13 $Y2=0
r282 111 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.225 $Y=0
+ $X2=7.31 $Y2=0
r283 110 147 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=7.395 $Y=0
+ $X2=8.05 $Y2=0
r284 110 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=0
+ $X2=7.31 $Y2=0
r285 108 141 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.285 $Y=0
+ $X2=6.21 $Y2=0
r286 108 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.285 $Y=0
+ $X2=6.37 $Y2=0
r287 107 144 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.455 $Y=0
+ $X2=7.13 $Y2=0
r288 107 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=0
+ $X2=6.37 $Y2=0
r289 105 138 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.29 $Y2=0
r290 105 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.43 $Y2=0
r291 104 141 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.515 $Y=0
+ $X2=6.21 $Y2=0
r292 104 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.515 $Y=0
+ $X2=5.43 $Y2=0
r293 102 135 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.37 $Y2=0
r294 102 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.49 $Y2=0
r295 101 138 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=4.575 $Y=0
+ $X2=5.29 $Y2=0
r296 101 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=0
+ $X2=4.49 $Y2=0
r297 99 132 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.465 $Y=0
+ $X2=3.45 $Y2=0
r298 99 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.55
+ $Y2=0
r299 98 135 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.635 $Y=0
+ $X2=4.37 $Y2=0
r300 98 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.55
+ $Y2=0
r301 94 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.01 $Y=0.085
+ $X2=12.01 $Y2=0
r302 94 96 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.01 $Y=0.085
+ $X2=12.01 $Y2=0.4
r303 90 124 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.07 $Y=0.085
+ $X2=11.07 $Y2=0
r304 90 92 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=11.07 $Y=0.085
+ $X2=11.07 $Y2=0.4
r305 86 121 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.13 $Y=0.085
+ $X2=10.13 $Y2=0
r306 86 88 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.13 $Y=0.085
+ $X2=10.13 $Y2=0.4
r307 82 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.19 $Y=0.085
+ $X2=9.19 $Y2=0
r308 82 84 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.19 $Y=0.085
+ $X2=9.19 $Y2=0.4
r309 78 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.25 $Y=0.085
+ $X2=8.25 $Y2=0
r310 78 80 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.25 $Y=0.085
+ $X2=8.25 $Y2=0.4
r311 74 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=0.085
+ $X2=7.31 $Y2=0
r312 74 76 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.31 $Y=0.085
+ $X2=7.31 $Y2=0.4
r313 70 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=0.085
+ $X2=6.37 $Y2=0
r314 70 72 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.37 $Y=0.085
+ $X2=6.37 $Y2=0.4
r315 66 106 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=0.085
+ $X2=5.43 $Y2=0
r316 66 68 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.43 $Y=0.085
+ $X2=5.43 $Y2=0.4
r317 62 103 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0
r318 62 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0.4
r319 58 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r320 58 60 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.4
r321 54 172 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r322 54 56 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.4
r323 53 169 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.67
+ $Y2=0
r324 52 172 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0 $X2=2.61
+ $Y2=0
r325 52 53 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.525 $Y=0
+ $X2=1.755 $Y2=0
r326 48 169 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r327 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.4
r328 47 166 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r329 46 169 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.67
+ $Y2=0
r330 46 47 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0
+ $X2=0.815 $Y2=0
r331 42 166 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r332 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.4
r333 13 96 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=11.875
+ $Y=0.235 $X2=12.01 $Y2=0.4
r334 12 92 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=10.885
+ $Y=0.235 $X2=11.07 $Y2=0.4
r335 11 88 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=0.235 $X2=10.13 $Y2=0.4
r336 10 84 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=9.005
+ $Y=0.235 $X2=9.19 $Y2=0.4
r337 9 80 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=8.065
+ $Y=0.235 $X2=8.25 $Y2=0.4
r338 8 76 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=7.125
+ $Y=0.235 $X2=7.31 $Y2=0.4
r339 7 72 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=6.185
+ $Y=0.235 $X2=6.37 $Y2=0.4
r340 6 68 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=5.245
+ $Y=0.235 $X2=5.43 $Y2=0.4
r341 5 64 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.49 $Y2=0.4
r342 4 60 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.4
r343 3 56 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.4
r344 2 50 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.4
r345 1 44 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

