* NGSPICE file created from sky130_fd_sc_hdll__a21boi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VPWR B1_N a_27_413# VPB phighvt w=420000u l=180000u
+  ad=5.355e+11p pd=4.23e+06u as=1.155e+11p ps=1.39e+06u
M1001 VPWR A1 a_338_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.75e+11p ps=5.15e+06u
M1002 VGND B1_N a_27_413# VNB nshort w=420000u l=150000u
+  ad=4.345e+11p pd=3.99e+06u as=1.533e+11p ps=1.57e+06u
M1003 a_434_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=2.665e+11p pd=2.12e+06u as=3.51e+11p ps=2.38e+06u
M1004 VGND A2 a_434_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y a_27_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_338_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_338_297# a_27_413# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.25e+11p ps=2.65e+06u
.ends

