* File: sky130_fd_sc_hdll__and4b_1.pxi.spice
* Created: Thu Aug 27 18:58:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND4B_1%A_N N_A_N_c_82_n N_A_N_c_83_n N_A_N_M1001_g
+ N_A_N_M1008_g A_N A_N N_A_N_c_81_n PM_SKY130_FD_SC_HDLL__AND4B_1%A_N
x_PM_SKY130_FD_SC_HDLL__AND4B_1%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1001_s
+ N_A_27_47#_c_116_n N_A_27_47#_c_124_n N_A_27_47#_c_125_n N_A_27_47#_M1006_g
+ N_A_27_47#_c_117_n N_A_27_47#_c_118_n N_A_27_47#_M1011_g N_A_27_47#_c_136_n
+ N_A_27_47#_c_126_n N_A_27_47#_c_119_n N_A_27_47#_c_120_n N_A_27_47#_c_127_n
+ N_A_27_47#_c_128_n N_A_27_47#_c_121_n N_A_27_47#_c_129_n N_A_27_47#_c_122_n
+ PM_SKY130_FD_SC_HDLL__AND4B_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND4B_1%B N_B_c_203_n N_B_c_204_n N_B_M1004_g
+ N_B_M1000_g B B B B N_B_c_202_n PM_SKY130_FD_SC_HDLL__AND4B_1%B
x_PM_SKY130_FD_SC_HDLL__AND4B_1%C N_C_c_247_n N_C_c_248_n N_C_M1009_g
+ N_C_M1002_g C C C C N_C_c_246_n PM_SKY130_FD_SC_HDLL__AND4B_1%C
x_PM_SKY130_FD_SC_HDLL__AND4B_1%D N_D_c_291_n N_D_c_292_n N_D_M1010_g
+ N_D_M1005_g D D D N_D_c_290_n PM_SKY130_FD_SC_HDLL__AND4B_1%D
x_PM_SKY130_FD_SC_HDLL__AND4B_1%A_213_413# N_A_213_413#_M1011_s
+ N_A_213_413#_M1006_d N_A_213_413#_M1009_d N_A_213_413#_c_333_n
+ N_A_213_413#_M1007_g N_A_213_413#_c_334_n N_A_213_413#_M1003_g
+ N_A_213_413#_c_335_n N_A_213_413#_c_339_n N_A_213_413#_c_340_n
+ N_A_213_413#_c_341_n N_A_213_413#_c_342_n N_A_213_413#_c_343_n
+ N_A_213_413#_c_348_n N_A_213_413#_c_344_n N_A_213_413#_c_345_n
+ N_A_213_413#_c_336_n PM_SKY130_FD_SC_HDLL__AND4B_1%A_213_413#
x_PM_SKY130_FD_SC_HDLL__AND4B_1%VPWR N_VPWR_M1001_d N_VPWR_M1004_d
+ N_VPWR_M1010_d N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n
+ VPWR N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_431_n N_VPWR_c_439_n
+ N_VPWR_c_440_n N_VPWR_c_441_n PM_SKY130_FD_SC_HDLL__AND4B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__AND4B_1%X N_X_M1003_d N_X_M1007_d N_X_c_494_n
+ N_X_c_492_n X X X N_X_c_493_n PM_SKY130_FD_SC_HDLL__AND4B_1%X
x_PM_SKY130_FD_SC_HDLL__AND4B_1%VGND N_VGND_M1008_d N_VGND_M1005_d VGND
+ N_VGND_c_516_n N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n
+ PM_SKY130_FD_SC_HDLL__AND4B_1%VGND
cc_1 VNB N_A_N_M1008_g 0.0399372f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A_N 0.017697f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A_N_c_81_n 0.0398594f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_27_47#_c_116_n 0.0431981f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_A_27_47#_c_117_n 0.0362928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_118_n 0.0169156f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_7 VNB N_A_27_47#_c_119_n 0.00740425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_120_n 0.00854299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_121_n 0.00315735f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_122_n 0.00235676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_M1000_g 0.0363534f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_12 VNB B 0.00981573f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_13 VNB N_B_c_202_n 0.0250337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_C_M1002_g 0.0297361f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_15 VNB C 0.00647762f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_16 VNB N_C_c_246_n 0.0239695f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_17 VNB N_D_M1005_g 0.0277765f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_18 VNB D 0.00923658f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_19 VNB N_D_c_290_n 0.0217962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_213_413#_c_333_n 0.0256657f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_21 VNB N_A_213_413#_c_334_n 0.0204561f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_213_413#_c_335_n 0.00873199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_213_413#_c_336_n 0.00295043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_431_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_492_n 0.0255948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_493_n 0.023848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_516_n 0.0151398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_517_n 0.0652024f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_29 VNB N_VGND_c_518_n 0.0231993f $X=-0.19 $Y=-0.24 $X2=0.267 $Y2=1.16
cc_30 VNB N_VGND_c_519_n 0.228833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_520_n 0.0113743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_N_c_82_n 0.0418932f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_33 VPB N_A_N_c_83_n 0.0258023f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_34 VPB A_N 0.0203025f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_35 VPB N_A_N_c_81_n 0.0102197f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_36 VPB N_A_27_47#_c_116_n 0.00382125f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_37 VPB N_A_27_47#_c_124_n 0.0357384f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_38 VPB N_A_27_47#_c_125_n 0.0244447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_126_n 0.00221628f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_127_n 0.00809874f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_128_n 0.00848141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_129_n 0.00946808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_122_n 4.77183e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_B_c_203_n 0.0299406f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_45 VPB N_B_c_204_n 0.025572f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_46 VPB B 0.00836374f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_47 VPB N_B_c_202_n 0.0197295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_C_c_247_n 0.0349738f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_49 VPB N_C_c_248_n 0.0245249f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_50 VPB C 0.00602051f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_51 VPB N_C_c_246_n 0.00339918f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_52 VPB N_D_c_291_n 0.0309521f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_53 VPB N_D_c_292_n 0.0224366f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_54 VPB D 0.00570973f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_55 VPB N_D_c_290_n 0.00318404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_213_413#_c_333_n 0.0285491f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_57 VPB N_A_213_413#_c_335_n 0.0117857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_213_413#_c_339_n 4.28953e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_213_413#_c_340_n 0.0245477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_213_413#_c_341_n 3.47697e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_213_413#_c_342_n 0.0043831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_213_413#_c_343_n 0.00116958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_213_413#_c_344_n 0.00207056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_213_413#_c_345_n 0.00615692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_213_413#_c_336_n 3.13322e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_432_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_433_n 0.0056146f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_68 VPB N_VPWR_c_434_n 0.0169709f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_69 VPB N_VPWR_c_435_n 0.00631622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_436_n 0.0151914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_437_n 0.0225084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_431_n 0.0487202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_439_n 0.00503031f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_440_n 0.0192631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_441_n 0.0137367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_X_c_494_n 0.00777218f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_77 VPB N_X_c_492_n 0.00999758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB X 0.035153f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_79 N_A_N_M1008_g N_A_27_47#_c_116_n 0.00859971f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_80 A_N N_A_27_47#_c_116_n 2.69498e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A_N_c_81_n N_A_27_47#_c_116_n 0.0210098f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_N_c_82_n N_A_27_47#_c_124_n 0.0124201f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_83 N_A_N_c_83_n N_A_27_47#_c_125_n 0.0240026f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_84 N_A_N_M1008_g N_A_27_47#_c_136_n 0.00482387f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_N_c_83_n N_A_27_47#_c_126_n 0.00605735f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_86 N_A_N_M1008_g N_A_27_47#_c_119_n 0.0173427f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_87 A_N N_A_27_47#_c_119_n 0.0082585f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_88 N_A_N_c_81_n N_A_27_47#_c_119_n 6.98058e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_89 A_N N_A_27_47#_c_120_n 0.0153899f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A_N_c_81_n N_A_27_47#_c_120_n 0.00135787f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_N_c_82_n N_A_27_47#_c_127_n 0.00922955f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_92 N_A_N_c_83_n N_A_27_47#_c_127_n 0.00977791f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_93 A_N N_A_27_47#_c_127_n 0.00829866f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_94 A_N N_A_27_47#_c_128_n 0.0162852f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A_N_c_81_n N_A_27_47#_c_128_n 6.55167e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_N_M1008_g N_A_27_47#_c_121_n 0.00396617f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_N_c_82_n N_A_27_47#_c_129_n 0.00660856f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_98 A_N N_A_27_47#_c_129_n 0.0211002f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_99 A_N N_A_27_47#_c_122_n 0.0210107f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A_N_c_81_n N_A_27_47#_c_122_n 0.00263949f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_N_M1008_g N_A_213_413#_c_335_n 0.00189887f $X=0.52 $Y=0.445 $X2=0
+ $Y2=0
cc_102 N_A_N_M1008_g N_A_213_413#_c_348_n 0.00162248f $X=0.52 $Y=0.445 $X2=0
+ $Y2=0
cc_103 N_A_N_c_83_n N_VPWR_c_432_n 0.0119443f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_104 N_A_N_c_83_n N_VPWR_c_436_n 0.00321743f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_105 N_A_N_c_83_n N_VPWR_c_431_n 0.00474836f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_106 N_A_N_M1008_g N_VGND_c_516_n 0.00199743f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_N_M1008_g N_VGND_c_519_n 0.00361213f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_N_M1008_g N_VGND_c_520_n 0.0124198f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_124_n N_B_c_203_n 0.00624609f $X=0.975 $Y=1.89 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_125_n N_B_c_204_n 0.0200768f $X=0.975 $Y=1.99 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_116_n N_B_M1000_g 0.0025596f $X=0.975 $Y=1.325 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_118_n N_B_M1000_g 0.0484094f $X=1.46 $Y=0.73 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_118_n B 0.00371347f $X=1.46 $Y=0.73 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_116_n N_B_c_202_n 0.00624609f $X=0.975 $Y=1.325 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_117_n N_B_c_202_n 0.00350435f $X=1.385 $Y=0.805 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_116_n N_A_213_413#_c_335_n 0.0100428f $X=0.975 $Y=1.325
+ $X2=0 $Y2=0
cc_117 N_A_27_47#_c_117_n N_A_213_413#_c_335_n 0.0142632f $X=1.385 $Y=0.805
+ $X2=0 $Y2=0
cc_118 N_A_27_47#_c_118_n N_A_213_413#_c_335_n 0.00265874f $X=1.46 $Y=0.73 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_c_119_n N_A_213_413#_c_335_n 0.00831715f $X=0.68 $Y=0.74 $X2=0
+ $Y2=0
cc_120 N_A_27_47#_c_127_n N_A_213_413#_c_335_n 0.00150574f $X=0.68 $Y=1.93 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_c_121_n N_A_213_413#_c_335_n 0.00750968f $X=0.765 $Y=0.995
+ $X2=0 $Y2=0
cc_122 N_A_27_47#_c_129_n N_A_213_413#_c_335_n 0.0236515f $X=0.765 $Y=1.845
+ $X2=0 $Y2=0
cc_123 N_A_27_47#_c_122_n N_A_213_413#_c_335_n 0.0243143f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_c_125_n N_A_213_413#_c_339_n 0.00602918f $X=0.975 $Y=1.99
+ $X2=0 $Y2=0
cc_125 N_A_27_47#_c_117_n N_A_213_413#_c_348_n 0.00225284f $X=1.385 $Y=0.805
+ $X2=0 $Y2=0
cc_126 N_A_27_47#_c_124_n N_A_213_413#_c_344_n 0.00135107f $X=0.975 $Y=1.89
+ $X2=0 $Y2=0
cc_127 N_A_27_47#_c_125_n N_A_213_413#_c_344_n 0.00120221f $X=0.975 $Y=1.99
+ $X2=0 $Y2=0
cc_128 N_A_27_47#_c_127_n N_A_213_413#_c_344_n 0.00789642f $X=0.68 $Y=1.93 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_125_n N_VPWR_c_432_n 0.00886721f $X=0.975 $Y=1.99 $X2=0
+ $Y2=0
cc_130 N_A_27_47#_c_126_n N_VPWR_c_432_n 0.0201996f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_131 N_A_27_47#_c_127_n N_VPWR_c_432_n 0.022702f $X=0.68 $Y=1.93 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_126_n N_VPWR_c_436_n 0.0120835f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_127_n N_VPWR_c_436_n 0.00247264f $X=0.68 $Y=1.93 $X2=0 $Y2=0
cc_134 N_A_27_47#_M1001_s N_VPWR_c_431_n 0.00369267f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_135 N_A_27_47#_c_125_n N_VPWR_c_431_n 0.0116975f $X=0.975 $Y=1.99 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_126_n N_VPWR_c_431_n 0.00664644f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_127_n N_VPWR_c_431_n 0.00541564f $X=0.68 $Y=1.93 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_125_n N_VPWR_c_440_n 0.00682361f $X=0.975 $Y=1.99 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_c_125_n N_VPWR_c_441_n 9.78895e-19 $X=0.975 $Y=1.99 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_c_119_n N_VGND_M1008_d 0.00183923f $X=0.68 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A_27_47#_c_136_n N_VGND_c_516_n 0.0120098f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_119_n N_VGND_c_516_n 0.00283814f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_116_n N_VGND_c_517_n 0.00441617f $X=0.975 $Y=1.325 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_c_117_n N_VGND_c_517_n 6.44498e-19 $X=1.385 $Y=0.805 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_c_118_n N_VGND_c_517_n 0.00585385f $X=1.46 $Y=0.73 $X2=0 $Y2=0
cc_146 N_A_27_47#_M1008_s N_VGND_c_519_n 0.00416008f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_c_116_n N_VGND_c_519_n 0.00608612f $X=0.975 $Y=1.325 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_118_n N_VGND_c_519_n 0.0119273f $X=1.46 $Y=0.73 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_136_n N_VGND_c_519_n 0.00663203f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_119_n N_VGND_c_519_n 0.00589722f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_116_n N_VGND_c_520_n 0.00102845f $X=0.975 $Y=1.325 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_118_n N_VGND_c_520_n 0.0028078f $X=1.46 $Y=0.73 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_136_n N_VGND_c_520_n 0.0157109f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_119_n N_VGND_c_520_n 0.021213f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_122_n N_VGND_c_520_n 0.00157757f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_156 N_B_c_203_n N_C_c_247_n 0.00406841f $X=1.585 $Y=1.89 $X2=0 $Y2=0
cc_157 B N_C_c_247_n 0.00160196f $X=1.88 $Y=0.425 $X2=0 $Y2=0
cc_158 N_B_c_202_n N_C_c_247_n 0.00322919f $X=1.82 $Y=1.3 $X2=0 $Y2=0
cc_159 N_B_c_204_n N_C_c_248_n 0.00758807f $X=1.585 $Y=1.99 $X2=0 $Y2=0
cc_160 N_B_M1000_g N_C_M1002_g 0.0198244f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_161 B N_C_M1002_g 0.00210655f $X=1.88 $Y=0.425 $X2=0 $Y2=0
cc_162 N_B_c_203_n C 3.71228e-19 $X=1.585 $Y=1.89 $X2=0 $Y2=0
cc_163 N_B_M1000_g C 0.00155379f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_164 B C 0.106143f $X=1.88 $Y=0.425 $X2=0 $Y2=0
cc_165 N_B_c_202_n C 3.01928e-19 $X=1.82 $Y=1.3 $X2=0 $Y2=0
cc_166 N_B_M1000_g N_C_c_246_n 0.00901707f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_167 B N_C_c_246_n 0.00283171f $X=1.88 $Y=0.425 $X2=0 $Y2=0
cc_168 N_B_M1000_g N_A_213_413#_c_335_n 0.00105034f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_169 B N_A_213_413#_c_335_n 0.059952f $X=1.88 $Y=0.425 $X2=0 $Y2=0
cc_170 N_B_c_202_n N_A_213_413#_c_335_n 0.0100282f $X=1.82 $Y=1.3 $X2=0 $Y2=0
cc_171 N_B_c_204_n N_A_213_413#_c_339_n 0.00650398f $X=1.585 $Y=1.99 $X2=0 $Y2=0
cc_172 N_B_c_203_n N_A_213_413#_c_340_n 0.0092494f $X=1.585 $Y=1.89 $X2=0 $Y2=0
cc_173 N_B_c_204_n N_A_213_413#_c_340_n 0.0123091f $X=1.585 $Y=1.99 $X2=0 $Y2=0
cc_174 B N_A_213_413#_c_340_n 0.0386926f $X=1.88 $Y=0.425 $X2=0 $Y2=0
cc_175 N_B_c_202_n N_A_213_413#_c_340_n 8.64548e-19 $X=1.82 $Y=1.3 $X2=0 $Y2=0
cc_176 N_B_c_204_n N_VPWR_c_432_n 9.36967e-19 $X=1.585 $Y=1.99 $X2=0 $Y2=0
cc_177 N_B_c_204_n N_VPWR_c_431_n 0.00560402f $X=1.585 $Y=1.99 $X2=0 $Y2=0
cc_178 N_B_c_204_n N_VPWR_c_440_n 0.00462245f $X=1.585 $Y=1.99 $X2=0 $Y2=0
cc_179 N_B_c_204_n N_VPWR_c_441_n 0.00979504f $X=1.585 $Y=1.99 $X2=0 $Y2=0
cc_180 N_B_M1000_g N_VGND_c_517_n 0.0038979f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_181 B N_VGND_c_517_n 0.0140961f $X=1.88 $Y=0.425 $X2=0 $Y2=0
cc_182 N_B_M1000_g N_VGND_c_519_n 0.00579689f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_183 B N_VGND_c_519_n 0.0159955f $X=1.88 $Y=0.425 $X2=0 $Y2=0
cc_184 B A_307_47# 0.00271511f $X=1.88 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_185 B A_379_47# 0.00582975f $X=1.88 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_186 N_C_c_247_n N_D_c_291_n 0.0141958f $X=2.445 $Y=1.89 $X2=0 $Y2=0
cc_187 C N_D_c_291_n 0.00110946f $X=2.35 $Y=0.425 $X2=0 $Y2=0
cc_188 N_C_c_248_n N_D_c_292_n 0.0235293f $X=2.445 $Y=1.99 $X2=0 $Y2=0
cc_189 N_C_M1002_g N_D_M1005_g 0.0297243f $X=2.47 $Y=0.445 $X2=0 $Y2=0
cc_190 C N_D_M1005_g 0.00536477f $X=2.35 $Y=0.425 $X2=0 $Y2=0
cc_191 N_C_c_247_n D 0.00109644f $X=2.445 $Y=1.89 $X2=0 $Y2=0
cc_192 N_C_M1002_g D 0.0010179f $X=2.47 $Y=0.445 $X2=0 $Y2=0
cc_193 C D 0.0827536f $X=2.35 $Y=0.425 $X2=0 $Y2=0
cc_194 N_C_c_246_n D 3.62814e-19 $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_195 C N_D_c_290_n 0.00191353f $X=2.35 $Y=0.425 $X2=0 $Y2=0
cc_196 N_C_c_246_n N_D_c_290_n 0.0175765f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_197 N_C_c_247_n N_A_213_413#_c_340_n 0.00348299f $X=2.445 $Y=1.89 $X2=0 $Y2=0
cc_198 N_C_c_248_n N_A_213_413#_c_340_n 0.0122757f $X=2.445 $Y=1.99 $X2=0 $Y2=0
cc_199 C N_A_213_413#_c_340_n 0.0216858f $X=2.35 $Y=0.425 $X2=0 $Y2=0
cc_200 N_C_c_246_n N_A_213_413#_c_340_n 0.0013504f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_201 N_C_c_248_n N_A_213_413#_c_341_n 0.00454072f $X=2.445 $Y=1.99 $X2=0 $Y2=0
cc_202 N_C_c_248_n N_VPWR_c_434_n 0.00462245f $X=2.445 $Y=1.99 $X2=0 $Y2=0
cc_203 N_C_c_248_n N_VPWR_c_431_n 0.00533157f $X=2.445 $Y=1.99 $X2=0 $Y2=0
cc_204 N_C_c_248_n N_VPWR_c_441_n 0.00955087f $X=2.445 $Y=1.99 $X2=0 $Y2=0
cc_205 N_C_M1002_g N_VGND_c_517_n 0.00599743f $X=2.47 $Y=0.445 $X2=0 $Y2=0
cc_206 C N_VGND_c_517_n 0.00974409f $X=2.35 $Y=0.425 $X2=0 $Y2=0
cc_207 N_C_M1002_g N_VGND_c_519_n 0.006162f $X=2.47 $Y=0.445 $X2=0 $Y2=0
cc_208 C N_VGND_c_519_n 0.00934269f $X=2.35 $Y=0.425 $X2=0 $Y2=0
cc_209 C A_379_47# 0.00237115f $X=2.35 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_210 C A_509_47# 0.00326822f $X=2.35 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_211 N_D_c_291_n N_A_213_413#_c_333_n 0.0223345f $X=2.95 $Y=1.89 $X2=0 $Y2=0
cc_212 N_D_c_292_n N_A_213_413#_c_333_n 0.00916453f $X=2.95 $Y=1.99 $X2=0 $Y2=0
cc_213 D N_A_213_413#_c_333_n 0.00188283f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_214 N_D_c_290_n N_A_213_413#_c_333_n 0.0160273f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_215 N_D_M1005_g N_A_213_413#_c_334_n 0.0207522f $X=2.975 $Y=0.445 $X2=0 $Y2=0
cc_216 D N_A_213_413#_c_334_n 0.00266835f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_217 N_D_c_292_n N_A_213_413#_c_341_n 0.00476323f $X=2.95 $Y=1.99 $X2=0 $Y2=0
cc_218 N_D_c_291_n N_A_213_413#_c_342_n 0.00339951f $X=2.95 $Y=1.89 $X2=0 $Y2=0
cc_219 N_D_c_292_n N_A_213_413#_c_342_n 0.0114971f $X=2.95 $Y=1.99 $X2=0 $Y2=0
cc_220 D N_A_213_413#_c_342_n 0.020514f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_221 N_D_c_291_n N_A_213_413#_c_343_n 0.00491721f $X=2.95 $Y=1.89 $X2=0 $Y2=0
cc_222 D N_A_213_413#_c_343_n 0.0287528f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_223 D N_A_213_413#_c_345_n 0.00124698f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_224 N_D_c_290_n N_A_213_413#_c_345_n 2.25801e-19 $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_225 D N_A_213_413#_c_336_n 0.0269012f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_226 N_D_c_290_n N_A_213_413#_c_336_n 0.0010463f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_227 N_D_c_292_n N_VPWR_c_433_n 0.00319717f $X=2.95 $Y=1.99 $X2=0 $Y2=0
cc_228 N_D_c_292_n N_VPWR_c_434_n 0.00523815f $X=2.95 $Y=1.99 $X2=0 $Y2=0
cc_229 N_D_c_292_n N_VPWR_c_431_n 0.00694721f $X=2.95 $Y=1.99 $X2=0 $Y2=0
cc_230 N_D_c_292_n N_VPWR_c_441_n 0.00108425f $X=2.95 $Y=1.99 $X2=0 $Y2=0
cc_231 D N_X_c_492_n 0.0059135f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_232 N_D_M1005_g N_X_c_493_n 8.59019e-19 $X=2.975 $Y=0.445 $X2=0 $Y2=0
cc_233 D N_X_c_493_n 0.00548267f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_234 N_D_M1005_g N_VGND_c_517_n 0.0152989f $X=2.975 $Y=0.445 $X2=0 $Y2=0
cc_235 D N_VGND_c_517_n 0.0103531f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_236 N_D_M1005_g N_VGND_c_519_n 0.00249993f $X=2.975 $Y=0.445 $X2=0 $Y2=0
cc_237 D N_VGND_c_519_n 0.0052956f $X=2.84 $Y=0.765 $X2=0 $Y2=0
cc_238 N_A_213_413#_c_342_n N_VPWR_M1010_d 0.00631886f $X=3.245 $Y=1.96 $X2=0
+ $Y2=0
cc_239 N_A_213_413#_c_343_n N_VPWR_M1010_d 0.00388543f $X=3.33 $Y=1.875 $X2=0
+ $Y2=0
cc_240 N_A_213_413#_c_339_n N_VPWR_c_432_n 0.012863f $X=1.285 $Y=2.3 $X2=0 $Y2=0
cc_241 N_A_213_413#_c_333_n N_VPWR_c_433_n 0.00329263f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_242 N_A_213_413#_c_342_n N_VPWR_c_433_n 0.01959f $X=3.245 $Y=1.96 $X2=0 $Y2=0
cc_243 N_A_213_413#_c_340_n N_VPWR_c_434_n 0.00397113f $X=2.63 $Y=1.96 $X2=0
+ $Y2=0
cc_244 N_A_213_413#_c_341_n N_VPWR_c_434_n 0.0116919f $X=2.715 $Y=2.3 $X2=0
+ $Y2=0
cc_245 N_A_213_413#_c_342_n N_VPWR_c_434_n 0.00401756f $X=3.245 $Y=1.96 $X2=0
+ $Y2=0
cc_246 N_A_213_413#_c_333_n N_VPWR_c_437_n 0.00681844f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_247 N_A_213_413#_c_342_n N_VPWR_c_437_n 3.57522e-19 $X=3.245 $Y=1.96 $X2=0
+ $Y2=0
cc_248 N_A_213_413#_M1006_d N_VPWR_c_431_n 0.00847461f $X=1.065 $Y=2.065 $X2=0
+ $Y2=0
cc_249 N_A_213_413#_M1009_d N_VPWR_c_431_n 0.00322491f $X=2.535 $Y=2.065 $X2=0
+ $Y2=0
cc_250 N_A_213_413#_c_333_n N_VPWR_c_431_n 0.0130776f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_251 N_A_213_413#_c_339_n N_VPWR_c_431_n 0.00646998f $X=1.285 $Y=2.3 $X2=0
+ $Y2=0
cc_252 N_A_213_413#_c_340_n N_VPWR_c_431_n 0.0162265f $X=2.63 $Y=1.96 $X2=0
+ $Y2=0
cc_253 N_A_213_413#_c_341_n N_VPWR_c_431_n 0.00644606f $X=2.715 $Y=2.3 $X2=0
+ $Y2=0
cc_254 N_A_213_413#_c_342_n N_VPWR_c_431_n 0.00821332f $X=3.245 $Y=1.96 $X2=0
+ $Y2=0
cc_255 N_A_213_413#_c_339_n N_VPWR_c_440_n 0.0118139f $X=1.285 $Y=2.3 $X2=0
+ $Y2=0
cc_256 N_A_213_413#_c_340_n N_VPWR_c_440_n 0.00447575f $X=2.63 $Y=1.96 $X2=0
+ $Y2=0
cc_257 N_A_213_413#_c_339_n N_VPWR_c_441_n 0.0126549f $X=1.285 $Y=2.3 $X2=0
+ $Y2=0
cc_258 N_A_213_413#_c_340_n N_VPWR_c_441_n 0.0483995f $X=2.63 $Y=1.96 $X2=0
+ $Y2=0
cc_259 N_A_213_413#_c_341_n N_VPWR_c_441_n 0.0137885f $X=2.715 $Y=2.3 $X2=0
+ $Y2=0
cc_260 N_A_213_413#_c_333_n N_X_c_494_n 0.0119045f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_213_413#_c_343_n N_X_c_494_n 0.0231758f $X=3.33 $Y=1.875 $X2=0 $Y2=0
cc_262 N_A_213_413#_c_333_n N_X_c_492_n 0.0016986f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_213_413#_c_334_n N_X_c_492_n 0.0129509f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A_213_413#_c_343_n N_X_c_492_n 0.00801916f $X=3.33 $Y=1.875 $X2=0 $Y2=0
cc_265 N_A_213_413#_c_336_n N_X_c_492_n 0.0233841f $X=3.45 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_213_413#_c_342_n X 0.0115472f $X=3.245 $Y=1.96 $X2=0 $Y2=0
cc_267 N_A_213_413#_c_334_n N_X_c_493_n 0.0128779f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_213_413#_c_336_n N_X_c_493_n 9.98652e-19 $X=3.45 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_213_413#_c_333_n N_VGND_c_517_n 6.13671e-19 $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_270 N_A_213_413#_c_334_n N_VGND_c_517_n 0.00594971f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_271 N_A_213_413#_c_348_n N_VGND_c_517_n 0.0143957f $X=1.25 $Y=0.42 $X2=0
+ $Y2=0
cc_272 N_A_213_413#_c_336_n N_VGND_c_517_n 0.00376991f $X=3.45 $Y=1.16 $X2=0
+ $Y2=0
cc_273 N_A_213_413#_c_334_n N_VGND_c_518_n 0.00491742f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_274 N_A_213_413#_M1011_s N_VGND_c_519_n 0.00244967f $X=1.125 $Y=0.235 $X2=0
+ $Y2=0
cc_275 N_A_213_413#_c_334_n N_VGND_c_519_n 0.00974775f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_276 N_A_213_413#_c_348_n N_VGND_c_519_n 0.00874023f $X=1.25 $Y=0.42 $X2=0
+ $Y2=0
cc_277 N_A_213_413#_c_348_n N_VGND_c_520_n 0.0130177f $X=1.25 $Y=0.42 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_431_n N_X_M1007_d 0.00430086f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_c_437_n X 0.0253796f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_c_431_n X 0.0137872f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_281 N_X_c_493_n N_VGND_c_517_n 0.0137469f $X=3.72 $Y=0.38 $X2=0 $Y2=0
cc_282 N_X_c_493_n N_VGND_c_518_n 0.0247744f $X=3.72 $Y=0.38 $X2=0 $Y2=0
cc_283 N_X_M1003_d N_VGND_c_519_n 0.00211564f $X=3.585 $Y=0.235 $X2=0 $Y2=0
cc_284 N_X_c_493_n N_VGND_c_519_n 0.0174216f $X=3.72 $Y=0.38 $X2=0 $Y2=0
cc_285 N_VGND_c_519_n A_307_47# 0.00664531f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_286 N_VGND_c_519_n A_379_47# 0.0103144f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_287 N_VGND_c_519_n A_509_47# 0.00937177f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
