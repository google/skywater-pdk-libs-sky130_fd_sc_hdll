* File: sky130_fd_sc_hdll__clkinvlp_2.pxi.spice
* Created: Thu Aug 27 19:03:10 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKINVLP_2%A N_A_M1001_g N_A_c_27_n N_A_M1002_g
+ N_A_c_28_n N_A_M1003_g N_A_c_30_n N_A_M1000_g N_A_c_31_n A A N_A_c_32_n
+ N_A_c_33_n PM_SKY130_FD_SC_HDLL__CLKINVLP_2%A
x_PM_SKY130_FD_SC_HDLL__CLKINVLP_2%VPWR N_VPWR_M1001_d N_VPWR_M1003_d
+ N_VPWR_c_67_n N_VPWR_c_68_n N_VPWR_c_69_n N_VPWR_c_70_n VPWR N_VPWR_c_71_n
+ N_VPWR_c_66_n PM_SKY130_FD_SC_HDLL__CLKINVLP_2%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKINVLP_2%Y N_Y_M1000_d N_Y_M1001_s Y Y Y Y N_Y_c_88_n
+ PM_SKY130_FD_SC_HDLL__CLKINVLP_2%Y
x_PM_SKY130_FD_SC_HDLL__CLKINVLP_2%VGND N_VGND_M1002_s N_VGND_c_109_n
+ N_VGND_c_110_n N_VGND_c_111_n VGND N_VGND_c_112_n N_VGND_c_113_n
+ PM_SKY130_FD_SC_HDLL__CLKINVLP_2%VGND
cc_1 VNB N_A_c_27_n 0.0223343f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=0.995
cc_2 VNB N_A_c_28_n 0.0124832f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.082
cc_3 VNB N_A_M1003_g 0.0119835f $X=-0.19 $Y=-0.24 $X2=1.135 $Y2=1.985
cc_4 VNB N_A_c_30_n 0.0234789f $X=-0.19 $Y=-0.24 $X2=1.185 $Y2=0.995
cc_5 VNB N_A_c_31_n 0.0146011f $X=-0.19 $Y=-0.24 $X2=1.135 $Y2=1.082
cc_6 VNB N_A_c_32_n 0.0517951f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_7 VNB N_A_c_33_n 0.00936522f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_8 VNB N_VPWR_c_66_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.372 $Y2=1.19
cc_9 VNB Y 0.00192599f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=0.61
cc_10 VNB N_Y_c_88_n 0.0228142f $X=-0.19 $Y=-0.24 $X2=0.372 $Y2=1.16
cc_11 VNB N_VGND_c_109_n 0.0238309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_110_n 0.0115308f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=0.61
cc_13 VNB N_VGND_c_111_n 0.00572238f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.082
cc_14 VNB N_VGND_c_112_n 0.0343864f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_15 VNB N_VGND_c_113_n 0.145349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VPB N_A_M1001_g 0.0291172f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.985
cc_17 VPB N_A_M1003_g 0.0333679f $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.985
cc_18 VPB N_A_c_32_n 0.0108532f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_19 VPB N_A_c_33_n 0.015867f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_20 VPB N_VPWR_c_67_n 0.0143479f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=0.995
cc_21 VPB N_VPWR_c_68_n 0.00228555f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=0.61
cc_22 VPB N_VPWR_c_69_n 0.0129807f $X=-0.19 $Y=1.305 $X2=0.75 $Y2=1.082
cc_23 VPB N_VPWR_c_70_n 0.0544286f $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.985
cc_24 VPB N_VPWR_c_71_n 0.0217884f $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.082
cc_25 VPB N_VPWR_c_66_n 0.0502546f $X=-0.19 $Y=1.305 $X2=0.372 $Y2=1.19
cc_26 VPB Y 0.00130058f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=0.61
cc_27 N_A_c_33_n N_VPWR_M1001_d 0.00456301f $X=0.515 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_28 N_A_M1001_g N_VPWR_c_68_n 0.0199547f $X=0.605 $Y=1.985 $X2=0 $Y2=0
cc_29 N_A_M1003_g N_VPWR_c_68_n 0.0013387f $X=1.135 $Y=1.985 $X2=0 $Y2=0
cc_30 N_A_c_32_n N_VPWR_c_68_n 8.71838e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_31 N_A_c_33_n N_VPWR_c_68_n 0.0239572f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_32 N_A_M1003_g N_VPWR_c_70_n 0.0270796f $X=1.135 $Y=1.985 $X2=0 $Y2=0
cc_33 N_A_M1001_g N_VPWR_c_71_n 0.00695524f $X=0.605 $Y=1.985 $X2=0 $Y2=0
cc_34 N_A_M1003_g N_VPWR_c_71_n 0.00648274f $X=1.135 $Y=1.985 $X2=0 $Y2=0
cc_35 N_A_M1001_g N_VPWR_c_66_n 0.0113395f $X=0.605 $Y=1.985 $X2=0 $Y2=0
cc_36 N_A_M1003_g N_VPWR_c_66_n 0.00972069f $X=1.135 $Y=1.985 $X2=0 $Y2=0
cc_37 N_A_c_27_n Y 0.00406934f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_38 N_A_c_28_n Y 0.0119713f $X=1.01 $Y=1.082 $X2=0 $Y2=0
cc_39 N_A_M1003_g Y 0.0510311f $X=1.135 $Y=1.985 $X2=0 $Y2=0
cc_40 N_A_c_30_n Y 0.0167373f $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_41 N_A_c_31_n Y 0.0111062f $X=1.135 $Y=1.082 $X2=0 $Y2=0
cc_42 N_A_c_32_n Y 0.0038034f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_43 N_A_c_33_n Y 0.0439713f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_44 N_A_c_27_n N_Y_c_88_n 0.00243717f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_45 N_A_c_28_n N_Y_c_88_n 6.96208e-19 $X=1.01 $Y=1.082 $X2=0 $Y2=0
cc_46 N_A_c_30_n N_Y_c_88_n 0.0158122f $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_47 N_A_c_27_n N_VGND_c_109_n 0.0108318f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_48 N_A_c_30_n N_VGND_c_109_n 8.79064e-19 $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_49 N_A_c_32_n N_VGND_c_109_n 0.00206864f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_50 N_A_c_33_n N_VGND_c_109_n 0.0177327f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_51 N_A_c_27_n N_VGND_c_112_n 0.00440246f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_52 N_A_c_30_n N_VGND_c_112_n 0.00306316f $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_53 N_A_c_27_n N_VGND_c_113_n 0.00842314f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A_c_30_n N_VGND_c_113_n 0.00443248f $X=1.185 $Y=0.995 $X2=0 $Y2=0
cc_55 N_VPWR_c_66_n N_Y_M1001_s 0.00419524f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_56 N_VPWR_c_70_n Y 0.0780892f $X=1.5 $Y=1.63 $X2=0 $Y2=0
cc_57 N_VPWR_c_71_n Y 0.0290092f $X=1.405 $Y=2.715 $X2=0 $Y2=0
cc_58 N_VPWR_c_66_n Y 0.0160096f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_59 N_Y_c_88_n N_VGND_c_109_n 0.0169367f $X=1.4 $Y=0.58 $X2=0 $Y2=0
cc_60 N_Y_c_88_n N_VGND_c_112_n 0.0375636f $X=1.4 $Y=0.58 $X2=0 $Y2=0
cc_61 N_Y_c_88_n N_VGND_c_113_n 0.0272658f $X=1.4 $Y=0.58 $X2=0 $Y2=0
cc_62 Y A_150_67# 0.00116151f $X=1.055 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_63 N_Y_c_88_n A_150_67# 0.00345979f $X=1.4 $Y=0.58 $X2=-0.19 $Y2=-0.24
