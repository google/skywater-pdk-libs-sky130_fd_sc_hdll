* File: sky130_fd_sc_hdll__or4bb_2.pxi.spice
* Created: Thu Aug 27 19:25:38 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%C_N N_C_N_c_99_n N_C_N_c_100_n N_C_N_M1010_g
+ N_C_N_M1001_g C_N C_N N_C_N_c_96_n N_C_N_c_97_n N_C_N_c_98_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_2%C_N
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%D_N N_D_N_c_129_n N_D_N_M1003_g N_D_N_c_130_n
+ N_D_N_M1011_g D_N D_N PM_SKY130_FD_SC_HDLL__OR4BB_2%D_N
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%A_216_93# N_A_216_93#_M1003_d
+ N_A_216_93#_M1011_d N_A_216_93#_c_169_n N_A_216_93#_c_170_n
+ N_A_216_93#_M1008_g N_A_216_93#_M1002_g N_A_216_93#_c_171_n
+ N_A_216_93#_c_164_n N_A_216_93#_c_165_n N_A_216_93#_c_166_n
+ N_A_216_93#_c_167_n N_A_216_93#_c_168_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_2%A_216_93#
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%A_27_410# N_A_27_410#_M1001_s
+ N_A_27_410#_M1010_s N_A_27_410#_M1015_g N_A_27_410#_c_233_n
+ N_A_27_410#_M1006_g N_A_27_410#_c_234_n N_A_27_410#_c_239_n
+ N_A_27_410#_c_240_n N_A_27_410#_c_241_n N_A_27_410#_c_242_n
+ N_A_27_410#_c_243_n N_A_27_410#_c_235_n N_A_27_410#_c_236_n
+ N_A_27_410#_c_245_n PM_SKY130_FD_SC_HDLL__OR4BB_2%A_27_410#
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%B N_B_c_326_n N_B_c_327_n N_B_c_329_n
+ N_B_c_330_n N_B_M1009_g N_B_M1012_g N_B_c_328_n B B
+ PM_SKY130_FD_SC_HDLL__OR4BB_2%B
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%A N_A_c_369_n N_A_M1000_g N_A_M1007_g A
+ N_A_c_371_n A PM_SKY130_FD_SC_HDLL__OR4BB_2%A
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%A_336_413# N_A_336_413#_M1002_d
+ N_A_336_413#_M1012_d N_A_336_413#_M1008_s N_A_336_413#_c_417_n
+ N_A_336_413#_M1004_g N_A_336_413#_c_408_n N_A_336_413#_M1013_g
+ N_A_336_413#_c_418_n N_A_336_413#_M1005_g N_A_336_413#_c_409_n
+ N_A_336_413#_M1014_g N_A_336_413#_c_419_n N_A_336_413#_c_432_n
+ N_A_336_413#_c_420_n N_A_336_413#_c_410_n N_A_336_413#_c_411_n
+ N_A_336_413#_c_421_n N_A_336_413#_c_429_n N_A_336_413#_c_521_p
+ N_A_336_413#_c_412_n N_A_336_413#_c_466_n N_A_336_413#_c_422_n
+ N_A_336_413#_c_413_n N_A_336_413#_c_423_n N_A_336_413#_c_414_n
+ N_A_336_413#_c_415_n N_A_336_413#_c_416_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_2%A_336_413#
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%VPWR N_VPWR_M1010_d N_VPWR_M1000_d
+ N_VPWR_M1005_d N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n N_VPWR_c_541_n
+ N_VPWR_c_542_n N_VPWR_c_543_n VPWR N_VPWR_c_544_n N_VPWR_c_545_n
+ N_VPWR_c_546_n N_VPWR_c_537_n PM_SKY130_FD_SC_HDLL__OR4BB_2%VPWR
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%X N_X_M1013_s N_X_M1004_s N_X_c_605_n
+ N_X_c_607_n N_X_c_603_n X PM_SKY130_FD_SC_HDLL__OR4BB_2%X
x_PM_SKY130_FD_SC_HDLL__OR4BB_2%VGND N_VGND_M1001_d N_VGND_M1002_s
+ N_VGND_M1015_d N_VGND_M1007_d N_VGND_M1014_d N_VGND_c_629_n N_VGND_c_630_n
+ N_VGND_c_631_n N_VGND_c_632_n N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n
+ N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n N_VGND_c_640_n
+ VGND N_VGND_c_641_n N_VGND_c_642_n N_VGND_c_643_n VGND
+ PM_SKY130_FD_SC_HDLL__OR4BB_2%VGND
cc_1 VNB N_C_N_c_96_n 0.0258704f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_2 VNB N_C_N_c_97_n 0.00825123f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_3 VNB N_C_N_c_98_n 0.0208838f $X=-0.19 $Y=-0.24 $X2=0.547 $Y2=0.995
cc_4 VNB N_D_N_c_129_n 0.019134f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_5 VNB N_D_N_c_130_n 0.0304902f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.26
cc_6 VNB D_N 0.0023568f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.675
cc_7 VNB N_A_216_93#_M1002_g 0.0343207f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_8 VNB N_A_216_93#_c_164_n 0.00470982f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_216_93#_c_165_n 7.21544e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_216_93#_c_166_n 0.0128829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_216_93#_c_167_n 0.00175f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_216_93#_c_168_n 0.0379272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_410#_M1015_g 0.0275893f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_14 VNB N_A_27_410#_c_233_n 0.0252977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_410#_c_234_n 0.0224941f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_16 VNB N_A_27_410#_c_235_n 6.93211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_410#_c_236_n 0.0187913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_c_326_n 0.00670451f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_19 VNB N_B_c_327_n 0.0210422f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.875
cc_20 VNB N_B_c_328_n 0.0158925f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.445
cc_21 VNB N_A_c_369_n 0.022998f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_22 VNB N_A_M1007_g 0.0293024f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.995
cc_23 VNB N_A_c_371_n 0.00453319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_336_413#_c_408_n 0.0176571f $X=-0.19 $Y=-0.24 $X2=0.547 $Y2=1.16
cc_25 VNB N_A_336_413#_c_409_n 0.0212176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_336_413#_c_410_n 0.0129372f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_336_413#_c_411_n 0.0047498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_336_413#_c_412_n 0.00328923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_336_413#_c_413_n 0.00149272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_336_413#_c_414_n 0.00260241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_336_413#_c_415_n 0.0018431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_336_413#_c_416_n 0.0526882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_537_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_603_n 8.19802e-19 $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_35 VNB N_VGND_c_629_n 0.015125f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_36 VNB N_VGND_c_630_n 0.020554f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.19
cc_37 VNB N_VGND_c_631_n 0.0119755f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_632_n 0.00206109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_633_n 0.0131265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_634_n 0.00870713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_635_n 0.0226869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_636_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_637_n 0.0149555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_638_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_639_n 0.00973217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_640_n 0.0135819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_641_n 0.021207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_642_n 0.00718038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_643_n 0.28542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VPB N_C_N_c_99_n 0.0336404f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.875
cc_51 VPB N_C_N_c_100_n 0.0286094f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.975
cc_52 VPB N_C_N_c_96_n 0.00432955f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_53 VPB N_C_N_c_97_n 0.0024706f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_54 VPB N_D_N_c_130_n 0.0315127f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_55 VPB D_N 5.16383e-19 $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.675
cc_56 VPB N_A_216_93#_c_169_n 0.0386139f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.675
cc_57 VPB N_A_216_93#_c_170_n 0.0307681f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_58 VPB N_A_216_93#_c_171_n 0.00893983f $X=-0.19 $Y=1.305 $X2=0.547 $Y2=0.995
cc_59 VPB N_A_216_93#_c_165_n 0.00417897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_216_93#_c_168_n 0.0105233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_410#_c_233_n 0.0265239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_410#_c_234_n 0.0263498f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_63 VPB N_A_27_410#_c_239_n 0.0164639f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_64 VPB N_A_27_410#_c_240_n 0.0216326f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.19
cc_65 VPB N_A_27_410#_c_241_n 0.00680513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_410#_c_242_n 0.00589342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_410#_c_243_n 0.00201281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_410#_c_235_n 9.16142e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_410#_c_245_n 0.0111036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_B_c_329_n 0.00604293f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.975
cc_71 VPB N_B_c_330_n 0.0511655f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_72 VPB N_B_M1009_g 0.0107583f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.995
cc_73 VPB B 0.0130977f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_c_369_n 0.0281529f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_75 VPB N_A_c_371_n 0.00333961f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_336_413#_c_417_n 0.0187074f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.445
cc_77 VPB N_A_336_413#_c_418_n 0.019582f $X=-0.19 $Y=1.305 $X2=0.547 $Y2=0.995
cc_78 VPB N_A_336_413#_c_419_n 0.00985638f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.53
cc_79 VPB N_A_336_413#_c_420_n 0.00256019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_336_413#_c_421_n 0.00407334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_336_413#_c_422_n 0.00156472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_336_413#_c_423_n 0.00139492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_336_413#_c_416_n 0.0272394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_538_n 0.0143673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_539_n 0.0113193f $X=-0.19 $Y=1.305 $X2=0.547 $Y2=0.995
cc_86 VPB N_VPWR_c_540_n 0.0131006f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_87 VPB N_VPWR_c_541_n 0.00940721f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.19
cc_88 VPB N_VPWR_c_542_n 0.0709048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_543_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_544_n 0.0145108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_545_n 0.0210157f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_546_n 0.00593769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_537_n 0.0747118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_X_c_603_n 0.00119494f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_95 N_C_N_c_98_n N_D_N_c_129_n 0.0105159f $X=0.547 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_96 N_C_N_c_99_n N_D_N_c_130_n 0.0219446f $X=0.495 $Y=1.875 $X2=0 $Y2=0
cc_97 N_C_N_c_100_n N_D_N_c_130_n 0.00196932f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_98 N_C_N_c_96_n N_D_N_c_130_n 0.0183318f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_99 N_C_N_c_97_n N_D_N_c_130_n 0.00929663f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_100 N_C_N_c_96_n D_N 2.91347e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_101 N_C_N_c_97_n D_N 0.0265431f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_102 N_C_N_c_97_n N_A_216_93#_c_171_n 0.0116733f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_103 N_C_N_c_96_n N_A_27_410#_c_234_n 0.0216334f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_104 N_C_N_c_97_n N_A_27_410#_c_234_n 0.0534696f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_105 N_C_N_c_98_n N_A_27_410#_c_234_n 0.00501087f $X=0.547 $Y=0.995 $X2=0
+ $Y2=0
cc_106 N_C_N_c_100_n N_A_27_410#_c_239_n 0.00559296f $X=0.495 $Y=1.975 $X2=0
+ $Y2=0
cc_107 N_C_N_c_99_n N_A_27_410#_c_240_n 0.00425397f $X=0.495 $Y=1.875 $X2=0
+ $Y2=0
cc_108 N_C_N_c_100_n N_A_27_410#_c_240_n 0.0121812f $X=0.495 $Y=1.975 $X2=0
+ $Y2=0
cc_109 N_C_N_c_96_n N_A_27_410#_c_240_n 3.38113e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_110 N_C_N_c_97_n N_A_27_410#_c_240_n 0.0318398f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_111 N_C_N_c_96_n N_A_27_410#_c_236_n 4.49664e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_112 N_C_N_c_98_n N_A_27_410#_c_236_n 0.00218147f $X=0.547 $Y=0.995 $X2=0
+ $Y2=0
cc_113 N_C_N_c_97_n N_VPWR_M1010_d 0.00436687f $X=0.53 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_114 N_C_N_c_100_n N_VPWR_c_538_n 0.0127593f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_115 N_C_N_c_100_n N_VPWR_c_544_n 0.00310301f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_116 N_C_N_c_100_n N_VPWR_c_537_n 0.00460685f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_117 N_C_N_c_97_n N_VGND_c_629_n 0.0108718f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_118 N_C_N_c_98_n N_VGND_c_629_n 0.00447091f $X=0.547 $Y=0.995 $X2=0 $Y2=0
cc_119 N_C_N_c_98_n N_VGND_c_635_n 0.00510437f $X=0.547 $Y=0.995 $X2=0 $Y2=0
cc_120 N_C_N_c_98_n N_VGND_c_643_n 0.00512902f $X=0.547 $Y=0.995 $X2=0 $Y2=0
cc_121 N_D_N_c_130_n N_A_216_93#_c_171_n 0.00834248f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_122 D_N N_A_216_93#_c_171_n 0.0173366f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_123 N_D_N_c_129_n N_A_216_93#_c_164_n 0.00406983f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_D_N_c_130_n N_A_216_93#_c_164_n 2.39076e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_125 D_N N_A_216_93#_c_164_n 0.00635704f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_126 N_D_N_c_130_n N_A_216_93#_c_165_n 0.00531552f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_127 D_N N_A_216_93#_c_165_n 0.00635704f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_128 N_D_N_c_129_n N_A_216_93#_c_166_n 0.00206399f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_129 N_D_N_c_130_n N_A_216_93#_c_166_n 0.00274492f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_130 D_N N_A_216_93#_c_166_n 0.0127706f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_131 N_D_N_c_130_n N_A_216_93#_c_167_n 5.83016e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_132 D_N N_A_216_93#_c_167_n 0.0144726f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_133 N_D_N_c_130_n N_A_216_93#_c_168_n 0.0119111f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_134 D_N N_A_216_93#_c_168_n 8.87853e-19 $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_135 N_D_N_c_130_n N_A_27_410#_c_240_n 0.0167468f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_136 D_N N_A_27_410#_c_240_n 0.00124584f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_137 N_D_N_c_130_n N_VPWR_c_542_n 0.0031102f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_138 N_D_N_c_130_n N_VPWR_c_537_n 0.00500987f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_139 N_D_N_c_129_n N_VGND_c_629_n 0.00291681f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_140 N_D_N_c_129_n N_VGND_c_630_n 0.00510437f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_141 N_D_N_c_129_n N_VGND_c_631_n 0.0030892f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_142 N_D_N_c_129_n N_VGND_c_643_n 0.00512902f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_216_93#_M1002_g N_A_27_410#_M1015_g 0.0246037f $X=2.065 $Y=0.445
+ $X2=0 $Y2=0
cc_144 N_A_216_93#_c_169_n N_A_27_410#_c_233_n 0.0229713f $X=2.04 $Y=1.89 $X2=0
+ $Y2=0
cc_145 N_A_216_93#_c_170_n N_A_27_410#_c_233_n 0.00116326f $X=2.04 $Y=1.99 $X2=0
+ $Y2=0
cc_146 N_A_216_93#_c_164_n N_A_27_410#_c_233_n 2.4865e-19 $X=1.605 $Y=1.075
+ $X2=0 $Y2=0
cc_147 N_A_216_93#_c_165_n N_A_27_410#_c_233_n 2.4865e-19 $X=1.605 $Y=1.525
+ $X2=0 $Y2=0
cc_148 N_A_216_93#_c_167_n N_A_27_410#_c_233_n 4.52975e-19 $X=1.77 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_216_93#_c_168_n N_A_27_410#_c_233_n 0.0219919f $X=2.065 $Y=1.16 $X2=0
+ $Y2=0
cc_150 N_A_216_93#_M1011_d N_A_27_410#_c_240_n 0.00258871f $X=1.12 $Y=1.485
+ $X2=0 $Y2=0
cc_151 N_A_216_93#_c_169_n N_A_27_410#_c_240_n 0.00101201f $X=2.04 $Y=1.89 $X2=0
+ $Y2=0
cc_152 N_A_216_93#_c_170_n N_A_27_410#_c_240_n 0.00744737f $X=2.04 $Y=1.99 $X2=0
+ $Y2=0
cc_153 N_A_216_93#_c_171_n N_A_27_410#_c_240_n 0.0449386f $X=1.51 $Y=1.61 $X2=0
+ $Y2=0
cc_154 N_A_216_93#_c_167_n N_A_27_410#_c_240_n 0.0045774f $X=1.77 $Y=1.16 $X2=0
+ $Y2=0
cc_155 N_A_216_93#_c_168_n N_A_27_410#_c_240_n 0.00315934f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_156 N_A_216_93#_c_169_n N_A_27_410#_c_241_n 0.0105998f $X=2.04 $Y=1.89 $X2=0
+ $Y2=0
cc_157 N_A_216_93#_c_171_n N_A_27_410#_c_241_n 0.00922297f $X=1.51 $Y=1.61 $X2=0
+ $Y2=0
cc_158 N_A_216_93#_c_169_n N_A_27_410#_c_242_n 0.0109553f $X=2.04 $Y=1.89 $X2=0
+ $Y2=0
cc_159 N_A_216_93#_c_169_n N_A_27_410#_c_243_n 0.00869215f $X=2.04 $Y=1.89 $X2=0
+ $Y2=0
cc_160 N_A_216_93#_c_171_n N_A_27_410#_c_243_n 0.0056179f $X=1.51 $Y=1.61 $X2=0
+ $Y2=0
cc_161 N_A_216_93#_c_165_n N_A_27_410#_c_243_n 0.00934447f $X=1.605 $Y=1.525
+ $X2=0 $Y2=0
cc_162 N_A_216_93#_c_167_n N_A_27_410#_c_243_n 0.00673601f $X=1.77 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_A_216_93#_c_168_n N_A_27_410#_c_243_n 0.00178889f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_164 N_A_216_93#_c_169_n N_A_27_410#_c_235_n 0.00171119f $X=2.04 $Y=1.89 $X2=0
+ $Y2=0
cc_165 N_A_216_93#_c_167_n N_A_27_410#_c_235_n 0.0056506f $X=1.77 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_A_216_93#_c_168_n N_A_27_410#_c_235_n 0.00173295f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_167 N_A_216_93#_c_170_n B 0.00308444f $X=2.04 $Y=1.99 $X2=0 $Y2=0
cc_168 N_A_216_93#_c_170_n N_A_336_413#_c_419_n 0.0121727f $X=2.04 $Y=1.99 $X2=0
+ $Y2=0
cc_169 N_A_216_93#_c_170_n N_A_336_413#_c_420_n 0.00679125f $X=2.04 $Y=1.99
+ $X2=0 $Y2=0
cc_170 N_A_216_93#_M1002_g N_A_336_413#_c_411_n 0.00249682f $X=2.065 $Y=0.445
+ $X2=0 $Y2=0
cc_171 N_A_216_93#_c_166_n N_A_336_413#_c_411_n 0.00739331f $X=1.265 $Y=0.66
+ $X2=0 $Y2=0
cc_172 N_A_216_93#_c_169_n N_A_336_413#_c_429_n 0.00151483f $X=2.04 $Y=1.89
+ $X2=0 $Y2=0
cc_173 N_A_216_93#_c_170_n N_VPWR_c_542_n 0.00451183f $X=2.04 $Y=1.99 $X2=0
+ $Y2=0
cc_174 N_A_216_93#_c_170_n N_VPWR_c_537_n 0.00874597f $X=2.04 $Y=1.99 $X2=0
+ $Y2=0
cc_175 N_A_216_93#_c_166_n N_VGND_M1002_s 4.10598e-19 $X=1.265 $Y=0.66 $X2=0
+ $Y2=0
cc_176 N_A_216_93#_c_166_n N_VGND_c_629_n 0.0101148f $X=1.265 $Y=0.66 $X2=0
+ $Y2=0
cc_177 N_A_216_93#_c_166_n N_VGND_c_630_n 0.0095527f $X=1.265 $Y=0.66 $X2=0
+ $Y2=0
cc_178 N_A_216_93#_M1002_g N_VGND_c_631_n 0.00831102f $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_A_216_93#_c_166_n N_VGND_c_631_n 0.0108829f $X=1.265 $Y=0.66 $X2=0
+ $Y2=0
cc_180 N_A_216_93#_c_167_n N_VGND_c_631_n 0.00711768f $X=1.77 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_A_216_93#_c_168_n N_VGND_c_631_n 0.00525518f $X=2.065 $Y=1.16 $X2=0
+ $Y2=0
cc_182 N_A_216_93#_M1002_g N_VGND_c_632_n 6.93631e-19 $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_183 N_A_216_93#_M1002_g N_VGND_c_637_n 0.00585385f $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_184 N_A_216_93#_M1002_g N_VGND_c_643_n 0.0121761f $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_185 N_A_216_93#_c_166_n N_VGND_c_643_n 0.0131649f $X=1.265 $Y=0.66 $X2=0
+ $Y2=0
cc_186 N_A_27_410#_M1015_g N_B_c_326_n 0.0128519f $X=2.55 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_187 N_A_27_410#_c_233_n N_B_c_327_n 0.0259242f $X=2.57 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_27_410#_c_235_n N_B_c_327_n 3.37553e-19 $X=2.485 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_27_410#_c_235_n N_B_c_329_n 4.70706e-19 $X=2.485 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_27_410#_c_233_n N_B_M1009_g 0.0359634f $X=2.57 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A_27_410#_c_242_n N_B_M1009_g 7.32223e-19 $X=2.4 $Y=1.5 $X2=0 $Y2=0
cc_192 N_A_27_410#_M1015_g N_B_c_328_n 0.012133f $X=2.55 $Y=0.445 $X2=0 $Y2=0
cc_193 N_A_27_410#_c_233_n N_A_c_371_n 0.00252948f $X=2.57 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_27_410#_c_235_n N_A_c_371_n 0.0187646f $X=2.485 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_27_410#_c_240_n N_A_336_413#_c_419_n 0.0273036f $X=1.87 $Y=1.95 $X2=0
+ $Y2=0
cc_196 N_A_27_410#_c_242_n N_A_336_413#_c_419_n 0.0049489f $X=2.4 $Y=1.5 $X2=0
+ $Y2=0
cc_197 N_A_27_410#_M1015_g N_A_336_413#_c_432_n 0.00511329f $X=2.55 $Y=0.445
+ $X2=0 $Y2=0
cc_198 N_A_27_410#_c_233_n N_A_336_413#_c_420_n 0.00198717f $X=2.57 $Y=1.41
+ $X2=0 $Y2=0
cc_199 N_A_27_410#_c_240_n N_A_336_413#_c_420_n 0.00508372f $X=1.87 $Y=1.95
+ $X2=0 $Y2=0
cc_200 N_A_27_410#_M1015_g N_A_336_413#_c_410_n 0.0127455f $X=2.55 $Y=0.445
+ $X2=0 $Y2=0
cc_201 N_A_27_410#_c_233_n N_A_336_413#_c_410_n 0.00345912f $X=2.57 $Y=1.41
+ $X2=0 $Y2=0
cc_202 N_A_27_410#_c_242_n N_A_336_413#_c_410_n 0.0012205f $X=2.4 $Y=1.5 $X2=0
+ $Y2=0
cc_203 N_A_27_410#_c_235_n N_A_336_413#_c_410_n 0.012923f $X=2.485 $Y=1.16 $X2=0
+ $Y2=0
cc_204 N_A_27_410#_c_233_n N_A_336_413#_c_411_n 2.86694e-19 $X=2.57 $Y=1.41
+ $X2=0 $Y2=0
cc_205 N_A_27_410#_c_242_n N_A_336_413#_c_411_n 0.00589573f $X=2.4 $Y=1.5 $X2=0
+ $Y2=0
cc_206 N_A_27_410#_c_233_n N_A_336_413#_c_421_n 0.0149855f $X=2.57 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_27_410#_c_242_n N_A_336_413#_c_421_n 0.00590782f $X=2.4 $Y=1.5 $X2=0
+ $Y2=0
cc_208 N_A_27_410#_c_233_n N_A_336_413#_c_429_n 2.30045e-19 $X=2.57 $Y=1.41
+ $X2=0 $Y2=0
cc_209 N_A_27_410#_c_240_n N_A_336_413#_c_429_n 0.00640417f $X=1.87 $Y=1.95
+ $X2=0 $Y2=0
cc_210 N_A_27_410#_c_241_n N_A_336_413#_c_429_n 0.0051505f $X=1.955 $Y=1.865
+ $X2=0 $Y2=0
cc_211 N_A_27_410#_c_242_n N_A_336_413#_c_429_n 0.0117409f $X=2.4 $Y=1.5 $X2=0
+ $Y2=0
cc_212 N_A_27_410#_c_242_n N_A_336_413#_c_423_n 0.00240533f $X=2.4 $Y=1.5 $X2=0
+ $Y2=0
cc_213 N_A_27_410#_c_240_n N_VPWR_M1010_d 0.00562672f $X=1.87 $Y=1.95 $X2=-0.19
+ $Y2=-0.24
cc_214 N_A_27_410#_c_239_n N_VPWR_c_538_n 0.0192602f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_215 N_A_27_410#_c_240_n N_VPWR_c_538_n 0.0265965f $X=1.87 $Y=1.95 $X2=0 $Y2=0
cc_216 N_A_27_410#_c_233_n N_VPWR_c_542_n 0.00393512f $X=2.57 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A_27_410#_c_240_n N_VPWR_c_542_n 0.0118526f $X=1.87 $Y=1.95 $X2=0 $Y2=0
cc_218 N_A_27_410#_c_239_n N_VPWR_c_544_n 0.017058f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_219 N_A_27_410#_c_240_n N_VPWR_c_544_n 0.00257955f $X=1.87 $Y=1.95 $X2=0
+ $Y2=0
cc_220 N_A_27_410#_c_233_n N_VPWR_c_537_n 0.00500987f $X=2.57 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_27_410#_c_239_n N_VPWR_c_537_n 0.00987673f $X=0.26 $Y=2.29 $X2=0
+ $Y2=0
cc_222 N_A_27_410#_c_240_n N_VPWR_c_537_n 0.0260532f $X=1.87 $Y=1.95 $X2=0 $Y2=0
cc_223 N_A_27_410#_c_242_n A_426_413# 0.00275594f $X=2.4 $Y=1.5 $X2=-0.19
+ $Y2=-0.24
cc_224 N_A_27_410#_c_236_n N_VGND_c_629_n 0.018587f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_225 N_A_27_410#_M1015_g N_VGND_c_632_n 0.0103553f $X=2.55 $Y=0.445 $X2=0
+ $Y2=0
cc_226 N_A_27_410#_c_236_n N_VGND_c_635_n 0.00972557f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_227 N_A_27_410#_M1015_g N_VGND_c_637_n 0.00199015f $X=2.55 $Y=0.445 $X2=0
+ $Y2=0
cc_228 N_A_27_410#_M1015_g N_VGND_c_643_n 0.00284206f $X=2.55 $Y=0.445 $X2=0
+ $Y2=0
cc_229 N_A_27_410#_c_236_n N_VGND_c_643_n 0.0107261f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_230 N_B_c_327_n N_A_c_369_n 0.0213315f $X=2.98 $Y=1.31 $X2=-0.19 $Y2=-0.24
cc_231 N_B_c_329_n N_A_c_369_n 0.00417671f $X=2.98 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_232 N_B_M1009_g N_A_c_369_n 0.0247568f $X=2.98 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_233 B N_A_c_369_n 6.06139e-19 $X=3.18 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_234 N_B_c_328_n N_A_M1007_g 0.0196004f $X=2.98 $Y=0.76 $X2=0 $Y2=0
cc_235 N_B_c_327_n N_A_c_371_n 0.0122623f $X=2.98 $Y=1.31 $X2=0 $Y2=0
cc_236 N_B_c_329_n N_A_c_371_n 0.00510764f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B_c_330_n N_A_336_413#_c_419_n 9.02506e-19 $X=2.98 $Y=2.035 $X2=0 $Y2=0
cc_238 B N_A_336_413#_c_419_n 0.0113771f $X=3.18 $Y=2.125 $X2=0 $Y2=0
cc_239 N_B_c_330_n N_A_336_413#_c_420_n 0.00275425f $X=2.98 $Y=2.035 $X2=0 $Y2=0
cc_240 B N_A_336_413#_c_420_n 0.00474738f $X=3.18 $Y=2.125 $X2=0 $Y2=0
cc_241 N_B_c_326_n N_A_336_413#_c_410_n 0.00630115f $X=2.98 $Y=0.86 $X2=0 $Y2=0
cc_242 N_B_c_328_n N_A_336_413#_c_410_n 0.00765134f $X=2.98 $Y=0.76 $X2=0 $Y2=0
cc_243 N_B_c_330_n N_A_336_413#_c_421_n 0.00109209f $X=2.98 $Y=2.035 $X2=0 $Y2=0
cc_244 N_B_M1009_g N_A_336_413#_c_421_n 0.0125693f $X=2.98 $Y=1.695 $X2=0 $Y2=0
cc_245 B N_A_336_413#_c_421_n 0.0385061f $X=3.18 $Y=2.125 $X2=0 $Y2=0
cc_246 N_B_M1009_g N_A_336_413#_c_423_n 0.00550607f $X=2.98 $Y=1.695 $X2=0 $Y2=0
cc_247 B N_A_336_413#_c_423_n 0.0138656f $X=3.18 $Y=2.125 $X2=0 $Y2=0
cc_248 N_B_c_330_n N_VPWR_c_539_n 0.00373437f $X=2.98 $Y=2.035 $X2=0 $Y2=0
cc_249 B N_VPWR_c_539_n 0.0239479f $X=3.18 $Y=2.125 $X2=0 $Y2=0
cc_250 N_B_c_330_n N_VPWR_c_542_n 0.00836618f $X=2.98 $Y=2.035 $X2=0 $Y2=0
cc_251 B N_VPWR_c_542_n 0.0427446f $X=3.18 $Y=2.125 $X2=0 $Y2=0
cc_252 N_B_c_330_n N_VPWR_c_537_n 0.011783f $X=2.98 $Y=2.035 $X2=0 $Y2=0
cc_253 B N_VPWR_c_537_n 0.0257296f $X=3.18 $Y=2.125 $X2=0 $Y2=0
cc_254 N_B_c_328_n N_VGND_c_632_n 0.00167196f $X=2.98 $Y=0.76 $X2=0 $Y2=0
cc_255 N_B_c_328_n N_VGND_c_639_n 6.85223e-19 $X=2.98 $Y=0.76 $X2=0 $Y2=0
cc_256 N_B_c_328_n N_VGND_c_640_n 0.00428022f $X=2.98 $Y=0.76 $X2=0 $Y2=0
cc_257 N_B_c_328_n N_VGND_c_643_n 0.00594333f $X=2.98 $Y=0.76 $X2=0 $Y2=0
cc_258 N_A_c_369_n N_A_336_413#_c_417_n 0.0154284f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_M1007_g N_A_336_413#_c_408_n 0.0180813f $X=3.49 $Y=0.445 $X2=0 $Y2=0
cc_260 N_A_c_371_n N_A_336_413#_c_410_n 0.0225698f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_c_371_n N_A_336_413#_c_421_n 0.0116453f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A_c_369_n N_A_336_413#_c_412_n 0.0034911f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_M1007_g N_A_336_413#_c_412_n 0.011693f $X=3.49 $Y=0.445 $X2=0 $Y2=0
cc_264 N_A_c_371_n N_A_336_413#_c_412_n 0.0204446f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_c_369_n N_A_336_413#_c_466_n 0.0141289f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A_c_371_n N_A_336_413#_c_466_n 0.0129269f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A_c_369_n N_A_336_413#_c_422_n 0.00348305f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_c_369_n N_A_336_413#_c_413_n 5.77159e-19 $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A_c_371_n N_A_336_413#_c_413_n 0.0146254f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_c_369_n N_A_336_413#_c_423_n 0.0110462f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A_c_371_n N_A_336_413#_c_423_n 0.0112473f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_c_369_n N_A_336_413#_c_414_n 0.00190284f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A_c_371_n N_A_336_413#_c_414_n 0.0271506f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_M1007_g N_A_336_413#_c_415_n 0.00353282f $X=3.49 $Y=0.445 $X2=0 $Y2=0
cc_275 N_A_c_369_n N_A_336_413#_c_416_n 0.0233474f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A_c_371_n N_A_336_413#_c_416_n 3.51189e-19 $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_c_369_n N_VPWR_c_539_n 0.00330158f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_c_369_n N_VPWR_c_542_n 0.00351015f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A_c_369_n N_VPWR_c_537_n 0.00445321f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A_M1007_g N_VGND_c_639_n 0.0105644f $X=3.49 $Y=0.445 $X2=0 $Y2=0
cc_281 N_A_M1007_g N_VGND_c_640_n 0.00199743f $X=3.49 $Y=0.445 $X2=0 $Y2=0
cc_282 N_A_M1007_g N_VGND_c_643_n 0.00284206f $X=3.49 $Y=0.445 $X2=0 $Y2=0
cc_283 N_A_336_413#_c_466_n N_VPWR_M1000_d 0.00563715f $X=3.765 $Y=1.58 $X2=0
+ $Y2=0
cc_284 N_A_336_413#_c_417_n N_VPWR_c_539_n 0.00482583f $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_285 N_A_336_413#_c_466_n N_VPWR_c_539_n 0.0204259f $X=3.765 $Y=1.58 $X2=0
+ $Y2=0
cc_286 N_A_336_413#_c_423_n N_VPWR_c_539_n 0.00726621f $X=3.31 $Y=1.58 $X2=0
+ $Y2=0
cc_287 N_A_336_413#_c_416_n N_VPWR_c_539_n 2.27534e-19 $X=4.475 $Y=1.202 $X2=0
+ $Y2=0
cc_288 N_A_336_413#_c_418_n N_VPWR_c_541_n 0.00840319f $X=4.475 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_336_413#_c_419_n N_VPWR_c_542_n 0.0304719f $X=2.26 $Y=2.29 $X2=0
+ $Y2=0
cc_290 N_A_336_413#_c_417_n N_VPWR_c_545_n 0.00702461f $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_291 N_A_336_413#_c_418_n N_VPWR_c_545_n 0.00597712f $X=4.475 $Y=1.41 $X2=0
+ $Y2=0
cc_292 N_A_336_413#_M1008_s N_VPWR_c_537_n 0.002265f $X=1.68 $Y=2.065 $X2=0
+ $Y2=0
cc_293 N_A_336_413#_c_417_n N_VPWR_c_537_n 0.0137694f $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_294 N_A_336_413#_c_418_n N_VPWR_c_537_n 0.0110832f $X=4.475 $Y=1.41 $X2=0
+ $Y2=0
cc_295 N_A_336_413#_c_419_n N_VPWR_c_537_n 0.027257f $X=2.26 $Y=2.29 $X2=0 $Y2=0
cc_296 N_A_336_413#_c_421_n N_VPWR_c_537_n 0.0102114f $X=3.225 $Y=1.87 $X2=0
+ $Y2=0
cc_297 N_A_336_413#_c_419_n A_426_413# 0.0046523f $X=2.26 $Y=2.29 $X2=-0.19
+ $Y2=-0.24
cc_298 N_A_336_413#_c_420_n A_426_413# 0.00311349f $X=2.345 $Y=2.205 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_336_413#_c_429_n A_426_413# 0.00379949f $X=2.43 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_300 N_A_336_413#_c_421_n A_532_297# 0.00442604f $X=3.225 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_301 N_A_336_413#_c_421_n A_614_297# 0.00197899f $X=3.225 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_302 N_A_336_413#_c_423_n A_614_297# 0.00482155f $X=3.31 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_303 N_A_336_413#_c_409_n N_X_c_605_n 0.00454228f $X=4.5 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A_336_413#_c_416_n N_X_c_605_n 0.00279746f $X=4.475 $Y=1.202 $X2=0
+ $Y2=0
cc_305 N_A_336_413#_c_417_n N_X_c_607_n 0.00842225f $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A_336_413#_c_418_n N_X_c_607_n 0.00369418f $X=4.475 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A_336_413#_c_466_n N_X_c_607_n 0.0111625f $X=3.765 $Y=1.58 $X2=0 $Y2=0
cc_308 N_A_336_413#_c_416_n N_X_c_607_n 0.00477572f $X=4.475 $Y=1.202 $X2=0
+ $Y2=0
cc_309 N_A_336_413#_c_417_n N_X_c_603_n 6.48952e-19 $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A_336_413#_c_408_n N_X_c_603_n 0.00179029f $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A_336_413#_c_418_n N_X_c_603_n 0.00270904f $X=4.475 $Y=1.41 $X2=0 $Y2=0
cc_312 N_A_336_413#_c_409_n N_X_c_603_n 0.00706836f $X=4.5 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A_336_413#_c_422_n N_X_c_603_n 0.00749371f $X=3.85 $Y=1.495 $X2=0 $Y2=0
cc_314 N_A_336_413#_c_414_n N_X_c_603_n 0.0190929f $X=3.955 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A_336_413#_c_415_n N_X_c_603_n 0.00666144f $X=3.902 $Y=0.995 $X2=0
+ $Y2=0
cc_316 N_A_336_413#_c_416_n N_X_c_603_n 0.0333631f $X=4.475 $Y=1.202 $X2=0 $Y2=0
cc_317 N_A_336_413#_c_418_n X 0.0138037f $X=4.475 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_336_413#_c_412_n N_VGND_M1007_d 0.00652347f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_319 N_A_336_413#_c_415_n N_VGND_M1007_d 6.98847e-19 $X=3.902 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_A_336_413#_c_432_n N_VGND_c_632_n 0.0125877f $X=2.275 $Y=0.47 $X2=0
+ $Y2=0
cc_321 N_A_336_413#_c_410_n N_VGND_c_632_n 0.0242276f $X=3.145 $Y=0.74 $X2=0
+ $Y2=0
cc_322 N_A_336_413#_c_409_n N_VGND_c_634_n 0.00971011f $X=4.5 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_336_413#_c_432_n N_VGND_c_637_n 0.00861358f $X=2.275 $Y=0.47 $X2=0
+ $Y2=0
cc_324 N_A_336_413#_c_410_n N_VGND_c_637_n 0.00309172f $X=3.145 $Y=0.74 $X2=0
+ $Y2=0
cc_325 N_A_336_413#_c_408_n N_VGND_c_639_n 0.00463088f $X=4.03 $Y=0.995 $X2=0
+ $Y2=0
cc_326 N_A_336_413#_c_521_p N_VGND_c_639_n 0.0135697f $X=3.23 $Y=0.47 $X2=0
+ $Y2=0
cc_327 N_A_336_413#_c_412_n N_VGND_c_639_n 0.0298327f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_328 N_A_336_413#_c_416_n N_VGND_c_639_n 3.3049e-19 $X=4.475 $Y=1.202 $X2=0
+ $Y2=0
cc_329 N_A_336_413#_c_410_n N_VGND_c_640_n 0.0035533f $X=3.145 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_A_336_413#_c_521_p N_VGND_c_640_n 0.00876148f $X=3.23 $Y=0.47 $X2=0
+ $Y2=0
cc_331 N_A_336_413#_c_412_n N_VGND_c_640_n 0.00283814f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_332 N_A_336_413#_c_408_n N_VGND_c_641_n 0.00585385f $X=4.03 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_A_336_413#_c_409_n N_VGND_c_641_n 0.00546121f $X=4.5 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_336_413#_M1002_d N_VGND_c_643_n 0.00494728f $X=2.14 $Y=0.235 $X2=0
+ $Y2=0
cc_335 N_A_336_413#_M1012_d N_VGND_c_643_n 0.00336566f $X=3.08 $Y=0.235 $X2=0
+ $Y2=0
cc_336 N_A_336_413#_c_408_n N_VGND_c_643_n 0.0111006f $X=4.03 $Y=0.995 $X2=0
+ $Y2=0
cc_337 N_A_336_413#_c_409_n N_VGND_c_643_n 0.010748f $X=4.5 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A_336_413#_c_432_n N_VGND_c_643_n 0.00625722f $X=2.275 $Y=0.47 $X2=0
+ $Y2=0
cc_339 N_A_336_413#_c_410_n N_VGND_c_643_n 0.0117669f $X=3.145 $Y=0.74 $X2=0
+ $Y2=0
cc_340 N_A_336_413#_c_521_p N_VGND_c_643_n 0.00625722f $X=3.23 $Y=0.47 $X2=0
+ $Y2=0
cc_341 N_A_336_413#_c_412_n N_VGND_c_643_n 0.00690419f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_537_n A_426_413# 0.00222986f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_343 N_VPWR_c_537_n N_X_M1004_s 0.00444633f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_344 N_VPWR_c_541_n N_X_c_603_n 0.0674594f $X=4.735 $Y=1.66 $X2=0 $Y2=0
cc_345 N_VPWR_c_545_n X 0.018822f $X=4.65 $Y=2.72 $X2=0 $Y2=0
cc_346 N_VPWR_c_537_n X 0.011161f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_347 N_VPWR_c_541_n N_VGND_c_634_n 0.00716889f $X=4.735 $Y=1.66 $X2=0 $Y2=0
cc_348 N_X_c_605_n N_VGND_c_634_n 0.0227154f $X=4.357 $Y=0.587 $X2=0 $Y2=0
cc_349 N_X_c_603_n N_VGND_c_634_n 0.00993153f $X=4.305 $Y=1.495 $X2=0 $Y2=0
cc_350 N_X_c_605_n N_VGND_c_641_n 0.00881626f $X=4.357 $Y=0.587 $X2=0 $Y2=0
cc_351 N_X_M1013_s N_VGND_c_643_n 0.00454589f $X=4.105 $Y=0.235 $X2=0 $Y2=0
cc_352 N_X_c_605_n N_VGND_c_643_n 0.0101156f $X=4.357 $Y=0.587 $X2=0 $Y2=0
