* File: sky130_fd_sc_hdll__ebufn_1.pxi.spice
* Created: Wed Sep  2 08:30:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__EBUFN_1%A N_A_c_63_n N_A_c_64_n N_A_M1001_g N_A_M1005_g
+ A A N_A_c_62_n PM_SKY130_FD_SC_HDLL__EBUFN_1%A
x_PM_SKY130_FD_SC_HDLL__EBUFN_1%TE_B N_TE_B_c_91_n N_TE_B_c_92_n N_TE_B_M1007_g
+ N_TE_B_c_88_n N_TE_B_M1006_g N_TE_B_c_93_n N_TE_B_M1003_g N_TE_B_c_89_n
+ N_TE_B_c_90_n TE_B TE_B PM_SKY130_FD_SC_HDLL__EBUFN_1%TE_B
x_PM_SKY130_FD_SC_HDLL__EBUFN_1%A_211_369# N_A_211_369#_M1006_d
+ N_A_211_369#_M1007_d N_A_211_369#_M1002_g N_A_211_369#_c_143_n
+ N_A_211_369#_c_139_n N_A_211_369#_c_144_n N_A_211_369#_c_140_n
+ N_A_211_369#_c_141_n N_A_211_369#_c_158_n N_A_211_369#_c_142_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_1%A_211_369#
x_PM_SKY130_FD_SC_HDLL__EBUFN_1%A_27_47# N_A_27_47#_M1005_s N_A_27_47#_M1001_s
+ N_A_27_47#_c_194_n N_A_27_47#_M1000_g N_A_27_47#_c_195_n N_A_27_47#_M1004_g
+ N_A_27_47#_c_196_n N_A_27_47#_c_206_n N_A_27_47#_c_197_n N_A_27_47#_c_223_n
+ N_A_27_47#_c_198_n N_A_27_47#_c_218_n N_A_27_47#_c_199_n N_A_27_47#_c_200_n
+ N_A_27_47#_c_201_n N_A_27_47#_c_202_n N_A_27_47#_c_203_n N_A_27_47#_c_204_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EBUFN_1%VPWR N_VPWR_M1001_d N_VPWR_M1003_s
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n VPWR N_VPWR_c_302_n
+ N_VPWR_c_303_n N_VPWR_c_298_n N_VPWR_c_305_n N_VPWR_c_306_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_1%VPWR
x_PM_SKY130_FD_SC_HDLL__EBUFN_1%Z N_Z_M1000_d N_Z_M1004_d Z Z Z Z Z Z Z
+ N_Z_c_350_n Z Z N_Z_c_346_n N_Z_c_348_n Z PM_SKY130_FD_SC_HDLL__EBUFN_1%Z
x_PM_SKY130_FD_SC_HDLL__EBUFN_1%VGND N_VGND_M1005_d N_VGND_M1002_s VGND
+ N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n
+ N_VGND_c_377_n PM_SKY130_FD_SC_HDLL__EBUFN_1%VGND
cc_1 VNB N_A_M1005_g 0.0379393f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A 0.0137853f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_c_62_n 0.0365501f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_TE_B_c_88_n 0.0300213f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_5 VNB N_TE_B_c_89_n 0.0159446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_TE_B_c_90_n 0.0653334f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_7 VNB N_A_211_369#_c_139_n 0.00738655f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_8 VNB N_A_211_369#_c_140_n 0.00536902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_211_369#_c_141_n 0.0210764f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_211_369#_c_142_n 0.0194452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_194_n 0.0172583f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_12 VNB N_A_27_47#_c_195_n 0.0237459f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_13 VNB N_A_27_47#_c_196_n 0.0132408f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_14 VNB N_A_27_47#_c_197_n 0.00348705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_198_n 0.0126163f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.53
cc_16 VNB N_A_27_47#_c_199_n 0.0224262f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_200_n 9.80023e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_201_n 0.0116929f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_202_n 0.00877432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_203_n 0.00450322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_204_n 0.00646242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_298_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB Z 0.00638732f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_24 VNB N_Z_c_346_n 0.0159232f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB Z 0.0241221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_372_n 0.0143912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_373_n 0.0169978f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.53
cc_28 VNB N_VGND_c_374_n 0.211356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_375_n 0.010096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_376_n 0.0341517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_377_n 0.0141533f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_c_63_n 0.0206487f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_33 VPB N_A_c_64_n 0.0279218f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_34 VPB A 0.016491f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_35 VPB N_A_c_62_n 0.00928613f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_36 VPB N_TE_B_c_91_n 0.0234188f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_37 VPB N_TE_B_c_92_n 0.0267598f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_38 VPB N_TE_B_c_93_n 0.0235775f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_TE_B_c_89_n 0.00188402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_TE_B_c_90_n 0.0335121f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_41 VPB TE_B 0.00610531f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_42 VPB N_A_211_369#_c_143_n 0.0055341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_211_369#_c_144_n 0.0152926f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_44 VPB N_A_211_369#_c_140_n 0.00552913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_211_369#_c_141_n 0.00791441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_195_n 0.0354728f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_47 VPB N_A_27_47#_c_206_n 0.0179778f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_48 VPB N_A_27_47#_c_197_n 0.0174098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_204_n 3.95116e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_299_n 4.18643e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_300_n 0.0165601f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_52 VPB N_VPWR_c_301_n 0.0058948f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_53 VPB N_VPWR_c_302_n 0.0194426f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_54 VPB N_VPWR_c_303_n 0.0438085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_298_n 0.0407245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_305_n 0.00496502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_306_n 0.00568265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_Z_c_348_n 0.0427352f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB Z 0.0103884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 N_A_c_63_n N_TE_B_c_91_n 0.011537f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_61 N_A_c_64_n N_TE_B_c_92_n 0.0329538f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_62 N_A_M1005_g N_TE_B_c_88_n 0.0195787f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_63 N_A_c_62_n N_TE_B_c_89_n 0.011537f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_c_62_n TE_B 4.42273e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_c_64_n N_A_27_47#_c_206_n 0.00593439f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_66 N_A_c_63_n N_A_27_47#_c_197_n 0.00970026f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_67 N_A_c_64_n N_A_27_47#_c_197_n 0.0267322f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_68 N_A_M1005_g N_A_27_47#_c_197_n 0.00969787f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_69 A N_A_27_47#_c_197_n 0.0690382f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_c_62_n N_A_27_47#_c_197_n 0.0114532f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_M1005_g N_A_27_47#_c_198_n 0.0162248f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_72 A N_A_27_47#_c_198_n 0.0218104f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_73 N_A_c_62_n N_A_27_47#_c_198_n 0.005262f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_M1005_g N_A_27_47#_c_218_n 5.0541e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A_c_64_n N_VPWR_c_299_n 0.0121612f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_76 N_A_c_64_n N_VPWR_c_302_n 0.00319306f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_77 N_A_c_64_n N_VPWR_c_298_n 0.00484792f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_78 N_A_M1005_g N_VGND_c_372_n 0.00196986f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_79 N_A_M1005_g N_VGND_c_374_n 0.00364793f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_80 N_A_M1005_g N_VGND_c_375_n 0.0126022f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_81 N_TE_B_c_92_n N_A_211_369#_c_143_n 0.00604845f $X=0.965 $Y=1.77 $X2=0
+ $Y2=0
cc_82 N_TE_B_c_93_n N_A_211_369#_c_143_n 0.00340357f $X=1.965 $Y=1.41 $X2=0
+ $Y2=0
cc_83 N_TE_B_c_88_n N_A_211_369#_c_139_n 0.00435552f $X=1.025 $Y=0.995 $X2=0
+ $Y2=0
cc_84 N_TE_B_c_90_n N_A_211_369#_c_139_n 0.0130656f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_85 N_TE_B_c_91_n N_A_211_369#_c_144_n 0.00421158f $X=0.965 $Y=1.67 $X2=0
+ $Y2=0
cc_86 N_TE_B_c_92_n N_A_211_369#_c_144_n 0.00600204f $X=0.965 $Y=1.77 $X2=0
+ $Y2=0
cc_87 N_TE_B_c_93_n N_A_211_369#_c_144_n 0.0243908f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_88 N_TE_B_c_90_n N_A_211_369#_c_144_n 0.0123106f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_89 TE_B N_A_211_369#_c_144_n 0.0405817f $X=1.02 $Y=1.105 $X2=0 $Y2=0
cc_90 N_TE_B_c_90_n N_A_211_369#_c_140_n 0.0164793f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_91 N_TE_B_c_90_n N_A_211_369#_c_141_n 0.0108561f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_92 N_TE_B_c_90_n N_A_211_369#_c_158_n 0.0250914f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_93 TE_B N_A_211_369#_c_158_n 0.0199562f $X=1.02 $Y=1.105 $X2=0 $Y2=0
cc_94 N_TE_B_c_92_n N_A_27_47#_c_197_n 0.00242329f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_95 N_TE_B_c_88_n N_A_27_47#_c_197_n 0.00207429f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_96 N_TE_B_c_89_n N_A_27_47#_c_197_n 0.00740247f $X=0.982 $Y=1.16 $X2=0 $Y2=0
cc_97 TE_B N_A_27_47#_c_197_n 0.0431252f $X=1.02 $Y=1.105 $X2=0 $Y2=0
cc_98 N_TE_B_c_88_n N_A_27_47#_c_223_n 0.0147309f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_99 N_TE_B_c_89_n N_A_27_47#_c_223_n 0.00256391f $X=0.982 $Y=1.16 $X2=0 $Y2=0
cc_100 N_TE_B_c_90_n N_A_27_47#_c_223_n 0.00303294f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_101 TE_B N_A_27_47#_c_223_n 0.0144816f $X=1.02 $Y=1.105 $X2=0 $Y2=0
cc_102 N_TE_B_c_88_n N_A_27_47#_c_218_n 0.00532102f $X=1.025 $Y=0.995 $X2=0
+ $Y2=0
cc_103 N_TE_B_c_90_n N_A_27_47#_c_199_n 0.00982463f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_104 TE_B N_A_27_47#_c_199_n 0.00160979f $X=1.02 $Y=1.105 $X2=0 $Y2=0
cc_105 N_TE_B_c_88_n N_A_27_47#_c_200_n 0.00778901f $X=1.025 $Y=0.995 $X2=0
+ $Y2=0
cc_106 N_TE_B_c_90_n N_A_27_47#_c_203_n 0.00310791f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_107 N_TE_B_c_92_n N_VPWR_c_299_n 0.00835522f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_108 N_TE_B_c_92_n N_VPWR_c_300_n 0.00642146f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_109 N_TE_B_c_92_n N_VPWR_c_301_n 0.00220651f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_110 N_TE_B_c_93_n N_VPWR_c_301_n 0.0114532f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_111 N_TE_B_c_93_n N_VPWR_c_303_n 0.0059915f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_112 N_TE_B_c_92_n N_VPWR_c_298_n 0.0121178f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_113 N_TE_B_c_93_n N_VPWR_c_298_n 0.011314f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_114 N_TE_B_c_93_n N_Z_c_350_n 0.0274649f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_115 N_TE_B_c_88_n N_VGND_c_374_n 0.00510711f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_116 N_TE_B_c_88_n N_VGND_c_375_n 0.00307718f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_117 N_TE_B_c_88_n N_VGND_c_376_n 0.00341702f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_211_369#_c_142_n N_A_27_47#_c_194_n 0.0388406f $X=2.58 $Y=0.995 $X2=0
+ $Y2=0
cc_119 N_A_211_369#_c_140_n N_A_27_47#_c_195_n 9.14502e-19 $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_120 N_A_211_369#_c_141_n N_A_27_47#_c_195_n 0.0388406f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_121 N_A_211_369#_c_139_n N_A_27_47#_c_197_n 0.00724176f $X=1.625 $Y=0.76
+ $X2=0 $Y2=0
cc_122 N_A_211_369#_c_144_n N_A_27_47#_c_197_n 0.0169015f $X=1.682 $Y=1.8 $X2=0
+ $Y2=0
cc_123 N_A_211_369#_M1006_d N_A_27_47#_c_223_n 0.00407554f $X=1.1 $Y=0.465 $X2=0
+ $Y2=0
cc_124 N_A_211_369#_c_139_n N_A_27_47#_c_223_n 0.0131399f $X=1.625 $Y=0.76 $X2=0
+ $Y2=0
cc_125 N_A_211_369#_M1006_d N_A_27_47#_c_218_n 0.00564702f $X=1.1 $Y=0.465 $X2=0
+ $Y2=0
cc_126 N_A_211_369#_c_139_n N_A_27_47#_c_199_n 0.0260704f $X=1.625 $Y=0.76 $X2=0
+ $Y2=0
cc_127 N_A_211_369#_c_140_n N_A_27_47#_c_199_n 0.00153568f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_128 N_A_211_369#_c_158_n N_A_27_47#_c_199_n 0.00349872f $X=1.682 $Y=1.2 $X2=0
+ $Y2=0
cc_129 N_A_211_369#_c_139_n N_A_27_47#_c_201_n 0.0080263f $X=1.625 $Y=0.76 $X2=0
+ $Y2=0
cc_130 N_A_211_369#_c_142_n N_A_27_47#_c_201_n 0.00460598f $X=2.58 $Y=0.995
+ $X2=0 $Y2=0
cc_131 N_A_211_369#_c_140_n N_A_27_47#_c_202_n 0.0425416f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_211_369#_c_141_n N_A_27_47#_c_202_n 0.00295767f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_A_211_369#_c_142_n N_A_27_47#_c_202_n 0.0118868f $X=2.58 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_A_211_369#_c_139_n N_A_27_47#_c_203_n 0.0150385f $X=1.625 $Y=0.76 $X2=0
+ $Y2=0
cc_135 N_A_211_369#_c_140_n N_A_27_47#_c_203_n 0.0181628f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_211_369#_c_140_n N_A_27_47#_c_204_n 0.0214816f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_211_369#_c_141_n N_A_27_47#_c_204_n 7.09784e-19 $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_211_369#_c_142_n N_A_27_47#_c_204_n 0.00342037f $X=2.58 $Y=0.995
+ $X2=0 $Y2=0
cc_139 N_A_211_369#_c_144_n N_VPWR_M1003_s 0.00628911f $X=1.682 $Y=1.8 $X2=0
+ $Y2=0
cc_140 N_A_211_369#_c_143_n N_VPWR_c_299_n 0.0176554f $X=1.2 $Y=2.265 $X2=0
+ $Y2=0
cc_141 N_A_211_369#_c_143_n N_VPWR_c_300_n 0.016801f $X=1.2 $Y=2.265 $X2=0 $Y2=0
cc_142 N_A_211_369#_c_144_n N_VPWR_c_300_n 0.00270145f $X=1.682 $Y=1.8 $X2=0
+ $Y2=0
cc_143 N_A_211_369#_c_143_n N_VPWR_c_301_n 0.0234344f $X=1.2 $Y=2.265 $X2=0
+ $Y2=0
cc_144 N_A_211_369#_c_144_n N_VPWR_c_301_n 0.0237891f $X=1.682 $Y=1.8 $X2=0
+ $Y2=0
cc_145 N_A_211_369#_M1007_d N_VPWR_c_298_n 0.00425925f $X=1.055 $Y=1.845 $X2=0
+ $Y2=0
cc_146 N_A_211_369#_c_143_n N_VPWR_c_298_n 0.00961964f $X=1.2 $Y=2.265 $X2=0
+ $Y2=0
cc_147 N_A_211_369#_c_144_n N_VPWR_c_298_n 0.00619214f $X=1.682 $Y=1.8 $X2=0
+ $Y2=0
cc_148 N_A_211_369#_c_144_n N_Z_c_350_n 0.0355366f $X=1.682 $Y=1.8 $X2=0 $Y2=0
cc_149 N_A_211_369#_c_140_n N_Z_c_350_n 0.0513857f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_211_369#_c_141_n N_Z_c_350_n 0.00687776f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_211_369#_c_142_n N_VGND_c_377_n 0.0178712f $X=2.58 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_197_n N_VPWR_M1001_d 0.00346171f $X=0.657 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_153 N_A_27_47#_c_206_n N_VPWR_c_299_n 0.0223193f $X=0.26 $Y=2.22 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_197_n N_VPWR_c_299_n 0.0168404f $X=0.657 $Y=1.785 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_c_206_n N_VPWR_c_302_n 0.0176987f $X=0.26 $Y=2.22 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_197_n N_VPWR_c_302_n 0.00204391f $X=0.657 $Y=1.785 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_195_n N_VPWR_c_303_n 0.00429453f $X=3.025 $Y=1.41 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_M1001_s N_VPWR_c_298_n 0.00247737f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_195_n N_VPWR_c_298_n 0.00850698f $X=3.025 $Y=1.41 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_206_n N_VPWR_c_298_n 0.00983733f $X=0.26 $Y=2.22 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_197_n N_VPWR_c_298_n 0.00516598f $X=0.657 $Y=1.785 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_194_n Z 6.56308e-19 $X=3 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_195_n N_Z_c_350_n 0.0671013f $X=3.025 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_202_n N_Z_c_350_n 0.0050271f $X=2.915 $Y=0.82 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_204_n N_Z_c_350_n 0.016899f $X=3.03 $Y=0.82 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_194_n N_Z_c_346_n 0.0085086f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_194_n Z 0.00115211f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_195_n Z 0.0137245f $X=3.025 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_204_n Z 0.0340861f $X=3.03 $Y=0.82 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_197_n N_VGND_M1005_d 0.00124624f $X=0.657 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_171 N_A_27_47#_c_223_n N_VGND_M1005_d 0.0042757f $X=1.065 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_172 N_A_27_47#_c_198_n N_VGND_M1005_d 0.00176688f $X=0.79 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_173 N_A_27_47#_c_202_n N_VGND_M1002_s 0.00313199f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_196_n N_VGND_c_372_n 0.0149234f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_198_n N_VGND_c_372_n 0.00263331f $X=0.79 $Y=0.72 $X2=0 $Y2=0
cc_176 N_A_27_47#_M1005_s N_VGND_c_374_n 0.00288498f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_196_n N_VGND_c_374_n 0.00962926f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_223_n N_VGND_c_374_n 0.00439315f $X=1.065 $Y=0.72 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_198_n N_VGND_c_374_n 0.00640771f $X=0.79 $Y=0.72 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_199_n N_VGND_c_374_n 0.0353877f $X=1.96 $Y=0.36 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_200_n N_VGND_c_374_n 0.00635703f $X=1.235 $Y=0.36 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_202_n N_VGND_c_374_n 0.00653798f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_204_n N_VGND_c_374_n 6.57368e-19 $X=3.03 $Y=0.82 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_196_n N_VGND_c_375_n 0.0127118f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_198_n N_VGND_c_375_n 0.0242074f $X=0.79 $Y=0.72 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_200_n N_VGND_c_375_n 0.0161129f $X=1.235 $Y=0.36 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_223_n N_VGND_c_376_n 0.0025586f $X=1.065 $Y=0.72 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_199_n N_VGND_c_376_n 0.0627f $X=1.96 $Y=0.36 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_200_n N_VGND_c_376_n 0.0119068f $X=1.235 $Y=0.36 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_202_n N_VGND_c_376_n 0.00249653f $X=2.915 $Y=0.82 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_194_n N_VGND_c_377_n 0.0219108f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_199_n N_VGND_c_377_n 0.0193047f $X=1.96 $Y=0.36 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_201_n N_VGND_c_377_n 0.00828285f $X=2.067 $Y=0.735 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_202_n N_VGND_c_377_n 0.0311374f $X=2.915 $Y=0.82 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_204_n N_VGND_c_377_n 0.0120156f $X=3.03 $Y=0.82 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_202_n A_543_47# 9.99318e-19 $X=2.915 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_197 N_VPWR_c_298_n A_411_297# 0.0095846f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_198 N_VPWR_c_298_n N_Z_M1004_d 0.00320814f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_301_n N_Z_c_350_n 0.0193455f $X=1.72 $Y=2.26 $X2=0 $Y2=0
cc_200 N_VPWR_c_303_n N_Z_c_350_n 0.0787848f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_201 N_VPWR_c_298_n N_Z_c_350_n 0.0449787f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_202 N_VPWR_c_303_n N_Z_c_348_n 0.0190186f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_203 N_VPWR_c_298_n N_Z_c_348_n 0.0103877f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_204 A_411_297# N_Z_c_350_n 0.0595985f $X=2.055 $Y=1.485 $X2=0.69 $Y2=2.72
cc_205 N_Z_c_346_n N_VGND_c_373_n 0.0230657f $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_206 N_Z_M1000_d N_VGND_c_374_n 0.00964791f $X=3.075 $Y=0.235 $X2=0 $Y2=0
cc_207 N_Z_c_346_n N_VGND_c_374_n 0.0126215f $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_208 N_VGND_c_377_n A_543_47# 0.00106602f $X=3.085 $Y=0.24 $X2=-0.19 $Y2=-0.24
