* NGSPICE file created from sky130_fd_sc_hdll__buf_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__buf_4 A VGND VNB VPB VPWR X
M1000 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=8.5e+11p ps=7.7e+06u
M1001 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=4.16e+11p pd=3.88e+06u as=5.85e+11p ps=5.7e+06u
M1002 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1007 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

