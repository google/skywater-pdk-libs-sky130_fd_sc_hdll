* File: sky130_fd_sc_hdll__dlrtn_4.pex.spice
* Created: Wed Sep  2 08:29:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%GATE_N 4 5 7 8 10 13 19 22 24
c39 19 0 2.42713e-19 $X=0.23 $Y=1.19
c40 13 0 3.98209e-20 $X=0.52 $Y=0.805
r41 22 25 39.7811 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.3 $Y=1.235
+ $X2=0.3 $Y2=1.4
r42 22 24 39.7811 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.3 $Y=1.235
+ $X2=0.3 $Y2=1.07
r43 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.3
+ $Y=1.235 $X2=0.3 $Y2=1.235
r44 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r45 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r46 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r47 4 5 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.33 $Y=1.665
+ $X2=0.495 $Y2=1.665
r48 4 25 59.9997 $w=2.1e-07 $l=1.9e-07 $layer=POLY_cond $X=0.33 $Y=1.59 $X2=0.33
+ $Y2=1.4
r49 1 13 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.33 $Y=0.805
+ $X2=0.52 $Y2=0.805
r50 1 24 59.9997 $w=2.1e-07 $l=1.9e-07 $layer=POLY_cond $X=0.33 $Y=0.88 $X2=0.33
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%A_27_363# 1 2 9 13 15 18 20 22 23 28 30 31
+ 32 36 37 39 42 44 45 48 50 52 53 59 60 64
c161 59 0 1.0603e-19 $X=3.365 $Y=1.87
c162 52 0 2.45073e-19 $X=3.22 $Y=1.87
c163 50 0 1.14507e-19 $X=3.21 $Y=0.915
c164 48 0 2.17725e-19 $X=2.945 $Y=0.9
c165 42 0 1.26282e-19 $X=3.21 $Y=1.575
c166 23 0 1.93796e-19 $X=0.965 $Y=1.59
c167 20 0 8.68433e-20 $X=3.42 $Y=1.99
c168 13 0 2.2873e-20 $X=0.965 $Y=1.74
c169 9 0 2.60437e-20 $X=0.94 $Y=0.445
r170 60 72 4.25306 $w=4.18e-07 $l=1.55e-07 $layer=LI1_cond $X=3.365 $Y=1.785
+ $X2=3.21 $Y2=1.785
r171 60 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.425
+ $Y=1.74 $X2=3.425 $Y2=1.74
r172 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.365 $Y=1.87
+ $X2=3.365 $Y2=1.87
r173 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=1.87
+ $X2=0.72 $Y2=1.87
r174 53 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.865 $Y=1.87
+ $X2=0.72 $Y2=1.87
r175 52 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.22 $Y=1.87
+ $X2=3.365 $Y2=1.87
r176 52 53 2.9146 $w=1.4e-07 $l=2.355e-06 $layer=MET1_cond $X=3.22 $Y=1.87
+ $X2=0.865 $Y2=1.87
r177 47 50 8.48326 $w=3.58e-07 $l=2.65e-07 $layer=LI1_cond $X=2.945 $Y=0.915
+ $X2=3.21 $Y2=0.915
r178 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.945
+ $Y=0.9 $X2=2.945 $Y2=0.9
r179 42 72 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=3.21 $Y=1.575
+ $X2=3.21 $Y2=1.785
r180 41 50 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=3.21 $Y2=0.915
r181 41 42 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=3.21 $Y2=1.575
r182 40 64 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.81 $Y=1.235
+ $X2=0.94 $Y2=1.235
r183 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.235 $X2=0.81 $Y2=1.235
r184 37 56 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.795
+ $X2=0.75 $Y2=1.88
r185 37 39 22.2541 $w=2.88e-07 $l=5.6e-07 $layer=LI1_cond $X=0.75 $Y=1.795
+ $X2=0.75 $Y2=1.235
r186 36 45 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=0.75 $Y=1.215
+ $X2=0.75 $Y2=1.07
r187 36 39 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=0.75 $Y=1.215
+ $X2=0.75 $Y2=1.235
r188 34 45 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.69 $Y=0.805
+ $X2=0.69 $Y2=1.07
r189 33 44 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=1.88
+ $X2=0.24 $Y2=1.88
r190 32 56 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.75 $Y2=1.88
r191 32 33 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.395 $Y2=1.88
r192 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.69 $Y2=0.805
r193 30 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.395 $Y2=0.72
r194 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.31 $Y=0.635
+ $X2=0.395 $Y2=0.72
r195 26 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.31 $Y=0.635
+ $X2=0.31 $Y2=0.445
r196 20 69 48.3784 $w=2.91e-07 $l=2.52488e-07 $layer=POLY_cond $X=3.42 $Y=1.99
+ $X2=3.425 $Y2=1.74
r197 20 22 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.42 $Y=1.99
+ $X2=3.42 $Y2=2.275
r198 16 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=0.735
+ $X2=2.945 $Y2=0.9
r199 16 18 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.945 $Y=0.735
+ $X2=2.945 $Y2=0.415
r200 13 23 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=1.59
r201 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r202 11 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.37
+ $X2=0.94 $Y2=1.235
r203 11 23 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.94 $Y=1.37
+ $X2=0.94 $Y2=1.59
r204 7 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.1
+ $X2=0.94 $Y2=1.235
r205 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.94 $Y=1.1 $X2=0.94
+ $Y2=0.445
r206 2 44 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r207 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%D 2 3 5 8 10 11 12
c45 12 0 5.01492e-20 $X=1.61 $Y=1.19
c46 2 0 1.74491e-19 $X=1.955 $Y=1.67
r47 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.16 $X2=1.6 $Y2=1.16
r48 10 15 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.855 $Y=1.16
+ $X2=1.6 $Y2=1.16
r49 10 11 3.18546 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.855 $Y=1.16
+ $X2=1.955 $Y2=1.16
r50 6 11 33.332 $w=1.75e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.955 $Y2=1.16
r51 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.98 $Y=0.995 $X2=1.98
+ $Y2=0.445
r52 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.955 $Y=1.77
+ $X2=1.955 $Y2=2.165
r53 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.955 $Y=1.67 $X2=1.955
+ $Y2=1.77
r54 1 11 33.332 $w=1.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.325
+ $X2=1.955 $Y2=1.16
r55 1 2 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=1.955 $Y=1.325
+ $X2=1.955 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%A_319_369# 1 2 8 9 11 14 17 20 23 27 30 32
c78 32 0 1.14507e-19 $X=2.4 $Y=0.765
c79 30 0 1.2579e-19 $X=2.4 $Y=0.93
c80 17 0 1.74491e-19 $X=1.72 $Y=1.99
r81 30 33 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=0.93 $X2=2.4
+ $Y2=1.095
r82 30 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=0.93 $X2=2.4
+ $Y2=0.765
r83 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=0.93 $X2=2.4 $Y2=0.93
r84 27 29 12.2997 $w=3.67e-07 $l=4.63249e-07 $layer=LI1_cond $X=2.03 $Y=0.72
+ $X2=2.4 $Y2=0.93
r85 26 27 8.64305 $w=3.67e-07 $l=2.6e-07 $layer=LI1_cond $X=1.77 $Y=0.72
+ $X2=2.03 $Y2=0.72
r86 20 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=1.495
+ $X2=2.03 $Y2=1.58
r87 19 27 5.25812 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=2.03 $Y=1.095
+ $X2=2.03 $Y2=0.72
r88 19 20 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.03 $Y=1.095 $X2=2.03
+ $Y2=1.495
r89 15 23 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.72 $Y=1.58
+ $X2=2.03 $Y2=1.58
r90 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.72 $Y2=1.99
r91 14 32 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.425 $Y=0.445
+ $X2=2.425 $Y2=0.765
r92 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=1.77
+ $X2=2.425 $Y2=2.165
r93 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.425 $Y=1.67 $X2=2.425
+ $Y2=1.77
r94 8 33 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.67
+ $X2=2.425 $Y2=1.095
r95 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.845 $X2=1.72 $Y2=1.99
r96 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.235 $X2=1.77 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%A_203_47# 1 2 8 9 11 12 16 20 24 26 27 30
+ 33 36 40
c114 40 0 3.47682e-19 $X=2.87 $Y=1.44
c115 9 0 1.43299e-19 $X=2.95 $Y=1.99
c116 2 0 1.13552e-19 $X=1.055 $Y=1.815
r117 39 41 43.3814 $w=3.15e-07 $l=1.95e-07 $layer=POLY_cond $X=2.892 $Y=1.44
+ $X2=2.892 $Y2=1.635
r118 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.44 $X2=2.87 $Y2=1.44
r119 36 39 21.9826 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=2.892 $Y=1.32
+ $X2=2.892 $Y2=1.44
r120 33 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.81 $Y=1.53
+ $X2=2.81 $Y2=1.53
r121 30 46 5.20126 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.53 $X2=1.2
+ $Y2=1.445
r122 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.18 $Y=1.53
+ $X2=1.18 $Y2=1.53
r123 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.325 $Y=1.53
+ $X2=1.18 $Y2=1.53
r124 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.665 $Y=1.53
+ $X2=2.81 $Y2=1.53
r125 26 27 1.65841 $w=1.4e-07 $l=1.34e-06 $layer=MET1_cond $X=2.665 $Y=1.53
+ $X2=1.325 $Y2=1.53
r126 22 30 2.13415 $w=2.68e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=1.58 $X2=1.2
+ $Y2=1.53
r127 22 24 16.2196 $w=2.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.2 $Y=1.58 $X2=1.2
+ $Y2=1.96
r128 20 46 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=1.15 $Y=0.445
+ $X2=1.15 $Y2=1.445
r129 14 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.465 $Y=1.245
+ $X2=3.465 $Y2=0.445
r130 13 36 20.1192 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=3.05 $Y=1.32
+ $X2=2.892 $Y2=1.32
r131 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.39 $Y=1.32
+ $X2=3.465 $Y2=1.245
r132 12 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.39 $Y=1.32
+ $X2=3.05 $Y2=1.32
r133 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.95 $Y=1.99
+ $X2=2.95 $Y2=2.275
r134 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.95 $Y=1.89 $X2=2.95
+ $Y2=1.99
r135 8 41 84.5522 $w=2e-07 $l=2.55e-07 $layer=POLY_cond $X=2.95 $Y=1.89 $X2=2.95
+ $Y2=1.635
r136 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r137 1 20 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.15 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%A_750_21# 1 2 9 11 13 14 16 17 19 20 22 23
+ 25 26 28 29 31 32 34 35 37 38 45 48 51 54 55 57 60 62 65 74
c157 74 0 1.09327e-19 $X=7.13 $Y=1.202
c158 55 0 1.1645e-19 $X=5.725 $Y=1.2
c159 9 0 1.26282e-19 $X=3.825 $Y=0.445
r160 74 75 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.13 $Y=1.202
+ $X2=7.155 $Y2=1.202
r161 73 74 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.71 $Y=1.202
+ $X2=7.13 $Y2=1.202
r162 72 73 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.685 $Y=1.202
+ $X2=6.71 $Y2=1.202
r163 71 72 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=6.215 $Y=1.202
+ $X2=6.685 $Y2=1.202
r164 70 71 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.19 $Y=1.202
+ $X2=6.215 $Y2=1.202
r165 67 68 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.745 $Y=1.202
+ $X2=5.77 $Y2=1.202
r166 64 65 7.4145 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.04 $Y=1.7
+ $X2=5.175 $Y2=1.7
r167 62 64 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.025 $Y=1.7
+ $X2=5.04 $Y2=1.7
r168 61 62 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=4.635 $Y=1.7
+ $X2=5.025 $Y2=1.7
r169 58 70 15.6324 $w=3.7e-07 $l=1.2e-07 $layer=POLY_cond $X=6.07 $Y=1.202
+ $X2=6.19 $Y2=1.202
r170 58 68 39.0811 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=6.07 $Y=1.202
+ $X2=5.77 $Y2=1.202
r171 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.07
+ $Y=1.16 $X2=6.07 $Y2=1.16
r172 55 57 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=5.725 $Y=1.2
+ $X2=6.07 $Y2=1.2
r173 53 55 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.64 $Y=1.325
+ $X2=5.725 $Y2=1.2
r174 53 54 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.64 $Y=1.325
+ $X2=5.64 $Y2=1.535
r175 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.555 $Y=1.62
+ $X2=5.64 $Y2=1.535
r176 51 65 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.555 $Y=1.62
+ $X2=5.175 $Y2=1.62
r177 48 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.635 $Y=1.535
+ $X2=4.635 $Y2=1.7
r178 48 60 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.635 $Y=1.535
+ $X2=4.635 $Y2=0.825
r179 43 60 7.25185 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=0.66
+ $X2=4.62 $Y2=0.825
r180 43 45 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.62 $Y=0.66
+ $X2=4.62 $Y2=0.38
r181 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=1.7 $X2=4.105 $Y2=1.7
r182 38 61 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=1.7
+ $X2=4.635 $Y2=1.7
r183 38 40 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.55 $Y=1.7
+ $X2=4.105 $Y2=1.7
r184 35 75 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.155 $Y=1.41
+ $X2=7.155 $Y2=1.202
r185 35 37 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.155 $Y=1.41
+ $X2=7.155 $Y2=1.985
r186 32 74 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.13 $Y=0.995
+ $X2=7.13 $Y2=1.202
r187 32 34 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.13 $Y=0.995
+ $X2=7.13 $Y2=0.56
r188 29 73 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.71 $Y=0.995
+ $X2=6.71 $Y2=1.202
r189 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.71 $Y=0.995
+ $X2=6.71 $Y2=0.56
r190 26 72 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.685 $Y=1.41
+ $X2=6.685 $Y2=1.202
r191 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.685 $Y=1.41
+ $X2=6.685 $Y2=1.985
r192 23 71 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.215 $Y=1.41
+ $X2=6.215 $Y2=1.202
r193 23 25 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.215 $Y=1.41
+ $X2=6.215 $Y2=1.985
r194 20 70 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.19 $Y=0.995
+ $X2=6.19 $Y2=1.202
r195 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.19 $Y=0.995
+ $X2=6.19 $Y2=0.56
r196 17 68 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.77 $Y=0.995
+ $X2=5.77 $Y2=1.202
r197 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.77 $Y=0.995
+ $X2=5.77 $Y2=0.56
r198 14 67 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.745 $Y=1.41
+ $X2=5.745 $Y2=1.202
r199 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.745 $Y=1.41
+ $X2=5.745 $Y2=1.985
r200 11 41 53.3563 $w=3.12e-07 $l=3.38452e-07 $layer=POLY_cond $X=3.9 $Y=1.99
+ $X2=4.005 $Y2=1.7
r201 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.9 $Y=1.99
+ $X2=3.9 $Y2=2.275
r202 7 41 78.6992 $w=3.12e-07 $l=5.07075e-07 $layer=POLY_cond $X=3.825 $Y=1.275
+ $X2=4.005 $Y2=1.7
r203 7 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.825 $Y=1.275
+ $X2=3.825 $Y2=0.445
r204 2 64 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=4.895
+ $Y=1.485 $X2=5.04 $Y2=1.755
r205 1 45 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.495
+ $Y=0.235 $X2=4.62 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%A_604_47# 1 2 7 9 11 14 16 18 22 27 29 30
+ 32 33
c91 30 0 2.92347e-19 $X=3.85 $Y=1.16
c92 29 0 1.43299e-19 $X=3.765 $Y=2.165
c93 9 0 1.92496e-19 $X=4.805 $Y=1.41
r94 35 36 9.46122 $w=2.45e-07 $l=1.9e-07 $layer=LI1_cond $X=3.575 $Y=1.16
+ $X2=3.765 $Y2=1.16
r95 33 39 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=4.295 $Y=1.16
+ $X2=4.295 $Y2=1.25
r96 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.16 $X2=4.295 $Y2=1.16
r97 30 36 3.97745 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=1.16
+ $X2=3.765 $Y2=1.16
r98 30 32 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.85 $Y=1.16
+ $X2=4.295 $Y2=1.16
r99 28 36 2.87745 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=1.325
+ $X2=3.765 $Y2=1.16
r100 28 29 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.765 $Y=1.325
+ $X2=3.765 $Y2=2.165
r101 27 35 2.87745 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=1.16
r102 26 27 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.575 $Y=0.565
+ $X2=3.575 $Y2=0.995
r103 22 26 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=3.49 $Y=0.422
+ $X2=3.575 $Y2=0.565
r104 22 24 11.5244 $w=2.83e-07 $l=2.85e-07 $layer=LI1_cond $X=3.49 $Y=0.422
+ $X2=3.205 $Y2=0.422
r105 18 29 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.68 $Y=2.275
+ $X2=3.765 $Y2=2.165
r106 18 20 25.93 $w=2.18e-07 $l=4.95e-07 $layer=LI1_cond $X=3.68 $Y=2.275
+ $X2=3.185 $Y2=2.275
r107 16 17 29.1618 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=4.805 $Y=1.25
+ $X2=4.805 $Y2=1.175
r108 14 17 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.83 $Y=0.56
+ $X2=4.83 $Y2=1.175
r109 9 16 53.8601 $w=2e-07 $l=1.6e-07 $layer=POLY_cond $X=4.805 $Y=1.41
+ $X2=4.805 $Y2=1.25
r110 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.805 $Y=1.41
+ $X2=4.805 $Y2=1.985
r111 8 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.43 $Y=1.25
+ $X2=4.295 $Y2=1.25
r112 7 16 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=4.705 $Y=1.25
+ $X2=4.805 $Y2=1.25
r113 7 8 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=4.705 $Y=1.25
+ $X2=4.43 $Y2=1.25
r114 2 20 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.065 $X2=3.185 $Y2=2.275
r115 1 24 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.235 $X2=3.205 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%RESET_B 1 3 4 6 7
r34 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.16 $X2=5.25 $Y2=1.16
r35 4 10 51.486 $w=2.55e-07 $l=2.62202e-07 $layer=POLY_cond $X=5.275 $Y=1.41
+ $X2=5.25 $Y2=1.16
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.275 $Y=1.41
+ $X2=5.275 $Y2=1.985
r37 1 10 39.2931 $w=2.55e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.25 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.235 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%VPWR 1 2 3 4 5 6 21 25 30 33 37 42 46 47
+ 49 50 52 53 54 56 61 85 86 89 92 97 100
c114 42 0 3.01823e-19 $X=5.51 $Y=1.97
c115 21 0 1.31521e-19 $X=0.73 $Y=2.22
r116 99 100 10.5224 $w=6.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.545 $Y=2.47
+ $X2=4.705 $Y2=2.47
r117 95 99 3.12409 $w=6.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.37 $Y=2.47
+ $X2=4.545 $Y2=2.47
r118 95 97 13.9143 $w=6.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.37 $Y=2.47
+ $X2=4.02 $Y2=2.47
r119 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r120 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r121 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r123 83 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r124 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r125 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r126 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r127 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r128 77 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r129 76 100 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=4.705 $Y2=2.72
r130 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r131 73 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r132 72 97 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.02 $Y2=2.72
r133 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r134 70 73 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r135 70 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r136 69 72 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r137 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r138 67 92 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.19 $Y2=2.72
r139 67 69 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.53 $Y2=2.72
r140 65 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 65 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r142 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 62 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.73 $Y2=2.72
r144 62 64 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r145 61 92 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.19 $Y2=2.72
r146 61 64 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.15 $Y2=2.72
r147 56 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.73 $Y2=2.72
r148 56 58 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.23 $Y2=2.72
r149 54 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r150 54 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r151 52 82 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.255 $Y=2.72
+ $X2=7.13 $Y2=2.72
r152 52 53 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=7.255 $Y=2.72
+ $X2=7.382 $Y2=2.72
r153 51 85 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.51 $Y=2.72 $X2=7.59
+ $Y2=2.72
r154 51 53 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=7.51 $Y=2.72
+ $X2=7.382 $Y2=2.72
r155 49 79 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.315 $Y=2.72
+ $X2=6.21 $Y2=2.72
r156 49 50 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.315 $Y=2.72
+ $X2=6.45 $Y2=2.72
r157 48 82 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=7.13 $Y2=2.72
r158 48 50 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=6.45 $Y2=2.72
r159 46 76 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.29 $Y2=2.72
r160 46 47 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.495 $Y2=2.72
r161 45 79 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=6.21 $Y2=2.72
r162 45 47 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=5.495 $Y2=2.72
r163 42 44 6.40424 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.51 $Y=1.97
+ $X2=5.51 $Y2=2.15
r164 37 40 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=7.382 $Y=1.66
+ $X2=7.382 $Y2=2.34
r165 35 53 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.382 $Y=2.635
+ $X2=7.382 $Y2=2.72
r166 35 40 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=7.382 $Y=2.635
+ $X2=7.382 $Y2=2.34
r167 31 50 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=2.635
+ $X2=6.45 $Y2=2.72
r168 31 33 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.45 $Y=2.635
+ $X2=6.45 $Y2=2
r169 30 44 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=5.495 $Y=2.34
+ $X2=5.495 $Y2=2.15
r170 28 47 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=2.635
+ $X2=5.495 $Y2=2.72
r171 28 30 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.495 $Y=2.635
+ $X2=5.495 $Y2=2.34
r172 23 92 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r173 23 25 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2
r174 19 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r175 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.22
r176 6 40 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.485 $X2=7.39 $Y2=2.34
r177 6 37 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.485 $X2=7.39 $Y2=1.66
r178 5 33 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.305
+ $Y=1.485 $X2=6.45 $Y2=2
r179 4 42 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.51 $Y2=1.97
r180 4 30 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.51 $Y2=2.34
r181 3 99 300 $w=1.7e-07 $l=6.62156e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.065 $X2=4.545 $Y2=2.3
r182 2 25 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.845 $X2=2.19 $Y2=2
r183 1 21 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%Q 1 2 3 4 15 19 21 23 24 27 29 31 34 35 38
+ 39 42
r72 47 49 1.33333 $w=7.32e-07 $l=8e-08 $layer=LI1_cond $X=6.835 $Y=1.58
+ $X2=6.835 $Y2=1.66
r73 42 47 6.5 $w=7.32e-07 $l=3.9e-07 $layer=LI1_cond $X=6.835 $Y=1.19 $X2=6.835
+ $Y2=1.58
r74 42 44 6.16667 $w=7.32e-07 $l=3.7e-07 $layer=LI1_cond $X=6.835 $Y=1.19
+ $X2=6.835 $Y2=0.82
r75 38 39 5.15594 $w=2.98e-07 $l=1.25e-07 $layer=LI1_cond $X=5.995 $Y=2
+ $X2=5.995 $Y2=1.875
r76 34 35 3.0866 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=2.34 $X2=5.98
+ $Y2=2.255
r77 29 49 3.8083 $w=7.32e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.92 $Y=1.665
+ $X2=6.835 $Y2=1.66
r78 29 31 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.92 $Y=1.665
+ $X2=6.92 $Y2=2.34
r79 25 44 5.14164 $w=7.32e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.92 $Y=0.735
+ $X2=6.835 $Y2=0.82
r80 25 27 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=6.92 $Y=0.735
+ $X2=6.92 $Y2=0.38
r81 23 44 9.61685 $w=1.7e-07 $l=4.3e-07 $layer=LI1_cond $X=6.405 $Y=0.82
+ $X2=6.835 $Y2=0.82
r82 23 24 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.405 $Y=0.82
+ $X2=6.195 $Y2=0.82
r83 22 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.145 $Y=1.58
+ $X2=6.02 $Y2=1.58
r84 21 47 9.61685 $w=1.7e-07 $l=4.3e-07 $layer=LI1_cond $X=6.405 $Y=1.58
+ $X2=6.835 $Y2=1.58
r85 21 22 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.405 $Y=1.58
+ $X2=6.145 $Y2=1.58
r86 19 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=1.665
+ $X2=6.02 $Y2=1.58
r87 19 39 9.68052 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=6.02 $Y=1.665
+ $X2=6.02 $Y2=1.875
r88 17 38 0.960369 $w=2.98e-07 $l=2.5e-08 $layer=LI1_cond $X=5.995 $Y=2.025
+ $X2=5.995 $Y2=2
r89 17 35 8.8354 $w=2.98e-07 $l=2.3e-07 $layer=LI1_cond $X=5.995 $Y=2.025
+ $X2=5.995 $Y2=2.255
r90 13 24 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=6.005 $Y=0.735
+ $X2=6.195 $Y2=0.82
r91 13 15 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=6.005 $Y=0.735
+ $X2=6.005 $Y2=0.38
r92 4 49 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.775
+ $Y=1.485 $X2=6.92 $Y2=1.66
r93 4 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.775
+ $Y=1.485 $X2=6.92 $Y2=2.34
r94 3 41 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=1.485 $X2=5.98 $Y2=1.66
r95 3 38 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=1.485 $X2=5.98 $Y2=2
r96 3 34 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=1.485 $X2=5.98 $Y2=2.34
r97 2 27 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.785
+ $Y=0.235 $X2=6.92 $Y2=0.38
r98 1 15 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.845
+ $Y=0.235 $X2=5.98 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_4%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45
+ 47 48 50 51 52 54 59 64 83 84 87 90 93
c119 84 0 3.98209e-20 $X=7.59 $Y=0
r120 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r121 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r122 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r123 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r124 81 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r125 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r126 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r127 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r128 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r129 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r130 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r131 72 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r132 71 74 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r133 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r134 69 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.035
+ $Y2=0
r135 69 71 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.37
+ $Y2=0
r136 68 94 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r137 68 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r138 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r139 65 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.19
+ $Y2=0
r140 65 67 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.53 $Y2=0
r141 64 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.87 $Y=0 $X2=4.035
+ $Y2=0
r142 64 67 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=3.87 $Y=0 $X2=2.53
+ $Y2=0
r143 63 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r144 63 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r145 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r146 60 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.73
+ $Y2=0
r147 60 62 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r148 59 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.19
+ $Y2=0
r149 59 62 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=1.15 $Y2=0
r150 54 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.73
+ $Y2=0
r151 54 56 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=0
+ $X2=0.23 $Y2=0
r152 52 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r153 52 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r154 50 80 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.255 $Y=0
+ $X2=7.13 $Y2=0
r155 50 51 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.255 $Y=0 $X2=7.36
+ $Y2=0
r156 49 83 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.465 $Y=0
+ $X2=7.59 $Y2=0
r157 49 51 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.465 $Y=0 $X2=7.36
+ $Y2=0
r158 47 77 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=0
+ $X2=6.21 $Y2=0
r159 47 48 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.375 $Y=0 $X2=6.48
+ $Y2=0
r160 46 80 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=6.585 $Y=0
+ $X2=7.13 $Y2=0
r161 46 48 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.585 $Y=0 $X2=6.48
+ $Y2=0
r162 44 74 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.29
+ $Y2=0
r163 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.48
+ $Y2=0
r164 43 77 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.645 $Y=0 $X2=6.21
+ $Y2=0
r165 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.645 $Y=0 $X2=5.48
+ $Y2=0
r166 39 51 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r167 39 41 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.38
r168 35 48 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.48 $Y=0.085
+ $X2=6.48 $Y2=0
r169 35 37 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=6.48 $Y=0.085
+ $X2=6.48 $Y2=0.38
r170 31 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r171 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.38
r172 27 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0.085
+ $X2=4.035 $Y2=0
r173 27 29 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=0.085
+ $X2=4.035 $Y2=0.445
r174 23 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0
r175 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0.36
r176 19 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r177 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r178 6 41 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.205
+ $Y=0.235 $X2=7.34 $Y2=0.38
r179 5 37 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=6.265
+ $Y=0.235 $X2=6.46 $Y2=0.38
r180 4 33 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=5.31
+ $Y=0.235 $X2=5.48 $Y2=0.38
r181 3 29 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.035 $Y2=0.445
r182 2 25 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.36
r183 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

