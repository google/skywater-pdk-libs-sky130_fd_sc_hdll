* File: sky130_fd_sc_hdll__and2b_1.pxi.spice
* Created: Wed Sep  2 08:21:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND2B_1%A_N N_A_N_c_57_n N_A_N_c_58_n N_A_N_M1000_g
+ N_A_N_M1006_g A_N A_N A_N N_A_N_c_56_n PM_SKY130_FD_SC_HDLL__AND2B_1%A_N
x_PM_SKY130_FD_SC_HDLL__AND2B_1%A_27_413# N_A_27_413#_M1006_d
+ N_A_27_413#_M1000_s N_A_27_413#_c_89_n N_A_27_413#_c_98_n N_A_27_413#_M1002_g
+ N_A_27_413#_c_90_n N_A_27_413#_M1003_g N_A_27_413#_c_99_n N_A_27_413#_c_100_n
+ N_A_27_413#_c_101_n N_A_27_413#_c_92_n N_A_27_413#_c_93_n N_A_27_413#_c_94_n
+ N_A_27_413#_c_95_n N_A_27_413#_c_96_n PM_SKY130_FD_SC_HDLL__AND2B_1%A_27_413#
x_PM_SKY130_FD_SC_HDLL__AND2B_1%B N_B_c_160_n N_B_M1007_g N_B_M1001_g B
+ PM_SKY130_FD_SC_HDLL__AND2B_1%B
x_PM_SKY130_FD_SC_HDLL__AND2B_1%A_225_413# N_A_225_413#_M1003_s
+ N_A_225_413#_M1002_d N_A_225_413#_c_191_n N_A_225_413#_M1005_g
+ N_A_225_413#_c_192_n N_A_225_413#_M1004_g N_A_225_413#_c_197_n
+ N_A_225_413#_c_193_n N_A_225_413#_c_194_n N_A_225_413#_c_195_n
+ N_A_225_413#_c_215_n PM_SKY130_FD_SC_HDLL__AND2B_1%A_225_413#
x_PM_SKY130_FD_SC_HDLL__AND2B_1%VPWR N_VPWR_M1000_d N_VPWR_M1007_d
+ N_VPWR_c_253_n VPWR N_VPWR_c_254_n N_VPWR_c_255_n N_VPWR_c_252_n
+ N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_259_n
+ PM_SKY130_FD_SC_HDLL__AND2B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__AND2B_1%X N_X_M1004_d N_X_M1005_d X X X N_X_c_291_n
+ N_X_c_290_n PM_SKY130_FD_SC_HDLL__AND2B_1%X
x_PM_SKY130_FD_SC_HDLL__AND2B_1%VGND N_VGND_M1006_s N_VGND_M1001_d
+ N_VGND_c_308_n N_VGND_c_309_n N_VGND_c_310_n VGND N_VGND_c_311_n
+ N_VGND_c_312_n N_VGND_c_313_n N_VGND_c_314_n
+ PM_SKY130_FD_SC_HDLL__AND2B_1%VGND
cc_1 VNB N_A_N_M1006_g 0.0385037f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A_N 0.0247288f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_A_N_c_56_n 0.035774f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_4 VNB N_A_27_413#_c_89_n 0.0111595f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_A_27_413#_c_90_n 0.0165653f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_6 VNB N_A_27_413#_M1003_g 0.0220462f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_7 VNB N_A_27_413#_c_92_n 0.00413025f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.19
cc_8 VNB N_A_27_413#_c_93_n 0.00377231f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.53
cc_9 VNB N_A_27_413#_c_94_n 0.00476028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_413#_c_95_n 0.00673088f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_413#_c_96_n 0.0431289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_160_n 0.0209835f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_13 VNB N_B_M1001_g 0.0386626f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_14 VNB N_A_225_413#_c_191_n 0.0272763f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_15 VNB N_A_225_413#_c_192_n 0.0197069f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_16 VNB N_A_225_413#_c_193_n 0.00538911f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_17 VNB N_A_225_413#_c_194_n 0.0168405f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=0.995
cc_18 VNB N_A_225_413#_c_195_n 0.00538806f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=0.85
cc_19 VNB N_VPWR_c_252_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB X 0.0240337f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_21 VNB N_X_c_290_n 0.0281254f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_22 VNB N_VGND_c_308_n 0.0114894f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_23 VNB N_VGND_c_309_n 0.0211579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_310_n 0.00319506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_311_n 0.0435704f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_26 VNB N_VGND_c_312_n 0.0232963f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_27 VNB N_VGND_c_313_n 0.187942f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.19
cc_28 VNB N_VGND_c_314_n 0.00702351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_A_N_c_57_n 0.042736f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_30 VPB N_A_N_c_58_n 0.0264662f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_31 VPB A_N 0.0149437f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_32 VPB N_A_N_c_56_n 0.00756804f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_33 VPB N_A_27_413#_c_89_n 0.0336024f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_34 VPB N_A_27_413#_c_98_n 0.0230839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_413#_c_99_n 0.00219961f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.325
cc_36 VPB N_A_27_413#_c_100_n 0.00861747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_413#_c_101_n 0.0109524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_413#_c_93_n 0.00955518f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.53
cc_39 VPB N_B_c_160_n 0.101141f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_40 VPB B 0.00737833f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_41 VPB N_A_225_413#_c_191_n 0.0367161f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_42 VPB N_A_225_413#_c_197_n 0.00640752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_225_413#_c_194_n 0.00812205f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=0.995
cc_44 VPB N_A_225_413#_c_195_n 0.00269355f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=0.85
cc_45 VPB N_VPWR_c_253_n 0.00285015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_254_n 0.015299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_255_n 0.0273184f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.19
cc_48 VPB N_VPWR_c_252_n 0.048528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_257_n 0.00580026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_258_n 0.0205261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_259_n 0.0196811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_X_c_291_n 0.0378767f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_53 VPB N_X_c_290_n 0.0144951f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_54 N_A_N_c_56_n N_A_27_413#_c_89_n 0.0116558f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_N_c_57_n N_A_27_413#_c_98_n 0.0116558f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_56 N_A_N_c_58_n N_A_27_413#_c_98_n 0.0130435f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_57 N_A_N_c_58_n N_A_27_413#_c_99_n 0.00550801f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_58 N_A_N_c_57_n N_A_27_413#_c_100_n 0.0126834f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_59 N_A_N_c_58_n N_A_27_413#_c_100_n 0.010017f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_60 A_N N_A_27_413#_c_100_n 0.00808417f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_61 A_N N_A_27_413#_c_101_n 0.0158932f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_62 N_A_N_c_56_n N_A_27_413#_c_101_n 6.27406e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_N_M1006_g N_A_27_413#_c_92_n 0.00520726f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_64 A_N N_A_27_413#_c_92_n 0.00267491f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_65 A_N N_A_27_413#_c_93_n 0.0302442f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_66 N_A_N_c_56_n N_A_27_413#_c_93_n 0.00879718f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_N_M1006_g N_A_27_413#_c_95_n 0.00323242f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_68 A_N N_A_27_413#_c_95_n 0.023149f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_69 N_A_N_M1006_g N_A_27_413#_c_96_n 0.0116558f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_70 A_N N_A_27_413#_c_96_n 2.43043e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_71 N_A_N_c_57_n N_A_225_413#_c_197_n 2.14247e-19 $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_72 N_A_N_c_58_n N_A_225_413#_c_197_n 5.64081e-19 $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_73 N_A_N_c_58_n N_VPWR_c_253_n 0.0129778f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_74 N_A_N_c_58_n N_VPWR_c_254_n 0.00321743f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_75 N_A_N_c_58_n N_VPWR_c_252_n 0.00482954f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_76 N_A_N_M1006_g N_VGND_c_309_n 0.00511692f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_77 A_N N_VGND_c_309_n 0.0225521f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_78 N_A_N_c_56_n N_VGND_c_309_n 0.0010017f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_N_M1006_g N_VGND_c_311_n 0.00585385f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_80 N_A_N_M1006_g N_VGND_c_313_n 0.0130277f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_81 A_N N_VGND_c_313_n 0.00193939f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_82 N_A_27_413#_c_89_n N_B_c_160_n 0.0284197f $X=1.035 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_27_413#_c_98_n N_B_c_160_n 0.0109994f $X=1.035 $Y=1.99 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_27_413#_c_90_n N_B_c_160_n 0.0076604f $X=1.485 $Y=0.88 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_27_413#_M1003_g N_B_M1001_g 0.0350627f $X=1.56 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A_27_413#_c_96_n N_B_M1001_g 0.00236933f $X=1.33 $Y=0.97 $X2=0 $Y2=0
cc_87 N_A_27_413#_c_89_n N_A_225_413#_c_197_n 0.0102023f $X=1.035 $Y=1.89 $X2=0
+ $Y2=0
cc_88 N_A_27_413#_c_98_n N_A_225_413#_c_197_n 0.0112053f $X=1.035 $Y=1.99 $X2=0
+ $Y2=0
cc_89 N_A_27_413#_c_100_n N_A_225_413#_c_197_n 0.019338f $X=0.665 $Y=1.9 $X2=0
+ $Y2=0
cc_90 N_A_27_413#_c_93_n N_A_225_413#_c_197_n 0.0238327f $X=0.782 $Y=1.785 $X2=0
+ $Y2=0
cc_91 N_A_27_413#_c_90_n N_A_225_413#_c_193_n 0.00648153f $X=1.485 $Y=0.88 $X2=0
+ $Y2=0
cc_92 N_A_27_413#_M1003_g N_A_225_413#_c_193_n 0.00585979f $X=1.56 $Y=0.445
+ $X2=0 $Y2=0
cc_93 N_A_27_413#_c_94_n N_A_225_413#_c_193_n 0.00680418f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_94 N_A_27_413#_c_95_n N_A_225_413#_c_193_n 0.0106118f $X=1.115 $Y=0.97 $X2=0
+ $Y2=0
cc_95 N_A_27_413#_c_89_n N_A_225_413#_c_194_n 0.00818837f $X=1.035 $Y=1.89 $X2=0
+ $Y2=0
cc_96 N_A_27_413#_c_90_n N_A_225_413#_c_194_n 0.00651805f $X=1.485 $Y=0.88 $X2=0
+ $Y2=0
cc_97 N_A_27_413#_c_93_n N_A_225_413#_c_194_n 0.0206051f $X=0.782 $Y=1.785 $X2=0
+ $Y2=0
cc_98 N_A_27_413#_c_95_n N_A_225_413#_c_194_n 0.0315093f $X=1.115 $Y=0.97 $X2=0
+ $Y2=0
cc_99 N_A_27_413#_c_96_n N_A_225_413#_c_194_n 0.00854961f $X=1.33 $Y=0.97 $X2=0
+ $Y2=0
cc_100 N_A_27_413#_M1003_g N_A_225_413#_c_215_n 0.00564898f $X=1.56 $Y=0.445
+ $X2=0 $Y2=0
cc_101 N_A_27_413#_c_94_n N_A_225_413#_c_215_n 0.0163154f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_102 N_A_27_413#_c_95_n N_A_225_413#_c_215_n 0.00236721f $X=1.115 $Y=0.97
+ $X2=0 $Y2=0
cc_103 N_A_27_413#_c_96_n N_A_225_413#_c_215_n 0.00712003f $X=1.33 $Y=0.97 $X2=0
+ $Y2=0
cc_104 N_A_27_413#_c_98_n N_VPWR_c_253_n 0.00471342f $X=1.035 $Y=1.99 $X2=0
+ $Y2=0
cc_105 N_A_27_413#_c_99_n N_VPWR_c_253_n 0.0194103f $X=0.26 $Y=2.225 $X2=0 $Y2=0
cc_106 N_A_27_413#_c_100_n N_VPWR_c_253_n 0.0287524f $X=0.665 $Y=1.9 $X2=0 $Y2=0
cc_107 N_A_27_413#_c_99_n N_VPWR_c_254_n 0.010445f $X=0.26 $Y=2.225 $X2=0 $Y2=0
cc_108 N_A_27_413#_c_100_n N_VPWR_c_254_n 0.00252438f $X=0.665 $Y=1.9 $X2=0
+ $Y2=0
cc_109 N_A_27_413#_M1000_s N_VPWR_c_252_n 0.00388418f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_110 N_A_27_413#_c_98_n N_VPWR_c_252_n 0.0111846f $X=1.035 $Y=1.99 $X2=0 $Y2=0
cc_111 N_A_27_413#_c_99_n N_VPWR_c_252_n 0.00640243f $X=0.26 $Y=2.225 $X2=0
+ $Y2=0
cc_112 N_A_27_413#_c_100_n N_VPWR_c_252_n 0.00582594f $X=0.665 $Y=1.9 $X2=0
+ $Y2=0
cc_113 N_A_27_413#_c_98_n N_VPWR_c_258_n 0.00646924f $X=1.035 $Y=1.99 $X2=0
+ $Y2=0
cc_114 N_A_27_413#_M1003_g N_VGND_c_310_n 0.00199455f $X=1.56 $Y=0.445 $X2=0
+ $Y2=0
cc_115 N_A_27_413#_M1003_g N_VGND_c_311_n 0.00388886f $X=1.56 $Y=0.445 $X2=0
+ $Y2=0
cc_116 N_A_27_413#_c_94_n N_VGND_c_311_n 0.0140003f $X=0.73 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_27_413#_M1006_d N_VGND_c_313_n 0.00388065f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_118 N_A_27_413#_M1003_g N_VGND_c_313_n 0.00686811f $X=1.56 $Y=0.445 $X2=0
+ $Y2=0
cc_119 N_A_27_413#_c_94_n N_VGND_c_313_n 0.00898311f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_120 N_A_27_413#_c_95_n N_VGND_c_313_n 0.0114982f $X=1.115 $Y=0.97 $X2=0 $Y2=0
cc_121 N_A_27_413#_c_96_n N_VGND_c_313_n 0.00704017f $X=1.33 $Y=0.97 $X2=0 $Y2=0
cc_122 N_B_c_160_n N_A_225_413#_c_191_n 0.014875f $X=1.525 $Y=1.99 $X2=0 $Y2=0
cc_123 N_B_M1001_g N_A_225_413#_c_191_n 0.0220121f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_124 B N_A_225_413#_c_191_n 0.00340151f $X=1.985 $Y=1.745 $X2=0 $Y2=0
cc_125 N_B_M1001_g N_A_225_413#_c_192_n 0.0212992f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_126 N_B_c_160_n N_A_225_413#_c_197_n 0.0113795f $X=1.525 $Y=1.99 $X2=0 $Y2=0
cc_127 B N_A_225_413#_c_197_n 0.0211295f $X=1.985 $Y=1.745 $X2=0 $Y2=0
cc_128 N_B_M1001_g N_A_225_413#_c_193_n 0.00561396f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_129 N_B_c_160_n N_A_225_413#_c_194_n 0.0430771f $X=1.525 $Y=1.99 $X2=0 $Y2=0
cc_130 N_B_M1001_g N_A_225_413#_c_194_n 0.0147879f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_131 B N_A_225_413#_c_194_n 0.0360408f $X=1.985 $Y=1.745 $X2=0 $Y2=0
cc_132 B N_A_225_413#_c_195_n 0.0103329f $X=1.985 $Y=1.745 $X2=0 $Y2=0
cc_133 B N_VPWR_M1007_d 0.00726586f $X=1.985 $Y=1.745 $X2=0 $Y2=0
cc_134 N_B_c_160_n N_VPWR_c_252_n 0.0144815f $X=1.525 $Y=1.99 $X2=0 $Y2=0
cc_135 B N_VPWR_c_252_n 0.0028364f $X=1.985 $Y=1.745 $X2=0 $Y2=0
cc_136 N_B_c_160_n N_VPWR_c_258_n 0.00742462f $X=1.525 $Y=1.99 $X2=0 $Y2=0
cc_137 N_B_c_160_n N_VPWR_c_259_n 0.00715641f $X=1.525 $Y=1.99 $X2=0 $Y2=0
cc_138 B N_VPWR_c_259_n 0.0429685f $X=1.985 $Y=1.745 $X2=0 $Y2=0
cc_139 N_B_c_160_n N_X_c_291_n 6.12275e-19 $X=1.525 $Y=1.99 $X2=0 $Y2=0
cc_140 B N_X_c_291_n 0.0265487f $X=1.985 $Y=1.745 $X2=0 $Y2=0
cc_141 N_B_M1001_g N_VGND_c_310_n 0.0197488f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_142 N_B_M1001_g N_VGND_c_311_n 0.00290915f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_143 N_B_M1001_g N_VGND_c_313_n 0.00534238f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A_225_413#_c_191_n N_VPWR_c_255_n 0.00482332f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_145 N_A_225_413#_M1002_d N_VPWR_c_252_n 0.0033624f $X=1.125 $Y=2.065 $X2=0
+ $Y2=0
cc_146 N_A_225_413#_c_191_n N_VPWR_c_252_n 0.00938119f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_147 N_A_225_413#_c_197_n N_VPWR_c_252_n 0.0122726f $X=1.28 $Y=2.225 $X2=0
+ $Y2=0
cc_148 N_A_225_413#_c_197_n N_VPWR_c_258_n 0.0158266f $X=1.28 $Y=2.225 $X2=0
+ $Y2=0
cc_149 N_A_225_413#_c_191_n N_VPWR_c_259_n 0.013221f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_150 N_A_225_413#_c_192_n X 0.00829818f $X=2.54 $Y=0.985 $X2=0 $Y2=0
cc_151 N_A_225_413#_c_191_n N_X_c_291_n 0.0342773f $X=2.515 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_225_413#_c_195_n N_X_c_291_n 0.00343613f $X=2.42 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_225_413#_c_191_n N_X_c_290_n 0.00637618f $X=2.515 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_225_413#_c_192_n N_X_c_290_n 0.0187814f $X=2.54 $Y=0.985 $X2=0 $Y2=0
cc_155 N_A_225_413#_c_195_n N_X_c_290_n 0.0225821f $X=2.42 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_225_413#_c_191_n N_VGND_c_310_n 9.07077e-19 $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_157 N_A_225_413#_c_192_n N_VGND_c_310_n 0.00356759f $X=2.54 $Y=0.985 $X2=0
+ $Y2=0
cc_158 N_A_225_413#_c_194_n N_VGND_c_310_n 0.0034384f $X=2.08 $Y=1.135 $X2=0
+ $Y2=0
cc_159 N_A_225_413#_c_195_n N_VGND_c_310_n 0.0161449f $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_160 N_A_225_413#_c_215_n N_VGND_c_310_n 0.00396157f $X=1.3 $Y=0.445 $X2=0
+ $Y2=0
cc_161 N_A_225_413#_c_215_n N_VGND_c_311_n 0.0177828f $X=1.3 $Y=0.445 $X2=0
+ $Y2=0
cc_162 N_A_225_413#_c_192_n N_VGND_c_312_n 0.00585385f $X=2.54 $Y=0.985 $X2=0
+ $Y2=0
cc_163 N_A_225_413#_M1003_s N_VGND_c_313_n 0.00284954f $X=1.175 $Y=0.235 $X2=0
+ $Y2=0
cc_164 N_A_225_413#_c_192_n N_VGND_c_313_n 0.0120647f $X=2.54 $Y=0.985 $X2=0
+ $Y2=0
cc_165 N_A_225_413#_c_215_n N_VGND_c_313_n 0.0145356f $X=1.3 $Y=0.445 $X2=0
+ $Y2=0
cc_166 N_VPWR_c_252_n N_X_M1005_d 0.00263275f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_167 N_VPWR_c_255_n N_X_c_291_n 0.0257166f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_168 N_VPWR_c_252_n N_X_c_291_n 0.0223143f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_169 N_VPWR_c_259_n N_X_c_291_n 0.017143f $X=2.275 $Y=2.485 $X2=0 $Y2=0
cc_170 X N_VGND_c_312_n 0.0263681f $X=2.875 $Y=0.425 $X2=0 $Y2=0
cc_171 N_X_M1004_d N_VGND_c_313_n 0.00558827f $X=2.615 $Y=0.235 $X2=0 $Y2=0
cc_172 X N_VGND_c_313_n 0.0143479f $X=2.875 $Y=0.425 $X2=0 $Y2=0
cc_173 N_VGND_c_313_n A_327_47# 0.0122415f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
