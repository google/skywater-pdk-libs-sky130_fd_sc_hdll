* NGSPICE file created from sky130_fd_sc_hdll__ebufn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__ebufn_4 A TE_B VGND VNB VPB VPWR Z
M1000 a_340_309# a_27_47# Z VPB phighvt w=1e+06u l=180000u
+  ad=1.9263e+12p pd=1.369e+07u as=5.8e+11p ps=5.16e+06u
M1001 Z a_27_47# a_413_47# VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=1.053e+12p ps=9.74e+06u
M1002 a_413_47# a_224_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.2475e+11p ps=6.13e+06u
M1003 a_413_47# a_27_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Z a_27_47# a_340_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_340_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=9.402e+11p ps=7.71e+06u
M1006 VGND a_224_47# a_413_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1008 VPWR TE_B a_340_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_224_47# TE_B VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1010 Z a_27_47# a_413_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_340_309# a_27_47# Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_340_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Z a_27_47# a_340_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_413_47# a_224_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_224_47# a_413_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR TE_B a_340_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_224_47# TE_B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1018 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1019 a_413_47# a_27_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

