* File: sky130_fd_sc_hdll__clkbuf_16.spice
* Created: Thu Aug 27 19:01:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkbuf_16.pex.spice"
.subckt sky130_fd_sc_hdll__clkbuf_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_A_118_297#_M1006_d N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.1323 PD=0.75 PS=1.47 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.2
+ SB=75009.3 A=0.063 P=1.14 MULT=1
MM1007 N_A_118_297#_M1006_d N_A_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75008.8 A=0.063 P=1.14 MULT=1
MM1011 N_A_118_297#_M1011_d N_A_M1011_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75008.3 A=0.063 P=1.14 MULT=1
MM1023 N_A_118_297#_M1011_d N_A_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0588 PD=0.75 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75007.9 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1023_s N_A_118_297#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0693 PD=0.7 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75007.4 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_118_297#_M1001_g N_X_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75007 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1001_d N_A_118_297#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.1
+ SB=75006.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_118_297#_M1005_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.5
+ SB=75006 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1005_d N_A_118_297#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75004
+ SB=75005.5 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_118_297#_M1017_g N_X_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75004.5
+ SB=75005 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1017_d N_A_118_297#_M1019_g N_X_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75005
+ SB=75004.6 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_118_297#_M1020_g N_X_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.0693 PD=0.745 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75005.5
+ SB=75004.1 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1020_d N_A_118_297#_M1021_g N_X_M1021_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.0693 PD=0.745 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75005.9
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_118_297#_M1024_g N_X_M1021_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75006.4
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1024_d N_A_118_297#_M1027_g N_X_M1027_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75006.9
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_A_118_297#_M1032_g N_X_M1027_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75007.4
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1032_d N_A_118_297#_M1033_g N_X_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75007.9
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_A_118_297#_M1036_g N_X_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75008.3
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1036_d N_A_118_297#_M1037_g N_X_M1037_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0798 PD=0.75 PS=0.8 NRD=0 NRS=14.28 M=1 R=2.8 SA=75008.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1039 N_VGND_M1039_d N_A_118_297#_M1039_g N_X_M1037_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0798 PD=1.37 PS=0.8 NRD=0 NRS=14.28 M=1 R=2.8 SA=75009.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_118_297#_M1013_d N_A_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90009.3 A=0.18 P=2.36 MULT=1
MM1014 N_A_118_297#_M1013_d N_A_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90008.8 A=0.18 P=2.36 MULT=1
MM1030 N_A_118_297#_M1030_d N_A_M1030_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90008.3 A=0.18 P=2.36 MULT=1
MM1034 N_A_118_297#_M1030_d N_A_M1034_g N_VPWR_M1034_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.6
+ SB=90007.9 A=0.18 P=2.36 MULT=1
MM1003 N_X_M1003_d N_A_118_297#_M1003_g N_VPWR_M1034_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.1
+ SB=90007.4 A=0.18 P=2.36 MULT=1
MM1004 N_X_M1003_d N_A_118_297#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.6
+ SB=90006.9 A=0.18 P=2.36 MULT=1
MM1008 N_X_M1008_d N_A_118_297#_M1008_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.1
+ SB=90006.4 A=0.18 P=2.36 MULT=1
MM1009 N_X_M1008_d N_A_118_297#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.5
+ SB=90005.9 A=0.18 P=2.36 MULT=1
MM1010 N_X_M1010_d N_A_118_297#_M1010_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90004
+ SB=90005.5 A=0.18 P=2.36 MULT=1
MM1015 N_X_M1010_d N_A_118_297#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90004.5
+ SB=90005 A=0.18 P=2.36 MULT=1
MM1016 N_X_M1016_d N_A_118_297#_M1016_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90005
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1018 N_X_M1016_d N_A_118_297#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.1475 PD=1.3 PS=1.295 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90005.5 SB=90004 A=0.18 P=2.36 MULT=1
MM1022 N_X_M1022_d N_A_118_297#_M1022_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.1475 PD=1.3 PS=1.295 NRD=1.9503 NRS=0.9653 M=1 R=5.55556
+ SA=90005.9 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1025 N_X_M1022_d N_A_118_297#_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90006.4
+ SB=90003.1 A=0.18 P=2.36 MULT=1
MM1026 N_X_M1026_d N_A_118_297#_M1026_g N_VPWR_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90006.9
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1028 N_X_M1026_d N_A_118_297#_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90007.4
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1029 N_X_M1029_d N_A_118_297#_M1029_g N_VPWR_M1028_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90007.9
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1031 N_X_M1029_d N_A_118_297#_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90008.3
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1035 N_X_M1035_d N_A_118_297#_M1035_g N_VPWR_M1031_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90008.8
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1038 N_X_M1035_d N_A_118_297#_M1038_g N_VPWR_M1038_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90009.3
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX40_noxref VNB VPB NWDIODE A=16.8525 P=24.21
*
.include "sky130_fd_sc_hdll__clkbuf_16.pxi.spice"
*
.ends
*
*
