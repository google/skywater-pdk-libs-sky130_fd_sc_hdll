* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand3b_4 A_N B C VGND VNB VPB VPWR Y
M1000 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.74e+12p pd=1.548e+07u as=2.61e+12p ps=2.322e+07u
M1001 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_225_47# B a_683_47# VNB nshort w=650000u l=150000u
+  ad=9.62e+11p pd=9.46e+06u as=8.645e+11p ps=7.86e+06u
M1004 a_683_47# B a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_225_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1006 Y a_27_47# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A_N a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1008 a_225_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C a_683_47# VNB nshort w=650000u l=150000u
+  ad=8.45e+11p pd=7.8e+06u as=0p ps=0u
M1012 a_683_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_225_47# B a_683_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y a_27_47# a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND C a_683_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_683_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1024 a_683_47# B a_225_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
