* File: sky130_fd_sc_hdll__inv_6.pex.spice
* Created: Thu Aug 27 19:09:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INV_6%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 38 39 40 61 64 68 72 76
c110 19 0 6.01499e-20 $X=1.905 $Y=1.41
r111 61 62 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=2.87 $Y2=1.202
r112 59 61 47.8071 $w=3.68e-07 $l=3.65e-07 $layer=POLY_cond $X=2.48 $Y=1.202
+ $X2=2.845 $Y2=1.202
r113 57 59 10.4783 $w=3.68e-07 $l=8e-08 $layer=POLY_cond $X=2.4 $Y=1.202
+ $X2=2.48 $Y2=1.202
r114 56 57 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.4 $Y2=1.202
r115 55 56 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=1.93 $Y=1.202
+ $X2=2.375 $Y2=1.202
r116 54 55 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r117 53 54 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.905 $Y2=1.202
r118 52 53 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r119 51 52 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.435 $Y2=1.202
r120 50 51 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r121 48 50 56.3207 $w=3.68e-07 $l=4.3e-07 $layer=POLY_cond $X=0.535 $Y=1.202
+ $X2=0.965 $Y2=1.202
r122 46 48 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.535 $Y2=1.202
r123 45 46 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r124 40 76 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=2.48 $Y=1.2
+ $X2=2.32 $Y2=1.2
r125 40 59 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.48
+ $Y=1.16 $X2=2.48 $Y2=1.16
r126 39 76 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=2.01 $Y=1.2
+ $X2=2.32 $Y2=1.2
r127 39 72 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.01 $Y=1.2
+ $X2=1.86 $Y2=1.2
r128 38 72 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=1.5 $Y=1.2 $X2=1.86
+ $Y2=1.2
r129 38 68 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=1.5 $Y=1.2 $X2=1.4
+ $Y2=1.2
r130 37 68 41.7184 $w=2.48e-07 $l=9.05e-07 $layer=LI1_cond $X=0.495 $Y=1.2
+ $X2=1.4 $Y2=1.2
r131 37 64 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.495 $Y=1.2
+ $X2=0.49 $Y2=1.2
r132 37 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.535
+ $Y=1.16 $X2=0.535 $Y2=1.16
r133 34 62 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=1.202
r134 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=0.56
r135 31 61 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r136 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r137 28 57 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.4 $Y2=1.202
r138 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.4 $Y2=0.56
r139 25 56 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r140 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r141 22 55 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r142 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r143 19 54 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r144 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r145 16 53 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r146 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r147 13 52 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r148 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r149 10 51 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r150 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r151 7 50 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r152 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r153 4 46 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r154 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r155 1 45 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r156 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_6%VPWR 1 2 3 4 13 15 19 23 25 29 33 36 37 38
+ 45 46 52 55
r57 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 43 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 43 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r64 40 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.14 $Y2=2.72
r65 40 42 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.99 $Y2=2.72
r66 38 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 38 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 36 42 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=3.08 $Y2=2.72
r70 35 45 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.45 $Y2=2.72
r71 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.08 $Y2=2.72
r72 31 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r73 31 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.34
r74 27 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r75 27 29 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r76 26 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72 $X2=1.2
+ $Y2=2.72
r77 25 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.14 $Y2=2.72
r78 25 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r79 21 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r80 21 23 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r81 20 49 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r82 19 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72 $X2=1.2
+ $Y2=2.72
r83 19 20 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r84 15 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r85 13 49 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.172 $Y2=2.72
r86 13 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r87 4 33 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2.34
r88 3 29 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r89 2 23 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r90 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r91 1 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_6%Y 1 2 3 4 5 6 19 21 25 27 28 29 33 37 39 45
+ 49 54 55 56 57 58 74 77 82
c108 82 0 6.01499e-20 $X=3.085 $Y=1.53
r109 64 70 28.0354 $w=1.78e-07 $l=4.55e-07 $layer=LI1_cond $X=3.065 $Y=0.815
+ $X2=2.61 $Y2=0.815
r110 58 82 0.291866 $w=1.88e-07 $l=5e-09 $layer=LI1_cond $X=3.08 $Y=1.59
+ $X2=3.085 $Y2=1.59
r111 58 65 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=3.08 $Y=1.59
+ $X2=3.065 $Y2=1.59
r112 58 65 0.720277 $w=3.98e-07 $l=2.5e-08 $layer=LI1_cond $X=3.065 $Y=1.47
+ $X2=3.065 $Y2=1.495
r113 57 58 8.0671 $w=3.98e-07 $l=2.8e-07 $layer=LI1_cond $X=3.065 $Y=1.19
+ $X2=3.065 $Y2=1.47
r114 56 74 0.308081 $w=1.78e-07 $l=5e-09 $layer=LI1_cond $X=3.08 $Y=0.815
+ $X2=3.085 $Y2=0.815
r115 56 64 0.924242 $w=1.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.08 $Y=0.815
+ $X2=3.065 $Y2=0.815
r116 56 57 7.77899 $w=3.98e-07 $l=2.7e-07 $layer=LI1_cond $X=3.065 $Y=0.92
+ $X2=3.065 $Y2=1.19
r117 56 64 0.432166 $w=3.98e-07 $l=1.5e-08 $layer=LI1_cond $X=3.065 $Y=0.92
+ $X2=3.065 $Y2=0.905
r118 47 70 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.61 $Y=0.725 $X2=2.61
+ $Y2=0.815
r119 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.61 $Y=0.725
+ $X2=2.61 $Y2=0.42
r120 43 65 28.0191 $w=1.88e-07 $l=4.8e-07 $layer=LI1_cond $X=2.585 $Y=1.59
+ $X2=3.065 $Y2=1.59
r121 43 77 11.2391 $w=1.88e-07 $l=1.9e-07 $layer=LI1_cond $X=2.585 $Y=1.59
+ $X2=2.395 $Y2=1.59
r122 43 45 19.8645 $w=3.78e-07 $l=6.55e-07 $layer=LI1_cond $X=2.585 $Y=1.685
+ $X2=2.585 $Y2=2.34
r123 42 54 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.645 $Y2=1.58
r124 42 77 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=2.395 $Y2=1.58
r125 40 55 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0.815
+ $X2=1.67 $Y2=0.815
r126 39 70 5.23737 $w=1.78e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0.815
+ $X2=2.61 $Y2=0.815
r127 39 40 47.4444 $w=1.78e-07 $l=7.7e-07 $layer=LI1_cond $X=2.525 $Y=0.815
+ $X2=1.755 $Y2=0.815
r128 35 55 1.54918 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.67 $Y=0.725 $X2=1.67
+ $Y2=0.815
r129 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.67 $Y=0.725
+ $X2=1.67 $Y2=0.42
r130 31 54 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=1.58
r131 31 33 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=2.34
r132 30 52 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.705 $Y2=1.58
r133 29 54 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=1.645 $Y2=1.58
r134 29 30 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=0.895 $Y2=1.58
r135 27 55 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0.815
+ $X2=1.67 $Y2=0.815
r136 27 28 47.4444 $w=1.78e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0.815
+ $X2=0.815 $Y2=0.815
r137 23 28 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.73 $Y=0.725
+ $X2=0.815 $Y2=0.815
r138 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=0.725
+ $X2=0.73 $Y2=0.42
r139 19 52 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.58
r140 19 21 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r141 6 43 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r142 6 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r143 5 54 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r144 5 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r145 4 52 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r146 4 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r147 3 49 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.42
r148 2 37 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.42
r149 1 25 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_6%VGND 1 2 3 4 13 15 17 21 23 27 31 33 35 42
+ 43 49 52 55 58
r58 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r59 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r60 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r61 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r62 43 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r63 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r64 40 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.015
+ $Y2=0
r65 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.45
+ $Y2=0
r66 39 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r67 39 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r68 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r69 36 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.14
+ $Y2=0
r70 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.53
+ $Y2=0
r71 35 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=3.015
+ $Y2=0
r72 35 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.53
+ $Y2=0
r73 33 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r74 33 58 0.0113817 $w=4.8e-07 $l=4e-08 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.19
+ $Y2=0
r75 33 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r76 29 55 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0
r77 29 31 11.5244 $w=2.98e-07 $l=3e-07 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0.385
r78 25 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r79 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.38
r80 24 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.2
+ $Y2=0
r81 23 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.14
+ $Y2=0
r82 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=1.285
+ $Y2=0
r83 19 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0
r84 19 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0.38
r85 18 46 4.1239 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r86 17 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.2
+ $Y2=0
r87 17 18 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.395
+ $Y2=0
r88 13 46 3.12417 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.262 $Y=0.085
+ $X2=0.197 $Y2=0
r89 13 15 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.262 $Y=0.085
+ $X2=0.262 $Y2=0.38
r90 4 31 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.385
r91 3 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r92 2 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r93 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends

