* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
M1000 a_357_297# B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=5.8e+11p ps=5.16e+06u
M1001 Y C2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1002 VGND C2 a_119_47# VNB nshort w=640000u l=150000u
+  ad=9.28e+11p pd=5.46e+06u as=1.344e+11p ps=1.7e+06u
M1003 Y B1 a_449_47# VNB nshort w=640000u l=150000u
+  ad=4.416e+11p pd=3.94e+06u as=1.344e+11p ps=1.7e+06u
M1004 a_117_297# B2 a_357_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_627_47# A1 Y VNB nshort w=640000u l=150000u
+  ad=2.432e+11p pd=2.04e+06u as=0p ps=0u
M1006 a_117_297# C1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_357_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.5e+11p ps=2.7e+06u
M1008 VGND A2 a_627_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_357_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_449_47# B2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_119_47# C1 Y VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
