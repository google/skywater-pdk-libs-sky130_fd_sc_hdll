* File: sky130_fd_sc_hdll__and2b_4.pex.spice
* Created: Wed Sep  2 08:22:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND2B_4%A_33_199# 1 2 7 9 10 12 14 15 16 19 26
r62 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.16 $X2=0.34 $Y2=1.16
r63 23 26 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.25 $Y=1.16 $X2=0.34
+ $Y2=1.16
r64 19 22 54.406 $w=2.13e-07 $l=1.015e-06 $layer=LI1_cond $X=3.832 $Y=0.68
+ $X2=3.832 $Y2=1.695
r65 17 22 11.7924 $w=2.13e-07 $l=2.2e-07 $layer=LI1_cond $X=3.832 $Y=1.915
+ $X2=3.832 $Y2=1.695
r66 15 17 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.725 $Y=2
+ $X2=3.832 $Y2=1.915
r67 15 16 221.166 $w=1.68e-07 $l=3.39e-06 $layer=LI1_cond $X=3.725 $Y=2
+ $X2=0.335 $Y2=2
r68 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.25 $Y=1.915
+ $X2=0.335 $Y2=2
r69 13 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.25 $Y=1.325
+ $X2=0.25 $Y2=1.16
r70 13 14 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.25 $Y=1.325
+ $X2=0.25 $Y2=1.915
r71 10 27 39.2524 $w=3.82e-07 $l=2.24332e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.38 $Y2=1.16
r72 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r73 7 27 45.1054 $w=3.82e-07 $l=3.02076e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.38 $Y2=1.16
r74 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r75 2 22 600 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_PDIFF $count=1 $X=3.62
+ $Y=1.485 $X2=3.815 $Y2=1.695
r76 1 19 182 $w=1.7e-07 $l=2.91419e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.465 $X2=3.81 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_4%B 1 3 4 6 7 11
r30 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r31 7 11 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=1.16 $X2=0.94
+ $Y2=1.16
r32 4 10 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.16
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r34 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.88 $Y=0.995
+ $X2=0.965 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.88 $Y=0.995 $X2=0.88
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_4%A_27_47# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 33 35 37 42 43 45 59
r114 59 60 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=2.975 $Y=1.202
+ $X2=3 $Y2=1.202
r115 58 59 61.062 $w=3.71e-07 $l=4.7e-07 $layer=POLY_cond $X=2.505 $Y=1.202
+ $X2=2.975 $Y2=1.202
r116 57 58 4.54717 $w=3.71e-07 $l=3.5e-08 $layer=POLY_cond $X=2.47 $Y=1.202
+ $X2=2.505 $Y2=1.202
r117 56 57 56.5148 $w=3.71e-07 $l=4.35e-07 $layer=POLY_cond $X=2.035 $Y=1.202
+ $X2=2.47 $Y2=1.202
r118 55 56 5.84636 $w=3.71e-07 $l=4.5e-08 $layer=POLY_cond $X=1.99 $Y=1.202
+ $X2=2.035 $Y2=1.202
r119 52 53 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=1.51 $Y=1.202
+ $X2=1.535 $Y2=1.202
r120 46 55 0.649596 $w=3.71e-07 $l=5e-09 $layer=POLY_cond $X=1.985 $Y=1.202
+ $X2=1.99 $Y2=1.202
r121 46 53 58.4636 $w=3.71e-07 $l=4.5e-07 $layer=POLY_cond $X=1.985 $Y=1.202
+ $X2=1.535 $Y2=1.202
r122 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.985
+ $Y=1.16 $X2=1.985 $Y2=1.16
r123 43 45 16.9665 $w=3.58e-07 $l=5.3e-07 $layer=LI1_cond $X=1.455 $Y=1.175
+ $X2=1.985 $Y2=1.175
r124 42 43 10.5932 $w=2.1e-07 $l=1.8e-07 $layer=LI1_cond $X=1.35 $Y=0.995
+ $X2=1.35 $Y2=1.175
r125 41 42 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=1.35 $Y=0.805
+ $X2=1.35 $Y2=0.995
r126 37 43 28.7021 $w=1.9e-07 $l=4.47e-07 $layer=LI1_cond $X=1.35 $Y=1.622
+ $X2=1.35 $Y2=1.175
r127 37 39 24.2248 $w=2.43e-07 $l=5.15e-07 $layer=LI1_cond $X=1.245 $Y=1.622
+ $X2=0.73 $Y2=1.622
r128 36 49 4.80081 $w=1.9e-07 $l=1.68e-07 $layer=LI1_cond $X=0.425 $Y=0.71
+ $X2=0.257 $Y2=0.71
r129 35 41 6.83868 $w=1.9e-07 $l=1.44914e-07 $layer=LI1_cond $X=1.245 $Y=0.71
+ $X2=1.35 $Y2=0.805
r130 35 36 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=1.245 $Y=0.71
+ $X2=0.425 $Y2=0.71
r131 31 49 2.71474 $w=3.35e-07 $l=9.5e-08 $layer=LI1_cond $X=0.257 $Y=0.615
+ $X2=0.257 $Y2=0.71
r132 31 33 8.0843 $w=3.33e-07 $l=2.35e-07 $layer=LI1_cond $X=0.257 $Y=0.615
+ $X2=0.257 $Y2=0.38
r133 28 60 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3 $Y=0.995 $X2=3
+ $Y2=1.202
r134 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3 $Y=0.995 $X2=3
+ $Y2=0.56
r135 25 59 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.975 $Y=1.41
+ $X2=2.975 $Y2=1.202
r136 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.975 $Y=1.41
+ $X2=2.975 $Y2=1.985
r137 22 58 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.505 $Y2=1.202
r138 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.505 $Y2=1.985
r139 19 57 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.47 $Y=0.995
+ $X2=2.47 $Y2=1.202
r140 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.47 $Y=0.995
+ $X2=2.47 $Y2=0.56
r141 16 56 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.035 $Y=1.41
+ $X2=2.035 $Y2=1.202
r142 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.035 $Y=1.41
+ $X2=2.035 $Y2=1.985
r143 13 55 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=1.202
r144 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=0.56
r145 10 53 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.202
r146 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.985
r147 7 52 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=1.202
r148 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.56
r149 2 39 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r150 1 49 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.72
r151 1 33 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_4%A_N 1 3 4 6 7
c30 4 0 1.30865e-19 $X=3.555 $Y=0.995
c31 1 0 1.71423e-19 $X=3.53 $Y=1.41
r32 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.16 $X2=3.42 $Y2=1.16
r33 4 10 38.5495 $w=3.2e-07 $l=2.08315e-07 $layer=POLY_cond $X=3.555 $Y=0.995
+ $X2=3.457 $Y2=1.16
r34 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.555 $Y=0.995
+ $X2=3.555 $Y2=0.675
r35 1 10 46.8073 $w=3.2e-07 $l=2.84165e-07 $layer=POLY_cond $X=3.53 $Y=1.41
+ $X2=3.457 $Y2=1.16
r36 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.53 $Y=1.41 $X2=3.53
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_4%VPWR 1 2 3 4 13 15 17 21 23 26 29 32 39 40
+ 46 49
r59 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 49 52 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.245 $Y=2.36
+ $X2=2.245 $Y2=2.72
r61 47 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r64 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 37 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 34 52 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.435 $Y=2.72
+ $X2=2.245 $Y2=2.72
r68 34 36 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.435 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 32 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 32 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 30 39 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.375 $Y=2.72
+ $X2=3.91 $Y2=2.72
r72 29 36 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=2.99 $Y2=2.72
r73 28 30 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.185 $Y=2.72
+ $X2=3.375 $Y2=2.72
r74 28 29 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.185 $Y=2.72
+ $X2=2.995 $Y2=2.72
r75 26 28 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.185 $Y=2.36
+ $X2=3.185 $Y2=2.72
r76 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=2.72
+ $X2=1.255 $Y2=2.72
r77 23 52 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.245 $Y2=2.72
r78 23 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.42 $Y2=2.72
r79 19 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=2.635
+ $X2=1.255 $Y2=2.72
r80 19 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.255 $Y=2.635
+ $X2=1.255 $Y2=2.36
r81 18 43 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r82 17 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=2.72
+ $X2=1.255 $Y2=2.72
r83 17 18 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.09 $Y=2.72
+ $X2=0.425 $Y2=2.72
r84 13 43 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r85 13 15 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2.34
r86 4 26 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.21 $Y2=2.36
r87 3 49 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=1.485 $X2=2.27 $Y2=2.36
r88 2 21 600 $w=1.7e-07 $l=9.69858e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.255 $Y2=2.36
r89 1 15 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_4%X 1 2 3 4 13 18 23 26 30 32
c47 32 0 1.30865e-19 $X=2.53 $Y=0.85
c48 23 0 1.71423e-19 $X=2.712 $Y=1.535
r49 30 32 0.558915 $w=5.33e-07 $l=2.5e-08 $layer=LI1_cond $X=2.712 $Y=0.825
+ $X2=2.712 $Y2=0.85
r50 26 30 2.44399 $w=5.35e-07 $l=1.05e-07 $layer=LI1_cond $X=2.712 $Y=0.72
+ $X2=2.712 $Y2=0.825
r51 26 32 0.670698 $w=5.33e-07 $l=3e-08 $layer=LI1_cond $X=2.712 $Y=0.88
+ $X2=2.712 $Y2=0.85
r52 23 26 14.6436 $w=5.33e-07 $l=6.55e-07 $layer=LI1_cond $X=2.712 $Y=1.535
+ $X2=2.712 $Y2=0.88
r53 23 25 2.44399 $w=5.35e-07 $l=1.05e-07 $layer=LI1_cond $X=2.712 $Y=1.535
+ $X2=2.712 $Y2=1.64
r54 21 26 25.356 $w=2.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.865 $Y=0.72
+ $X2=2.445 $Y2=0.72
r55 20 21 0.0965754 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=1.77 $Y=0.72
+ $X2=1.865 $Y2=0.72
r56 18 20 3.50239 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=1.77 $Y=0.66 $X2=1.77
+ $Y2=0.72
r57 13 25 6.21471 $w=2.1e-07 $l=2.67e-07 $layer=LI1_cond $X=2.445 $Y=1.64
+ $X2=2.712 $Y2=1.64
r58 13 15 34.0649 $w=2.08e-07 $l=6.45e-07 $layer=LI1_cond $X=2.445 $Y=1.64
+ $X2=1.8 $Y2=1.64
r59 4 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.595
+ $Y=1.485 $X2=2.74 $Y2=1.62
r60 3 15 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.625
+ $Y=1.485 $X2=1.8 $Y2=1.62
r61 2 26 182 $w=1.7e-07 $l=5.92431e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.235 $X2=2.735 $Y2=0.74
r62 1 18 182 $w=1.7e-07 $l=5.09166e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.77 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_4%VGND 1 2 3 12 14 16 17 23 25 35 36 39 43
r60 43 46 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.225
+ $Y2=0.36
r61 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r62 40 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r63 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r64 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r65 33 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r66 33 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r67 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r68 30 43 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.225
+ $Y2=0
r69 30 32 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.99
+ $Y2=0
r70 28 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r71 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r72 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r73 25 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.69
+ $Y2=0
r74 23 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r75 19 35 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.91
+ $Y2=0
r76 17 32 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=0 $X2=2.99
+ $Y2=0
r77 16 21 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.185
+ $Y2=0.36
r78 16 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.375
+ $Y2=0
r79 16 17 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=2.995
+ $Y2=0
r80 15 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r81 14 43 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.225
+ $Y2=0
r82 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.385
+ $Y2=0
r83 10 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r84 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.36
r85 3 21 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.235 $X2=3.21 $Y2=0.36
r86 2 46 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.235 $X2=2.25 $Y2=0.36
r87 1 12 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=0.955
+ $Y=0.235 $X2=1.22 $Y2=0.36
.ends

