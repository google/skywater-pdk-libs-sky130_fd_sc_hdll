* File: sky130_fd_sc_hdll__nor3_4.pxi.spice
* Created: Wed Sep  2 08:40:28 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR3_4%A N_A_c_92_n N_A_M1004_g N_A_c_98_n N_A_M1003_g
+ N_A_c_93_n N_A_M1013_g N_A_c_99_n N_A_M1009_g N_A_c_94_n N_A_M1014_g
+ N_A_c_100_n N_A_M1012_g N_A_c_101_n N_A_M1016_g N_A_c_95_n N_A_M1020_g A
+ N_A_c_96_n N_A_c_97_n PM_SKY130_FD_SC_HDLL__NOR3_4%A
x_PM_SKY130_FD_SC_HDLL__NOR3_4%B N_B_c_164_n N_B_M1005_g N_B_c_172_n N_B_M1001_g
+ N_B_c_165_n N_B_M1007_g N_B_c_173_n N_B_M1018_g N_B_c_174_n N_B_M1019_g
+ N_B_c_166_n N_B_M1011_g N_B_c_167_n N_B_M1022_g N_B_c_168_n N_B_M1017_g
+ N_B_c_176_n N_B_c_177_n N_B_c_178_n N_B_c_179_n N_B_c_169_n N_B_c_170_n B
+ N_B_c_171_n B PM_SKY130_FD_SC_HDLL__NOR3_4%B
x_PM_SKY130_FD_SC_HDLL__NOR3_4%C N_C_c_290_n N_C_M1000_g N_C_c_295_n N_C_M1006_g
+ N_C_c_291_n N_C_M1002_g N_C_c_296_n N_C_M1010_g N_C_c_292_n N_C_M1008_g
+ N_C_c_297_n N_C_M1015_g N_C_c_298_n N_C_M1021_g N_C_c_293_n N_C_M1023_g C
+ N_C_c_311_n N_C_c_294_n PM_SKY130_FD_SC_HDLL__NOR3_4%C
x_PM_SKY130_FD_SC_HDLL__NOR3_4%A_27_297# N_A_27_297#_M1003_s N_A_27_297#_M1009_s
+ N_A_27_297#_M1016_s N_A_27_297#_M1018_s N_A_27_297#_M1022_s
+ N_A_27_297#_c_379_n N_A_27_297#_c_427_p N_A_27_297#_c_380_n
+ N_A_27_297#_c_413_p N_A_27_297#_c_381_n N_A_27_297#_c_382_n
+ N_A_27_297#_c_415_p N_A_27_297#_c_416_p N_A_27_297#_c_443_p
+ N_A_27_297#_c_383_n N_A_27_297#_c_396_n N_A_27_297#_c_398_n
+ N_A_27_297#_c_400_n N_A_27_297#_c_420_p N_A_27_297#_c_401_n
+ PM_SKY130_FD_SC_HDLL__NOR3_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR3_4%VPWR N_VPWR_M1003_d N_VPWR_M1012_d N_VPWR_c_472_n
+ N_VPWR_c_473_n N_VPWR_c_474_n VPWR N_VPWR_c_475_n N_VPWR_c_471_n
+ N_VPWR_c_477_n N_VPWR_c_478_n VPWR PM_SKY130_FD_SC_HDLL__NOR3_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR3_4%A_497_297# N_A_497_297#_M1001_d
+ N_A_497_297#_M1019_d N_A_497_297#_M1010_s N_A_497_297#_M1021_s
+ N_A_497_297#_c_551_n N_A_497_297#_c_552_n N_A_497_297#_c_580_n
+ N_A_497_297#_c_566_n N_A_497_297#_c_568_n N_A_497_297#_c_553_n
+ N_A_497_297#_c_588_n N_A_497_297#_c_589_n
+ PM_SKY130_FD_SC_HDLL__NOR3_4%A_497_297#
x_PM_SKY130_FD_SC_HDLL__NOR3_4%Y N_Y_M1004_s N_Y_M1014_s N_Y_M1005_d N_Y_M1011_d
+ N_Y_M1002_d N_Y_M1023_d N_Y_M1006_d N_Y_M1015_d N_Y_c_632_n N_Y_c_617_n
+ N_Y_c_618_n N_Y_c_643_n N_Y_c_619_n N_Y_c_647_n N_Y_c_620_n N_Y_c_663_n
+ N_Y_c_621_n N_Y_c_667_n N_Y_c_699_n N_Y_c_622_n N_Y_c_630_n N_Y_c_708_n
+ N_Y_c_623_n N_Y_c_624_n N_Y_c_625_n N_Y_c_626_n N_Y_c_680_n N_Y_c_627_n
+ N_Y_c_682_n N_Y_c_628_n Y PM_SKY130_FD_SC_HDLL__NOR3_4%Y
x_PM_SKY130_FD_SC_HDLL__NOR3_4%VGND N_VGND_M1004_d N_VGND_M1013_d N_VGND_M1020_d
+ N_VGND_M1007_s N_VGND_M1000_s N_VGND_M1008_s N_VGND_M1017_s N_VGND_c_799_n
+ N_VGND_c_800_n N_VGND_c_801_n N_VGND_c_802_n N_VGND_c_803_n N_VGND_c_804_n
+ N_VGND_c_805_n N_VGND_c_806_n N_VGND_c_807_n N_VGND_c_808_n N_VGND_c_809_n
+ N_VGND_c_810_n N_VGND_c_811_n N_VGND_c_812_n N_VGND_c_813_n N_VGND_c_814_n
+ N_VGND_c_815_n N_VGND_c_816_n N_VGND_c_817_n VGND N_VGND_c_818_n
+ N_VGND_c_819_n N_VGND_c_820_n PM_SKY130_FD_SC_HDLL__NOR3_4%VGND
cc_1 VNB N_A_c_92_n 0.0218461f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_93_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_3 VNB N_A_c_94_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_4 VNB N_A_c_95_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_5 VNB N_A_c_96_n 0.0200187f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_6 VNB N_A_c_97_n 0.0801694f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_7 VNB N_B_c_164_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_B_c_165_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_9 VNB N_B_c_166_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_10 VNB N_B_c_167_n 0.0295f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_11 VNB N_B_c_168_n 0.0200445f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_12 VNB N_B_c_169_n 0.00679719f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_13 VNB N_B_c_170_n 0.00146858f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.202
cc_14 VNB N_B_c_171_n 0.0545376f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_C_c_290_n 0.0164927f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_16 VNB N_C_c_291_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_17 VNB N_C_c_292_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_18 VNB N_C_c_293_n 0.0173889f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_19 VNB N_C_c_294_n 0.0741172f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.202
cc_20 VNB N_VPWR_c_471_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_21 VNB N_Y_c_617_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.202
cc_22 VNB N_Y_c_618_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_23 VNB N_Y_c_619_n 0.00447396f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.202
cc_24 VNB N_Y_c_620_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.18
cc_25 VNB N_Y_c_621_n 0.0030003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_622_n 0.00275958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_623_n 0.019284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_624_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_625_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_626_n 0.00253348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_627_n 0.00251836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_628_n 0.00397012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB Y 0.0219404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_799_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_35 VNB N_VGND_c_800_n 0.0334656f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_36 VNB N_VGND_c_801_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_802_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_38 VNB N_VGND_c_803_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=1.202
cc_39 VNB N_VGND_c_804_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_40 VNB N_VGND_c_805_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_806_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_807_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_808_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_809_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_810_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_811_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_812_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_813_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_814_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_815_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_816_n 0.0192745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_817_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_818_n 0.014725f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_819_n 0.31689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_820_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VPB N_A_c_98_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_57 VPB N_A_c_99_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_58 VPB N_A_c_100_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_59 VPB N_A_c_101_n 0.0161064f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_60 VPB N_A_c_97_n 0.048391f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_61 VPB N_B_c_172_n 0.0164231f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_62 VPB N_B_c_173_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_63 VPB N_B_c_174_n 0.0161042f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.995
cc_64 VPB N_B_c_167_n 0.0315461f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_65 VPB N_B_c_176_n 0.0021681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_B_c_177_n 0.0077831f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_67 VPB N_B_c_178_n 2.85754e-19 $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_68 VPB N_B_c_179_n 0.00119741f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_69 VPB N_B_c_171_n 0.0328562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_C_c_295_n 0.0164077f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_71 VPB N_C_c_296_n 0.0158625f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_72 VPB N_C_c_297_n 0.0158724f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_73 VPB N_C_c_298_n 0.0159787f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_74 VPB N_C_c_294_n 0.0465936f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.202
cc_75 VPB N_A_27_297#_c_379_n 0.00371848f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_76 VPB N_A_27_297#_c_380_n 0.00196267f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_77 VPB N_A_27_297#_c_381_n 0.00201678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_297#_c_382_n 0.00416269f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_79 VPB N_A_27_297#_c_383_n 0.00151002f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_80 VPB N_VPWR_c_472_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_81 VPB N_VPWR_c_473_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.995
cc_82 VPB N_VPWR_c_474_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_83 VPB N_VPWR_c_475_n 0.114889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_471_n 0.0496483f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_85 VPB N_VPWR_c_477_n 0.0244347f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_86 VPB N_VPWR_c_478_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_87 VPB N_A_497_297#_c_551_n 0.00196267f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_88 VPB N_A_497_297#_c_552_n 0.0026013f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_89 VPB N_A_497_297#_c_553_n 0.00173525f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_90 VPB N_Y_c_630_n 0.014771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB Y 0.0270229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 N_A_c_95_n N_B_c_164_n 0.0243397f $X=1.95 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_93 N_A_c_101_n N_B_c_172_n 0.00971598f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_c_96_n N_B_c_169_n 0.0121231f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_c_97_n N_B_c_169_n 2.62535e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_96 N_A_c_96_n N_B_c_171_n 2.62535e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_c_97_n N_B_c_171_n 0.0243397f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_98 N_A_c_96_n N_A_27_297#_c_379_n 0.021852f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_c_98_n N_A_27_297#_c_380_n 0.0158351f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_c_99_n N_A_27_297#_c_380_n 0.0156273f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_96_n N_A_27_297#_c_380_n 0.0487385f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_c_97_n N_A_27_297#_c_380_n 0.00837544f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_103 N_A_c_100_n N_A_27_297#_c_381_n 0.0156273f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_c_101_n N_A_27_297#_c_381_n 0.0155666f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_c_96_n N_A_27_297#_c_381_n 0.0480109f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_c_97_n N_A_27_297#_c_381_n 0.00816971f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_107 N_A_c_96_n N_A_27_297#_c_383_n 0.0204509f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_c_97_n N_A_27_297#_c_383_n 0.00656533f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_109 N_A_c_98_n N_VPWR_c_472_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_c_99_n N_VPWR_c_472_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_99_n N_VPWR_c_473_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_c_100_n N_VPWR_c_473_n 0.00702461f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_c_100_n N_VPWR_c_474_n 0.00300743f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_c_101_n N_VPWR_c_474_n 0.00300743f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_c_101_n N_VPWR_c_475_n 0.00702461f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_c_98_n N_VPWR_c_471_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_c_99_n N_VPWR_c_471_n 0.0124092f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_c_100_n N_VPWR_c_471_n 0.0124092f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_101_n N_VPWR_c_471_n 0.0124344f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_98_n N_VPWR_c_477_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_c_92_n N_Y_c_632_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_c_93_n N_Y_c_632_n 0.00686626f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_c_94_n N_Y_c_632_n 5.45498e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_c_93_n N_Y_c_617_n 0.00901745f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_94_n N_Y_c_617_n 0.00901745f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_96_n N_Y_c_617_n 0.0398926f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_c_97_n N_Y_c_617_n 0.00345541f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_128 N_A_c_92_n N_Y_c_618_n 0.00266157f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_c_93_n N_Y_c_618_n 0.00116636f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_96_n N_Y_c_618_n 0.0307014f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_c_97_n N_Y_c_618_n 0.00358305f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_132 N_A_c_93_n N_Y_c_643_n 5.24597e-19 $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_94_n N_Y_c_643_n 0.00651696f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_95_n N_Y_c_619_n 0.0106151f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_96_n N_Y_c_619_n 0.0118017f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_95_n N_Y_c_647_n 5.32212e-19 $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_94_n N_Y_c_624_n 0.00119564f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_c_96_n N_Y_c_624_n 0.030835f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_c_97_n N_Y_c_624_n 0.00486271f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_140 N_A_c_92_n N_VGND_c_800_n 0.00496762f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_c_96_n N_VGND_c_800_n 0.0233945f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_c_92_n N_VGND_c_801_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_c_93_n N_VGND_c_801_n 0.00423334f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_c_93_n N_VGND_c_802_n 0.00379224f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_94_n N_VGND_c_802_n 0.00276126f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_95_n N_VGND_c_803_n 0.00268723f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_94_n N_VGND_c_808_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_c_95_n N_VGND_c_808_n 0.00437852f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_c_92_n N_VGND_c_819_n 0.0106014f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_c_93_n N_VGND_c_819_n 0.006093f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_c_94_n N_VGND_c_819_n 0.00608558f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_c_95_n N_VGND_c_819_n 0.00615622f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B_c_166_n N_C_c_290_n 0.0172799f $X=3.36 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_154 N_B_c_174_n N_C_c_295_n 0.00950644f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B_c_176_n N_C_c_295_n 8.60137e-19 $X=4 $Y=1.445 $X2=0 $Y2=0
cc_156 N_B_c_178_n N_C_c_295_n 0.00126614f $X=4.085 $Y=1.53 $X2=0 $Y2=0
cc_157 N_B_c_176_n N_C_c_296_n 7.76481e-19 $X=4 $Y=1.445 $X2=0 $Y2=0
cc_158 N_B_c_177_n N_C_c_296_n 0.0123908f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_159 N_B_c_177_n N_C_c_297_n 0.0118911f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_160 N_B_c_167_n N_C_c_298_n 0.0377754f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_161 N_B_c_177_n N_C_c_298_n 0.011848f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_162 N_B_c_179_n N_C_c_298_n 6.53633e-19 $X=5.63 $Y=1.445 $X2=0 $Y2=0
cc_163 N_B_c_168_n N_C_c_293_n 0.0104094f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B_c_167_n N_C_c_311_n 2.50769e-19 $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B_c_177_n N_C_c_311_n 0.0752208f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_166 N_B_c_169_n N_C_c_311_n 0.0168497f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_167 N_B_c_170_n N_C_c_311_n 0.0124922f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B_c_167_n N_C_c_294_n 0.0248037f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B_c_176_n N_C_c_294_n 0.0104489f $X=4 $Y=1.445 $X2=0 $Y2=0
cc_170 N_B_c_177_n N_C_c_294_n 0.0185005f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_171 N_B_c_179_n N_C_c_294_n 0.00195024f $X=5.63 $Y=1.445 $X2=0 $Y2=0
cc_172 N_B_c_169_n N_C_c_294_n 0.0268928f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_173 N_B_c_170_n N_C_c_294_n 9.05613e-19 $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B_c_171_n N_C_c_294_n 0.0172799f $X=3.335 $Y=1.202 $X2=0 $Y2=0
cc_175 N_B_c_172_n N_A_27_297#_c_382_n 2.98195e-19 $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_176 N_B_c_172_n N_A_27_297#_c_396_n 0.0212527f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_177 N_B_c_173_n N_A_27_297#_c_396_n 0.0155785f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_178 N_B_c_172_n N_A_27_297#_c_398_n 3.44206e-19 $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B_c_173_n N_A_27_297#_c_398_n 0.0023925f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B_c_167_n N_A_27_297#_c_400_n 0.00315098f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_181 N_B_c_174_n N_A_27_297#_c_401_n 0.00378027f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B_c_167_n N_A_27_297#_c_401_n 0.00170122f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B_c_177_n N_A_27_297#_c_401_n 0.00147363f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_184 N_B_c_178_n N_A_27_297#_c_401_n 3.67354e-19 $X=4.085 $Y=1.53 $X2=0 $Y2=0
cc_185 N_B_c_172_n N_VPWR_c_475_n 0.00429453f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B_c_173_n N_VPWR_c_475_n 0.00429453f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_187 N_B_c_174_n N_VPWR_c_475_n 0.00702461f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B_c_167_n N_VPWR_c_475_n 0.00702461f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_189 N_B_c_172_n N_VPWR_c_471_n 0.00609021f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_190 N_B_c_173_n N_VPWR_c_471_n 0.00536044f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B_c_174_n N_VPWR_c_471_n 0.00625464f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B_c_167_n N_VPWR_c_471_n 0.00686589f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B_c_177_n N_A_497_297#_M1010_s 0.00183837f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_194 N_B_c_177_n N_A_497_297#_M1021_s 0.00183837f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_195 N_B_c_173_n N_A_497_297#_c_551_n 0.0117691f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B_c_174_n N_A_497_297#_c_551_n 0.0116631f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B_c_169_n N_A_497_297#_c_551_n 0.0487385f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_198 N_B_c_171_n N_A_497_297#_c_551_n 0.00816971f $X=3.335 $Y=1.202 $X2=0
+ $Y2=0
cc_199 N_B_c_178_n N_A_497_297#_c_552_n 0.00226124f $X=4.085 $Y=1.53 $X2=0 $Y2=0
cc_200 N_B_c_169_n N_A_497_297#_c_552_n 0.0214236f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_201 N_B_c_172_n N_A_497_297#_c_553_n 2.98195e-19 $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_169_n N_A_497_297#_c_553_n 0.0197909f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_203 N_B_c_171_n N_A_497_297#_c_553_n 0.00648575f $X=3.335 $Y=1.202 $X2=0
+ $Y2=0
cc_204 N_B_c_177_n N_Y_M1006_d 4.37662e-19 $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_205 N_B_c_178_n N_Y_M1006_d 0.0017553f $X=4.085 $Y=1.53 $X2=0 $Y2=0
cc_206 N_B_c_177_n N_Y_M1015_d 0.00183401f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_207 N_B_c_164_n N_Y_c_619_n 0.00865686f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_208 N_B_c_169_n N_Y_c_619_n 0.00826974f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_209 N_B_c_164_n N_Y_c_647_n 0.00644736f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B_c_165_n N_Y_c_647_n 0.00693563f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B_c_166_n N_Y_c_647_n 5.34196e-19 $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B_c_165_n N_Y_c_620_n 0.00929182f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B_c_166_n N_Y_c_620_n 0.00650032f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B_c_169_n N_Y_c_620_n 0.0400808f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_215 N_B_c_171_n N_Y_c_620_n 0.00468948f $X=3.335 $Y=1.202 $X2=0 $Y2=0
cc_216 N_B_c_165_n N_Y_c_663_n 5.69266e-19 $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B_c_166_n N_Y_c_663_n 0.00857123f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B_c_177_n N_Y_c_621_n 0.00519546f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_219 N_B_c_169_n N_Y_c_621_n 0.0260084f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_220 N_B_c_177_n N_Y_c_667_n 0.0360776f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_221 N_B_c_167_n N_Y_c_630_n 0.01732f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_222 N_B_c_177_n N_Y_c_630_n 0.0324187f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_223 N_B_c_170_n N_Y_c_630_n 0.00420776f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_224 N_B_c_167_n N_Y_c_623_n 0.00469442f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B_c_168_n N_Y_c_623_n 0.0126624f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B_c_170_n N_Y_c_623_n 0.0190977f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_227 N_B_c_164_n N_Y_c_625_n 0.00116636f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B_c_165_n N_Y_c_625_n 0.00116636f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B_c_169_n N_Y_c_625_n 0.0307014f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_230 N_B_c_171_n N_Y_c_625_n 0.00358305f $X=3.335 $Y=1.202 $X2=0 $Y2=0
cc_231 N_B_c_166_n N_Y_c_626_n 0.00269873f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B_c_169_n N_Y_c_626_n 0.0315242f $X=3.915 $Y=1.18 $X2=0 $Y2=0
cc_233 N_B_c_177_n N_Y_c_680_n 0.00317598f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_234 N_B_c_178_n N_Y_c_680_n 0.0108404f $X=4.085 $Y=1.53 $X2=0 $Y2=0
cc_235 N_B_c_177_n N_Y_c_682_n 0.0131392f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_236 N_B_c_167_n N_Y_c_628_n 0.00188952f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B_c_177_n N_Y_c_628_n 0.00867931f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_238 N_B_c_170_n N_Y_c_628_n 0.0057042f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_239 N_B_c_167_n Y 0.020908f $X=5.685 $Y=1.41 $X2=0 $Y2=0
cc_240 N_B_c_168_n Y 0.00291891f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B_c_177_n Y 0.00839911f $X=5.545 $Y=1.53 $X2=0 $Y2=0
cc_242 N_B_c_179_n Y 0.00710913f $X=5.63 $Y=1.445 $X2=0 $Y2=0
cc_243 N_B_c_170_n Y 0.016408f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_244 N_B_c_164_n N_VGND_c_803_n 0.00268723f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_245 N_B_c_165_n N_VGND_c_804_n 0.00385467f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_246 N_B_c_166_n N_VGND_c_804_n 0.00365402f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_247 N_B_c_168_n N_VGND_c_807_n 0.00438629f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B_c_164_n N_VGND_c_810_n 0.00423334f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B_c_165_n N_VGND_c_810_n 0.00423334f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B_c_166_n N_VGND_c_812_n 0.00396605f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B_c_168_n N_VGND_c_816_n 0.00437852f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B_c_164_n N_VGND_c_819_n 0.00587047f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_253 N_B_c_165_n N_VGND_c_819_n 0.00620835f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_254 N_B_c_166_n N_VGND_c_819_n 0.00583042f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_255 N_B_c_168_n N_VGND_c_819_n 0.00715937f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_256 N_C_c_298_n N_A_27_297#_c_400_n 2.84537e-19 $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_257 N_C_c_295_n N_A_27_297#_c_401_n 0.0097459f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_258 N_C_c_296_n N_A_27_297#_c_401_n 0.00403222f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_259 N_C_c_297_n N_A_27_297#_c_401_n 0.00403222f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_260 N_C_c_298_n N_A_27_297#_c_401_n 0.00404951f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_261 N_C_c_295_n N_VPWR_c_475_n 0.00429453f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_262 N_C_c_296_n N_VPWR_c_475_n 0.00429453f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_263 N_C_c_297_n N_VPWR_c_475_n 0.00429453f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_264 N_C_c_298_n N_VPWR_c_475_n 0.00429453f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_265 N_C_c_295_n N_VPWR_c_471_n 0.00549531f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_266 N_C_c_296_n N_VPWR_c_471_n 0.0054701f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_267 N_C_c_297_n N_VPWR_c_471_n 0.0054701f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_268 N_C_c_298_n N_VPWR_c_471_n 0.00549531f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_269 N_C_c_295_n N_A_497_297#_c_552_n 2.98195e-19 $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_270 N_C_c_295_n N_A_497_297#_c_566_n 0.0089518f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_271 N_C_c_296_n N_A_497_297#_c_566_n 0.00966052f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_272 N_C_c_297_n N_A_497_297#_c_568_n 0.00961745f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_273 N_C_c_298_n N_A_497_297#_c_568_n 0.00966501f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_274 N_C_c_290_n N_Y_c_663_n 0.00686626f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_275 N_C_c_291_n N_Y_c_663_n 5.45498e-19 $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_276 N_C_c_290_n N_Y_c_621_n 0.00901745f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_277 N_C_c_291_n N_Y_c_621_n 0.00997702f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_278 N_C_c_311_n N_Y_c_621_n 0.00266908f $X=5.04 $Y=1.16 $X2=0 $Y2=0
cc_279 N_C_c_294_n N_Y_c_621_n 0.00345343f $X=5.215 $Y=1.202 $X2=0 $Y2=0
cc_280 N_C_c_296_n N_Y_c_667_n 0.0109083f $X=4.275 $Y=1.41 $X2=0 $Y2=0
cc_281 N_C_c_297_n N_Y_c_667_n 0.0109083f $X=4.745 $Y=1.41 $X2=0 $Y2=0
cc_282 N_C_c_290_n N_Y_c_699_n 5.24597e-19 $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_283 N_C_c_291_n N_Y_c_699_n 0.00651696f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_284 N_C_c_292_n N_Y_c_699_n 0.00693563f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_285 N_C_c_293_n N_Y_c_699_n 5.34196e-19 $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_286 N_C_c_292_n N_Y_c_622_n 0.00928691f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_287 N_C_c_293_n N_Y_c_622_n 0.00649747f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_288 N_C_c_311_n N_Y_c_622_n 0.040146f $X=5.04 $Y=1.16 $X2=0 $Y2=0
cc_289 N_C_c_294_n N_Y_c_622_n 0.0046868f $X=5.215 $Y=1.202 $X2=0 $Y2=0
cc_290 N_C_c_298_n N_Y_c_630_n 0.0106623f $X=5.215 $Y=1.41 $X2=0 $Y2=0
cc_291 N_C_c_292_n N_Y_c_708_n 5.69266e-19 $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_292 N_C_c_293_n N_Y_c_708_n 0.00857123f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_293 N_C_c_290_n N_Y_c_626_n 0.00112787f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_294 N_C_c_294_n N_Y_c_680_n 6.87638e-19 $X=5.215 $Y=1.202 $X2=0 $Y2=0
cc_295 N_C_c_291_n N_Y_c_627_n 0.00116508f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_296 N_C_c_292_n N_Y_c_627_n 0.00116508f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_297 N_C_c_311_n N_Y_c_627_n 0.0307598f $X=5.04 $Y=1.16 $X2=0 $Y2=0
cc_298 N_C_c_294_n N_Y_c_627_n 0.00358038f $X=5.215 $Y=1.202 $X2=0 $Y2=0
cc_299 N_C_c_293_n N_Y_c_628_n 0.0027131f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_300 N_C_c_311_n N_Y_c_628_n 0.00609668f $X=5.04 $Y=1.16 $X2=0 $Y2=0
cc_301 N_C_c_290_n N_VGND_c_805_n 0.00379224f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_302 N_C_c_291_n N_VGND_c_805_n 0.00276126f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_303 N_C_c_292_n N_VGND_c_806_n 0.00385467f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_304 N_C_c_293_n N_VGND_c_806_n 0.00365402f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_305 N_C_c_290_n N_VGND_c_812_n 0.00423334f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_306 N_C_c_291_n N_VGND_c_814_n 0.00423334f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_307 N_C_c_292_n N_VGND_c_814_n 0.00423334f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_308 N_C_c_293_n N_VGND_c_816_n 0.00396605f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_309 N_C_c_290_n N_VGND_c_819_n 0.00599324f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_310 N_C_c_291_n N_VGND_c_819_n 0.00597024f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_311 N_C_c_292_n N_VGND_c_819_n 0.00620835f $X=4.72 $Y=0.995 $X2=0 $Y2=0
cc_312 N_C_c_293_n N_VGND_c_819_n 0.00594864f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A_27_297#_c_380_n N_VPWR_M1003_d 0.00187091f $X=1.095 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_314 N_A_27_297#_c_381_n N_VPWR_M1012_d 0.00187091f $X=2.035 $Y=1.54 $X2=0
+ $Y2=0
cc_315 N_A_27_297#_c_380_n N_VPWR_c_472_n 0.0143191f $X=1.095 $Y=1.54 $X2=0
+ $Y2=0
cc_316 N_A_27_297#_c_413_p N_VPWR_c_473_n 0.0149311f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_317 N_A_27_297#_c_381_n N_VPWR_c_474_n 0.0143191f $X=2.035 $Y=1.54 $X2=0
+ $Y2=0
cc_318 N_A_27_297#_c_415_p N_VPWR_c_475_n 0.015002f $X=2.16 $Y=2.085 $X2=0 $Y2=0
cc_319 N_A_27_297#_c_416_p N_VPWR_c_475_n 0.0149886f $X=3.1 $Y=2.085 $X2=0 $Y2=0
cc_320 N_A_27_297#_c_396_n N_VPWR_c_475_n 0.040548f $X=2.975 $Y=2.275 $X2=0
+ $Y2=0
cc_321 N_A_27_297#_c_398_n N_VPWR_c_475_n 2.34313e-19 $X=2.98 $Y=2.2 $X2=0 $Y2=0
cc_322 N_A_27_297#_c_400_n N_VPWR_c_475_n 6.77819e-19 $X=5.89 $Y=2.21 $X2=0
+ $Y2=0
cc_323 N_A_27_297#_c_420_p N_VPWR_c_475_n 0.0154637f $X=5.89 $Y=2.21 $X2=0 $Y2=0
cc_324 N_A_27_297#_c_401_n N_VPWR_c_475_n 0.00231517f $X=5.695 $Y=2.2 $X2=0
+ $Y2=0
cc_325 N_A_27_297#_M1003_s N_VPWR_c_471_n 0.00358889f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_326 N_A_27_297#_M1009_s N_VPWR_c_471_n 0.00370124f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_327 N_A_27_297#_M1016_s N_VPWR_c_471_n 0.00297222f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_328 N_A_27_297#_M1018_s N_VPWR_c_471_n 0.00138294f $X=2.955 $Y=1.485 $X2=0
+ $Y2=0
cc_329 N_A_27_297#_M1022_s N_VPWR_c_471_n 0.00113892f $X=5.775 $Y=1.485 $X2=0
+ $Y2=0
cc_330 N_A_27_297#_c_427_p N_VPWR_c_471_n 0.00974347f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_331 N_A_27_297#_c_413_p N_VPWR_c_471_n 0.00955092f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_332 N_A_27_297#_c_415_p N_VPWR_c_471_n 0.00962794f $X=2.16 $Y=2.085 $X2=0
+ $Y2=0
cc_333 N_A_27_297#_c_416_p N_VPWR_c_471_n 0.00270511f $X=3.1 $Y=2.085 $X2=0
+ $Y2=0
cc_334 N_A_27_297#_c_396_n N_VPWR_c_471_n 0.0151721f $X=2.975 $Y=2.275 $X2=0
+ $Y2=0
cc_335 N_A_27_297#_c_398_n N_VPWR_c_471_n 0.0347312f $X=2.98 $Y=2.2 $X2=0 $Y2=0
cc_336 N_A_27_297#_c_400_n N_VPWR_c_471_n 0.0351309f $X=5.89 $Y=2.21 $X2=0 $Y2=0
cc_337 N_A_27_297#_c_420_p N_VPWR_c_471_n 0.00228824f $X=5.89 $Y=2.21 $X2=0
+ $Y2=0
cc_338 N_A_27_297#_c_401_n N_VPWR_c_471_n 0.233713f $X=5.695 $Y=2.2 $X2=0 $Y2=0
cc_339 N_A_27_297#_c_427_p N_VPWR_c_477_n 0.0165369f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_340 N_A_27_297#_c_396_n N_A_497_297#_M1001_d 0.00309975f $X=2.975 $Y=2.275
+ $X2=-0.19 $Y2=1.305
cc_341 N_A_27_297#_c_398_n N_A_497_297#_M1001_d 0.00142656f $X=2.98 $Y=2.2
+ $X2=-0.19 $Y2=1.305
cc_342 N_A_27_297#_c_401_n N_A_497_297#_M1019_d 0.00108334f $X=5.695 $Y=2.2
+ $X2=0 $Y2=0
cc_343 N_A_27_297#_c_401_n N_A_497_297#_M1010_s 4.4742e-19 $X=5.695 $Y=2.2 $X2=0
+ $Y2=0
cc_344 N_A_27_297#_c_401_n N_A_497_297#_M1021_s 4.72165e-19 $X=5.695 $Y=2.2
+ $X2=0 $Y2=0
cc_345 N_A_27_297#_M1018_s N_A_497_297#_c_551_n 0.00183202f $X=2.955 $Y=1.485
+ $X2=0 $Y2=0
cc_346 N_A_27_297#_c_443_p N_A_497_297#_c_551_n 0.0138782f $X=3.1 $Y=1.96 $X2=0
+ $Y2=0
cc_347 N_A_27_297#_c_396_n N_A_497_297#_c_551_n 0.00349887f $X=2.975 $Y=2.275
+ $X2=0 $Y2=0
cc_348 N_A_27_297#_c_398_n N_A_497_297#_c_551_n 0.00440098f $X=2.98 $Y=2.2 $X2=0
+ $Y2=0
cc_349 N_A_27_297#_c_401_n N_A_497_297#_c_551_n 0.00676646f $X=5.695 $Y=2.2
+ $X2=0 $Y2=0
cc_350 N_A_27_297#_c_416_p N_A_497_297#_c_580_n 0.00395971f $X=3.1 $Y=2.085
+ $X2=0 $Y2=0
cc_351 N_A_27_297#_c_398_n N_A_497_297#_c_580_n 6.17524e-19 $X=2.98 $Y=2.2 $X2=0
+ $Y2=0
cc_352 N_A_27_297#_c_401_n N_A_497_297#_c_580_n 0.026552f $X=5.695 $Y=2.2 $X2=0
+ $Y2=0
cc_353 N_A_27_297#_c_401_n N_A_497_297#_c_566_n 0.0104158f $X=5.695 $Y=2.2 $X2=0
+ $Y2=0
cc_354 N_A_27_297#_c_401_n N_A_497_297#_c_568_n 0.00664335f $X=5.695 $Y=2.2
+ $X2=0 $Y2=0
cc_355 N_A_27_297#_c_382_n N_A_497_297#_c_553_n 0.00226124f $X=2.16 $Y=1.625
+ $X2=0 $Y2=0
cc_356 N_A_27_297#_c_396_n N_A_497_297#_c_553_n 0.0139523f $X=2.975 $Y=2.275
+ $X2=0 $Y2=0
cc_357 N_A_27_297#_c_398_n N_A_497_297#_c_553_n 0.00351885f $X=2.98 $Y=2.2 $X2=0
+ $Y2=0
cc_358 N_A_27_297#_c_401_n N_A_497_297#_c_588_n 0.0189729f $X=5.695 $Y=2.2 $X2=0
+ $Y2=0
cc_359 N_A_27_297#_c_400_n N_A_497_297#_c_589_n 0.00170527f $X=5.89 $Y=2.21
+ $X2=0 $Y2=0
cc_360 N_A_27_297#_c_420_p N_A_497_297#_c_589_n 0.00471166f $X=5.89 $Y=2.21
+ $X2=0 $Y2=0
cc_361 N_A_27_297#_c_401_n N_A_497_297#_c_589_n 0.0159469f $X=5.695 $Y=2.2 $X2=0
+ $Y2=0
cc_362 N_A_27_297#_c_401_n N_Y_M1006_d 0.00394772f $X=5.695 $Y=2.2 $X2=0 $Y2=0
cc_363 N_A_27_297#_c_401_n N_Y_M1015_d 0.00337752f $X=5.695 $Y=2.2 $X2=0 $Y2=0
cc_364 N_A_27_297#_c_381_n N_Y_c_619_n 3.18413e-19 $X=2.035 $Y=1.54 $X2=0 $Y2=0
cc_365 N_A_27_297#_c_382_n N_Y_c_619_n 0.00936521f $X=2.16 $Y=1.625 $X2=0 $Y2=0
cc_366 N_A_27_297#_c_401_n N_Y_c_667_n 0.0121827f $X=5.695 $Y=2.2 $X2=0 $Y2=0
cc_367 N_A_27_297#_M1022_s N_Y_c_630_n 0.0087808f $X=5.775 $Y=1.485 $X2=0 $Y2=0
cc_368 N_A_27_297#_c_400_n N_Y_c_630_n 0.0119586f $X=5.89 $Y=2.21 $X2=0 $Y2=0
cc_369 N_A_27_297#_c_420_p N_Y_c_630_n 0.0142669f $X=5.89 $Y=2.21 $X2=0 $Y2=0
cc_370 N_A_27_297#_c_401_n N_Y_c_630_n 0.0115553f $X=5.695 $Y=2.2 $X2=0 $Y2=0
cc_371 N_A_27_297#_c_401_n N_Y_c_680_n 0.00762843f $X=5.695 $Y=2.2 $X2=0 $Y2=0
cc_372 N_A_27_297#_c_400_n N_Y_c_682_n 0.00186067f $X=5.89 $Y=2.21 $X2=0 $Y2=0
cc_373 N_A_27_297#_c_401_n N_Y_c_682_n 0.00762843f $X=5.695 $Y=2.2 $X2=0 $Y2=0
cc_374 N_VPWR_c_471_n N_A_497_297#_M1001_d 0.00178143f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_375 N_VPWR_c_471_n N_A_497_297#_M1019_d 0.00139285f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_471_n N_A_497_297#_M1010_s 0.00129629f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_471_n N_A_497_297#_M1021_s 0.00134113f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_475_n N_A_497_297#_c_580_n 0.015002f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_379 N_VPWR_c_471_n N_A_497_297#_c_580_n 0.00271607f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_475_n N_A_497_297#_c_566_n 0.0386815f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_471_n N_A_497_297#_c_566_n 0.00614936f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_475_n N_A_497_297#_c_568_n 0.0386815f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_471_n N_A_497_297#_c_568_n 0.00615735f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_475_n N_A_497_297#_c_588_n 0.0143076f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_471_n N_A_497_297#_c_588_n 0.00252432f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_475_n N_A_497_297#_c_589_n 0.0143076f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_471_n N_A_497_297#_c_589_n 0.00252432f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_471_n N_Y_M1006_d 0.00130999f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_389 N_VPWR_c_471_n N_Y_M1015_d 0.00130546f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_471_n N_Y_c_630_n 0.0128562f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_391 N_A_497_297#_c_566_n N_Y_M1006_d 0.00330238f $X=4.385 $Y=2.38 $X2=0 $Y2=0
cc_392 N_A_497_297#_c_568_n N_Y_M1015_d 0.00330238f $X=5.325 $Y=2.38 $X2=0 $Y2=0
cc_393 N_A_497_297#_M1010_s N_Y_c_667_n 0.00335211f $X=4.365 $Y=1.485 $X2=0
+ $Y2=0
cc_394 N_A_497_297#_c_566_n N_Y_c_667_n 0.00400368f $X=4.385 $Y=2.38 $X2=0 $Y2=0
cc_395 N_A_497_297#_c_568_n N_Y_c_667_n 0.00400368f $X=5.325 $Y=2.38 $X2=0 $Y2=0
cc_396 N_A_497_297#_c_588_n N_Y_c_667_n 0.0123695f $X=4.51 $Y=2.3 $X2=0 $Y2=0
cc_397 N_A_497_297#_M1021_s N_Y_c_630_n 0.00361964f $X=5.305 $Y=1.485 $X2=0
+ $Y2=0
cc_398 N_A_497_297#_c_568_n N_Y_c_630_n 0.00383094f $X=5.325 $Y=2.38 $X2=0 $Y2=0
cc_399 N_A_497_297#_c_589_n N_Y_c_630_n 0.0117216f $X=5.45 $Y=2.3 $X2=0 $Y2=0
cc_400 N_A_497_297#_c_566_n N_Y_c_680_n 0.0105164f $X=4.385 $Y=2.38 $X2=0 $Y2=0
cc_401 N_A_497_297#_c_568_n N_Y_c_682_n 0.0105164f $X=5.325 $Y=2.38 $X2=0 $Y2=0
cc_402 N_Y_c_617_n N_VGND_M1013_d 0.00251047f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_403 N_Y_c_619_n N_VGND_M1020_d 0.00162089f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_404 N_Y_c_620_n N_VGND_M1007_s 0.00348805f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_405 N_Y_c_621_n N_VGND_M1000_s 0.00251047f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_406 N_Y_c_622_n N_VGND_M1008_s 0.00348805f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_407 N_Y_c_623_n N_VGND_M1017_s 0.00315681f $X=6.055 $Y=0.815 $X2=0 $Y2=0
cc_408 N_Y_c_618_n N_VGND_c_800_n 0.00835456f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_409 N_Y_c_632_n N_VGND_c_801_n 0.0223596f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_410 N_Y_c_617_n N_VGND_c_801_n 0.00266636f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_411 N_Y_c_632_n N_VGND_c_802_n 0.0183628f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_412 N_Y_c_617_n N_VGND_c_802_n 0.0127273f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_413 N_Y_c_619_n N_VGND_c_803_n 0.0122559f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_414 N_Y_c_647_n N_VGND_c_804_n 0.0183628f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_415 N_Y_c_620_n N_VGND_c_804_n 0.0131987f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_416 N_Y_c_663_n N_VGND_c_804_n 0.0223967f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_417 N_Y_c_663_n N_VGND_c_805_n 0.0183628f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_418 N_Y_c_621_n N_VGND_c_805_n 0.0127273f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_419 N_Y_c_699_n N_VGND_c_806_n 0.0183628f $X=4.51 $Y=0.39 $X2=0 $Y2=0
cc_420 N_Y_c_622_n N_VGND_c_806_n 0.0131987f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_421 N_Y_c_708_n N_VGND_c_806_n 0.0223967f $X=5.45 $Y=0.39 $X2=0 $Y2=0
cc_422 N_Y_c_623_n N_VGND_c_807_n 0.0127273f $X=6.055 $Y=0.815 $X2=0 $Y2=0
cc_423 N_Y_c_617_n N_VGND_c_808_n 0.00198695f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_424 N_Y_c_643_n N_VGND_c_808_n 0.0231806f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_425 N_Y_c_619_n N_VGND_c_808_n 0.00254521f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_426 N_Y_c_619_n N_VGND_c_810_n 0.00198695f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_427 N_Y_c_647_n N_VGND_c_810_n 0.0223596f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_428 N_Y_c_620_n N_VGND_c_810_n 0.00266636f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_429 N_Y_c_620_n N_VGND_c_812_n 0.00199443f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_430 N_Y_c_663_n N_VGND_c_812_n 0.0222529f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_431 N_Y_c_621_n N_VGND_c_812_n 0.00266636f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_432 N_Y_c_621_n N_VGND_c_814_n 0.00198695f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_433 N_Y_c_699_n N_VGND_c_814_n 0.0223596f $X=4.51 $Y=0.39 $X2=0 $Y2=0
cc_434 N_Y_c_622_n N_VGND_c_814_n 0.00266636f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_435 N_Y_c_622_n N_VGND_c_816_n 0.00199443f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_436 N_Y_c_708_n N_VGND_c_816_n 0.023074f $X=5.45 $Y=0.39 $X2=0 $Y2=0
cc_437 N_Y_c_623_n N_VGND_c_816_n 0.00254521f $X=6.055 $Y=0.815 $X2=0 $Y2=0
cc_438 N_Y_c_623_n N_VGND_c_818_n 0.00565615f $X=6.055 $Y=0.815 $X2=0 $Y2=0
cc_439 N_Y_M1004_s N_VGND_c_819_n 0.0025535f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_440 N_Y_M1014_s N_VGND_c_819_n 0.00304143f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_441 N_Y_M1005_d N_VGND_c_819_n 0.0025535f $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_442 N_Y_M1011_d N_VGND_c_819_n 0.00215201f $X=3.435 $Y=0.235 $X2=0 $Y2=0
cc_443 N_Y_M1002_d N_VGND_c_819_n 0.0025535f $X=4.325 $Y=0.235 $X2=0 $Y2=0
cc_444 N_Y_M1023_d N_VGND_c_819_n 0.00263993f $X=5.315 $Y=0.235 $X2=0 $Y2=0
cc_445 N_Y_c_632_n N_VGND_c_819_n 0.0141302f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_446 N_Y_c_617_n N_VGND_c_819_n 0.00972452f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_447 N_Y_c_643_n N_VGND_c_819_n 0.0143352f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_448 N_Y_c_619_n N_VGND_c_819_n 0.0094839f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_449 N_Y_c_647_n N_VGND_c_819_n 0.0141302f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_450 N_Y_c_620_n N_VGND_c_819_n 0.0100158f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_451 N_Y_c_663_n N_VGND_c_819_n 0.0139016f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_452 N_Y_c_621_n N_VGND_c_819_n 0.00972452f $X=4.295 $Y=0.815 $X2=0 $Y2=0
cc_453 N_Y_c_699_n N_VGND_c_819_n 0.0141302f $X=4.51 $Y=0.39 $X2=0 $Y2=0
cc_454 N_Y_c_622_n N_VGND_c_819_n 0.0100158f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_455 N_Y_c_708_n N_VGND_c_819_n 0.0141066f $X=5.45 $Y=0.39 $X2=0 $Y2=0
cc_456 N_Y_c_623_n N_VGND_c_819_n 0.0151477f $X=6.055 $Y=0.815 $X2=0 $Y2=0
