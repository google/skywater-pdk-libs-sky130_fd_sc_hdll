* File: sky130_fd_sc_hdll__a211o_4.pex.spice
* Created: Wed Sep  2 08:15:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A211O_4%A_79_204# 1 2 3 4 13 15 18 20 22 25 27 29
+ 32 34 36 39 41 52 54 55 56 57 59 63 65 67 69 70 71 72 74 79 91
c159 70 0 1.95691e-19 $X=2.545 $Y=1.505
c160 69 0 1.19052e-19 $X=2.502 $Y=1.185
c161 52 0 1.61215e-19 $X=2.507 $Y=1.045
c162 39 0 9.43382e-20 $X=2.42 $Y=0.56
r163 91 92 66.4119 $w=3.52e-07 $l=4.85e-07 $layer=POLY_cond $X=1.935 $Y=1.215
+ $X2=2.42 $Y2=1.215
r164 88 89 57.5114 $w=3.52e-07 $l=4.2e-07 $layer=POLY_cond $X=1.455 $Y=1.215
+ $X2=1.875 $Y2=1.215
r165 87 88 8.21591 $w=3.52e-07 $l=6e-08 $layer=POLY_cond $X=1.395 $Y=1.215
+ $X2=1.455 $Y2=1.215
r166 86 87 57.5114 $w=3.52e-07 $l=4.2e-07 $layer=POLY_cond $X=0.975 $Y=1.215
+ $X2=1.395 $Y2=1.215
r167 85 86 8.21591 $w=3.52e-07 $l=6e-08 $layer=POLY_cond $X=0.915 $Y=1.215
+ $X2=0.975 $Y2=1.215
r168 79 81 10.6146 $w=3.78e-07 $l=3.5e-07 $layer=LI1_cond $X=5.85 $Y=0.36
+ $X2=5.85 $Y2=0.71
r169 74 76 10.0081 $w=3.78e-07 $l=3.3e-07 $layer=LI1_cond $X=4.23 $Y=0.38
+ $X2=4.23 $Y2=0.71
r170 70 71 9.11278 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=2.545 $Y=1.505
+ $X2=2.545 $Y2=1.675
r171 68 76 4.80115 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.42 $Y=0.71
+ $X2=4.23 $Y2=0.71
r172 67 81 4.80115 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=5.66 $Y=0.71
+ $X2=5.85 $Y2=0.71
r173 67 68 72.3828 $w=1.88e-07 $l=1.24e-06 $layer=LI1_cond $X=5.66 $Y=0.71
+ $X2=4.42 $Y2=0.71
r174 66 72 6.34807 $w=1.9e-07 $l=1.23e-07 $layer=LI1_cond $X=3.27 $Y=0.71
+ $X2=3.147 $Y2=0.71
r175 65 76 4.80115 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.04 $Y=0.71
+ $X2=4.23 $Y2=0.71
r176 65 66 44.9474 $w=1.88e-07 $l=7.7e-07 $layer=LI1_cond $X=4.04 $Y=0.71
+ $X2=3.27 $Y2=0.71
r177 61 72 0.445202 $w=2.45e-07 $l=9.5e-08 $layer=LI1_cond $X=3.147 $Y=0.615
+ $X2=3.147 $Y2=0.71
r178 61 63 6.115 $w=2.43e-07 $l=1.3e-07 $layer=LI1_cond $X=3.147 $Y=0.615
+ $X2=3.147 $Y2=0.485
r179 57 59 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=2.705 $Y=1.955
+ $X2=3.695 $Y2=1.955
r180 55 72 6.34807 $w=1.9e-07 $l=1.22e-07 $layer=LI1_cond $X=3.025 $Y=0.71
+ $X2=3.147 $Y2=0.71
r181 55 56 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=3.025 $Y=0.71
+ $X2=2.62 $Y2=0.71
r182 54 57 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=2.617 $Y=1.87
+ $X2=2.705 $Y2=1.955
r183 54 71 12.3584 $w=1.73e-07 $l=1.95e-07 $layer=LI1_cond $X=2.617 $Y=1.87
+ $X2=2.617 $Y2=1.675
r184 52 69 6.06507 $w=2.3e-07 $l=1.42478e-07 $layer=LI1_cond $X=2.507 $Y=1.045
+ $X2=2.502 $Y2=1.185
r185 51 56 6.87974 $w=1.9e-07 $l=1.5331e-07 $layer=LI1_cond $X=2.507 $Y=0.805
+ $X2=2.62 $Y2=0.71
r186 51 52 12.2927 $w=2.23e-07 $l=2.4e-07 $layer=LI1_cond $X=2.507 $Y=0.805
+ $X2=2.507 $Y2=1.045
r187 49 69 6.06507 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=2.502 $Y=1.325
+ $X2=2.502 $Y2=1.185
r188 49 70 8.82722 $w=2.33e-07 $l=1.8e-07 $layer=LI1_cond $X=2.502 $Y=1.325
+ $X2=2.502 $Y2=1.505
r189 48 91 3.4233 $w=3.52e-07 $l=2.5e-08 $layer=POLY_cond $X=1.91 $Y=1.215
+ $X2=1.935 $Y2=1.215
r190 48 89 4.79261 $w=3.52e-07 $l=3.5e-08 $layer=POLY_cond $X=1.91 $Y=1.215
+ $X2=1.875 $Y2=1.215
r191 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.91
+ $Y=1.16 $X2=1.91 $Y2=1.16
r192 44 85 17.1165 $w=3.52e-07 $l=1.25e-07 $layer=POLY_cond $X=0.79 $Y=1.215
+ $X2=0.915 $Y2=1.215
r193 44 83 40.3949 $w=3.52e-07 $l=2.95e-07 $layer=POLY_cond $X=0.79 $Y=1.215
+ $X2=0.495 $Y2=1.215
r194 43 47 46.0977 $w=2.78e-07 $l=1.12e-06 $layer=LI1_cond $X=0.79 $Y=1.185
+ $X2=1.91 $Y2=1.185
r195 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.79
+ $Y=1.16 $X2=0.79 $Y2=1.16
r196 41 69 0.644758 $w=2.8e-07 $l=1.17e-07 $layer=LI1_cond $X=2.385 $Y=1.185
+ $X2=2.502 $Y2=1.185
r197 41 47 19.5504 $w=2.78e-07 $l=4.75e-07 $layer=LI1_cond $X=2.385 $Y=1.185
+ $X2=1.91 $Y2=1.185
r198 37 92 22.7654 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.42 $Y=1.02
+ $X2=2.42 $Y2=1.215
r199 37 39 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.42 $Y=1.02
+ $X2=2.42 $Y2=0.56
r200 34 91 18.4407 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=1.935 $Y=1.41
+ $X2=1.935 $Y2=1.215
r201 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.935 $Y=1.41
+ $X2=1.935 $Y2=1.985
r202 30 89 22.7654 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.875 $Y=1.02
+ $X2=1.875 $Y2=1.215
r203 30 32 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.875 $Y=1.02
+ $X2=1.875 $Y2=0.56
r204 27 88 18.4407 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.215
r205 27 29 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r206 23 87 22.7654 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.395 $Y=1.02
+ $X2=1.395 $Y2=1.215
r207 23 25 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.395 $Y=1.02
+ $X2=1.395 $Y2=0.56
r208 20 86 18.4407 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.215
r209 20 22 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.985
r210 16 85 22.7654 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.915 $Y=1.02
+ $X2=0.915 $Y2=1.215
r211 16 18 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.915 $Y=1.02
+ $X2=0.915 $Y2=0.56
r212 13 83 18.4407 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.215
r213 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r214 4 59 600 $w=1.7e-07 $l=5.39815e-07 $layer=licon1_PDIFF $count=1 $X=3.545
+ $Y=1.485 $X2=3.695 $Y2=1.955
r215 3 79 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=5.685
+ $Y=0.235 $X2=5.875 $Y2=0.36
r216 2 74 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=4.035
+ $Y=0.235 $X2=4.235 $Y2=0.38
r217 1 63 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.98
+ $Y=0.235 $X2=3.12 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_4%B1 3 5 7 8 10 11 13 14 17 20 23 29
c89 29 0 1.86691e-19 $X=4.41 $Y=1.16
c90 20 0 9.43382e-20 $X=2.875 $Y=1.16
c91 8 0 1.47328e-19 $X=4.455 $Y=1.41
c92 5 0 1.61215e-19 $X=2.975 $Y=1.41
c93 3 0 1.04186e-19 $X=2.905 $Y=0.56
r94 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.41
+ $Y=1.16 $X2=4.41 $Y2=1.16
r95 23 29 7.35129 $w=5.48e-07 $l=2.85e-07 $layer=LI1_cond $X=4.435 $Y=1.445
+ $X2=4.435 $Y2=1.16
r96 20 22 18.6163 $w=2.7e-07 $l=4.12e-07 $layer=LI1_cond $X=2.947 $Y=1.16
+ $X2=2.947 $Y2=1.572
r97 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.875
+ $Y=1.16 $X2=2.875 $Y2=1.16
r98 15 22 1.08521 $w=2.55e-07 $l=1.58e-07 $layer=LI1_cond $X=3.105 $Y=1.572
+ $X2=2.947 $Y2=1.572
r99 15 17 36.607 $w=2.53e-07 $l=8.1e-07 $layer=LI1_cond $X=3.105 $Y=1.572
+ $X2=3.915 $Y2=1.572
r100 14 23 4.29494 $w=2.55e-07 $l=1.9e-07 $layer=LI1_cond $X=4.245 $Y=1.572
+ $X2=4.435 $Y2=1.572
r101 14 17 14.914 $w=2.53e-07 $l=3.3e-07 $layer=LI1_cond $X=4.245 $Y=1.572
+ $X2=3.915 $Y2=1.572
r102 11 28 40.1936 $w=3.54e-07 $l=2.25278e-07 $layer=POLY_cond $X=4.55 $Y=0.985
+ $X2=4.435 $Y2=1.16
r103 11 13 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.55 $Y=0.985
+ $X2=4.55 $Y2=0.56
r104 8 28 45.6582 $w=3.54e-07 $l=2.59808e-07 $layer=POLY_cond $X=4.455 $Y=1.41
+ $X2=4.435 $Y2=1.16
r105 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.455 $Y=1.41
+ $X2=4.455 $Y2=1.985
r106 5 21 45.7096 $w=3.52e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.975 $Y=1.41
+ $X2=2.9 $Y2=1.16
r107 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.975 $Y=1.41
+ $X2=2.975 $Y2=1.985
r108 1 21 35.3842 $w=3.52e-07 $l=1.42478e-07 $layer=POLY_cond $X=2.905 $Y=1.02
+ $X2=2.9 $Y2=1.16
r109 1 3 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.905 $Y=1.02
+ $X2=2.905 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_4%C1 1 3 4 6 7 9 10 12 13 20 23
c46 13 0 1.04186e-19 $X=3.83 $Y=1.105
r47 20 21 3.05838 $w=3.94e-07 $l=2.5e-08 $layer=POLY_cond $X=3.935 $Y=1.2
+ $X2=3.96 $Y2=1.2
r48 18 20 12.8452 $w=3.94e-07 $l=1.05e-07 $layer=POLY_cond $X=3.83 $Y=1.2
+ $X2=3.935 $Y2=1.2
r49 16 18 45.8756 $w=3.94e-07 $l=3.75e-07 $layer=POLY_cond $X=3.455 $Y=1.2
+ $X2=3.83 $Y2=1.2
r50 15 16 9.7868 $w=3.94e-07 $l=8e-08 $layer=POLY_cond $X=3.375 $Y=1.2 $X2=3.455
+ $Y2=1.2
r51 13 23 14.9023 $w=2.88e-07 $l=3.75e-07 $layer=LI1_cond $X=3.83 $Y=1.13
+ $X2=3.455 $Y2=1.13
r52 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.83
+ $Y=1.16 $X2=3.83 $Y2=1.16
r53 10 21 25.4929 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.96 $Y=0.99
+ $X2=3.96 $Y2=1.2
r54 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.96 $Y=0.99
+ $X2=3.96 $Y2=0.56
r55 7 20 21.1025 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.935 $Y=1.41
+ $X2=3.935 $Y2=1.2
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.935 $Y=1.41
+ $X2=3.935 $Y2=1.985
r57 4 16 21.1025 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.455 $Y=1.41
+ $X2=3.455 $Y2=1.2
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.455 $Y=1.41
+ $X2=3.455 $Y2=1.985
r59 1 15 25.4929 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.375 $Y=0.99
+ $X2=3.375 $Y2=1.2
r60 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.375 $Y=0.99
+ $X2=3.375 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_4%A2 1 3 6 8 10 11 13 16 19 21 24 26 32 36
c72 11 0 1.56978e-19 $X=6.595 $Y=1.41
c73 6 0 1.86691e-19 $X=5.18 $Y=0.56
r74 26 32 2.76019 $w=3.2e-07 $l=9.5e-08 $layer=LI1_cond $X=6.285 $Y=1.605
+ $X2=6.285 $Y2=1.51
r75 26 36 15.9107 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=6.125 $Y=1.605
+ $X2=5.755 $Y2=1.605
r76 26 32 1.18846 $w=3.18e-07 $l=3.3e-08 $layer=LI1_cond $X=6.285 $Y=1.477
+ $X2=6.285 $Y2=1.51
r77 25 26 5.65417 $w=3.18e-07 $l=1.57e-07 $layer=LI1_cond $X=6.285 $Y=1.32
+ $X2=6.285 $Y2=1.477
r78 24 36 25.1005 $w=1.88e-07 $l=4.3e-07 $layer=LI1_cond $X=5.325 $Y=1.605
+ $X2=5.755 $Y2=1.605
r79 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.16 $X2=6.66 $Y2=1.16
r80 19 25 6.82572 $w=3e-07 $l=2.22711e-07 $layer=LI1_cond $X=6.445 $Y=1.17
+ $X2=6.285 $Y2=1.32
r81 19 21 8.25918 $w=2.98e-07 $l=2.15e-07 $layer=LI1_cond $X=6.445 $Y=1.17
+ $X2=6.66 $Y2=1.17
r82 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.11
+ $Y=1.16 $X2=5.11 $Y2=1.16
r83 14 24 7.85115 $w=1.9e-07 $l=2.32702e-07 $layer=LI1_cond $X=5.135 $Y=1.51
+ $X2=5.325 $Y2=1.605
r84 14 16 10.6146 $w=3.78e-07 $l=3.5e-07 $layer=LI1_cond $X=5.135 $Y=1.51
+ $X2=5.135 $Y2=1.16
r85 11 22 45.6837 $w=3.53e-07 $l=2.91548e-07 $layer=POLY_cond $X=6.595 $Y=1.41
+ $X2=6.685 $Y2=1.16
r86 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.595 $Y=1.41
+ $X2=6.595 $Y2=1.985
r87 8 22 36.7715 $w=3.53e-07 $l=1.99374e-07 $layer=POLY_cond $X=6.57 $Y=1.01
+ $X2=6.685 $Y2=1.16
r88 8 10 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.57 $Y=1.01 $X2=6.57
+ $Y2=0.56
r89 4 17 35.9216 $w=3.75e-07 $l=1.60935e-07 $layer=POLY_cond $X=5.18 $Y=1.02
+ $X2=5.135 $Y2=1.16
r90 4 6 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=5.18 $Y=1.02 $X2=5.18
+ $Y2=0.56
r91 1 17 45.2166 $w=3.75e-07 $l=2.91548e-07 $layer=POLY_cond $X=5.045 $Y=1.41
+ $X2=5.135 $Y2=1.16
r92 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.045 $Y=1.41
+ $X2=5.045 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_4%A1 3 5 7 8 10 13 15 22 25
c46 15 0 3.16013e-19 $X=5.66 $Y=1.105
r47 22 23 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=6.115 $Y=1.215
+ $X2=6.14 $Y2=1.215
r48 20 22 54.8027 $w=3.65e-07 $l=4.15e-07 $layer=POLY_cond $X=5.7 $Y=1.215
+ $X2=6.115 $Y2=1.215
r49 18 20 8.58356 $w=3.65e-07 $l=6.5e-08 $layer=POLY_cond $X=5.635 $Y=1.215
+ $X2=5.7 $Y2=1.215
r50 17 18 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=5.61 $Y=1.215
+ $X2=5.635 $Y2=1.215
r51 15 25 4.64695 $w=3.08e-07 $l=1.25e-07 $layer=LI1_cond $X=5.7 $Y=1.175
+ $X2=5.575 $Y2=1.175
r52 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.7
+ $Y=1.16 $X2=5.7 $Y2=1.16
r53 11 23 23.6381 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=6.14 $Y=1.02
+ $X2=6.14 $Y2=1.215
r54 11 13 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=6.14 $Y=1.02
+ $X2=6.14 $Y2=0.56
r55 8 22 19.2931 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=6.115 $Y=1.41
+ $X2=6.115 $Y2=1.215
r56 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.115 $Y=1.41
+ $X2=6.115 $Y2=1.985
r57 5 18 19.2931 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=5.635 $Y=1.41
+ $X2=5.635 $Y2=1.215
r58 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.635 $Y=1.41
+ $X2=5.635 $Y2=1.985
r59 1 17 23.6381 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=5.61 $Y=1.02
+ $X2=5.61 $Y2=1.215
r60 1 3 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=5.61 $Y=1.02 $X2=5.61
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_4%VPWR 1 2 3 4 5 16 18 22 24 28 30 32 34 39
+ 49 50 56 59 62 69
c107 1 0 1.48954e-19 $X=0.135 $Y=1.485
r108 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r109 69 72 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=6.33 $Y=2.36
+ $X2=6.33 $Y2=2.72
r110 66 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r112 62 65 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.26 $Y=2.36
+ $X2=5.26 $Y2=2.72
r113 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r114 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r115 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r116 50 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.21 $Y2=2.72
r117 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r118 47 72 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.52 $Y=2.72
+ $X2=6.33 $Y2=2.72
r119 47 49 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.52 $Y=2.72
+ $X2=7.13 $Y2=2.72
r120 46 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r121 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r122 43 46 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r123 43 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 42 45 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r125 42 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r126 40 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.26 $Y=2.72
+ $X2=2.135 $Y2=2.72
r127 40 42 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.26 $Y=2.72
+ $X2=2.53 $Y2=2.72
r128 39 65 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.07 $Y=2.72
+ $X2=5.26 $Y2=2.72
r129 39 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.07 $Y=2.72
+ $X2=4.83 $Y2=2.72
r130 38 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r131 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r132 35 53 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r133 35 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r134 34 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.05 $Y=2.72
+ $X2=1.215 $Y2=2.72
r135 34 37 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.05 $Y=2.72
+ $X2=0.69 $Y2=2.72
r136 32 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r137 32 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r138 31 65 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.45 $Y=2.72
+ $X2=5.26 $Y2=2.72
r139 30 72 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.14 $Y=2.72
+ $X2=6.33 $Y2=2.72
r140 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.14 $Y=2.72
+ $X2=5.45 $Y2=2.72
r141 26 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=2.635
+ $X2=2.135 $Y2=2.72
r142 26 28 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.135 $Y=2.635
+ $X2=2.135 $Y2=2
r143 25 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=2.72
+ $X2=1.215 $Y2=2.72
r144 24 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.01 $Y=2.72
+ $X2=2.135 $Y2=2.72
r145 24 25 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.01 $Y=2.72
+ $X2=1.38 $Y2=2.72
r146 20 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.635
+ $X2=1.215 $Y2=2.72
r147 20 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.215 $Y=2.635
+ $X2=1.215 $Y2=1.96
r148 16 53 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r149 16 18 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=1.96
r150 5 69 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.485 $X2=6.355 $Y2=2.36
r151 4 62 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=5.135
+ $Y=1.485 $X2=5.285 $Y2=2.36
r152 3 28 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.025
+ $Y=1.485 $X2=2.17 $Y2=2
r153 2 22 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=1.485 $X2=1.215 $Y2=1.96
r154 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_4%X 1 2 3 4 13 15 16 19 21 25 27 31 35 38 39
+ 40 43
c65 40 0 1.48954e-19 $X=0.23 $Y=0.85
r66 40 43 3.30224 $w=2.55e-07 $l=1.2e-07 $layer=LI1_cond $X=0.212 $Y=0.755
+ $X2=0.212 $Y2=0.875
r67 40 43 1.35582 $w=2.53e-07 $l=3e-08 $layer=LI1_cond $X=0.212 $Y=0.905
+ $X2=0.212 $Y2=0.875
r68 37 40 26.6644 $w=2.53e-07 $l=5.9e-07 $layer=LI1_cond $X=0.212 $Y=1.495
+ $X2=0.212 $Y2=0.905
r69 33 35 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=2.135 $Y=0.615
+ $X2=2.135 $Y2=0.42
r70 29 31 8.75598 $w=1.88e-07 $l=1.5e-07 $layer=LI1_cond $X=1.695 $Y=1.705
+ $X2=1.695 $Y2=1.855
r71 28 39 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=1.275 $Y=0.745
+ $X2=1.18 $Y2=0.745
r72 27 33 7.11373 $w=2.6e-07 $l=1.69115e-07 $layer=LI1_cond $X=2.045 $Y=0.745
+ $X2=2.135 $Y2=0.615
r73 27 28 34.13 $w=2.58e-07 $l=7.7e-07 $layer=LI1_cond $X=2.045 $Y=0.745
+ $X2=1.275 $Y2=0.745
r74 23 39 2.34704 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=1.18 $Y=0.615
+ $X2=1.18 $Y2=0.745
r75 23 25 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.18 $Y=0.615
+ $X2=1.18 $Y2=0.42
r76 22 38 4.64301 $w=2.1e-07 $l=9.3e-08 $layer=LI1_cond $X=0.83 $Y=1.6 $X2=0.737
+ $Y2=1.6
r77 21 29 6.83868 $w=2.1e-07 $l=1.44914e-07 $layer=LI1_cond $X=1.6 $Y=1.6
+ $X2=1.695 $Y2=1.705
r78 21 22 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=1.6 $Y=1.6 $X2=0.83
+ $Y2=1.6
r79 17 38 1.80272 $w=1.85e-07 $l=1.05e-07 $layer=LI1_cond $X=0.737 $Y=1.705
+ $X2=0.737 $Y2=1.6
r80 17 19 8.99263 $w=1.83e-07 $l=1.5e-07 $layer=LI1_cond $X=0.737 $Y=1.705
+ $X2=0.737 $Y2=1.855
r81 16 37 6.89985 $w=2.1e-07 $l=1.72696e-07 $layer=LI1_cond $X=0.34 $Y=1.6
+ $X2=0.212 $Y2=1.495
r82 15 38 4.64301 $w=2.1e-07 $l=9.2e-08 $layer=LI1_cond $X=0.645 $Y=1.6
+ $X2=0.737 $Y2=1.6
r83 15 16 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=0.645 $Y=1.6
+ $X2=0.34 $Y2=1.6
r84 14 40 3.52239 $w=2.4e-07 $l=1.28e-07 $layer=LI1_cond $X=0.34 $Y=0.755
+ $X2=0.212 $Y2=0.755
r85 13 39 4.08801 $w=2.5e-07 $l=9.98749e-08 $layer=LI1_cond $X=1.085 $Y=0.755
+ $X2=1.18 $Y2=0.745
r86 13 14 35.7738 $w=2.38e-07 $l=7.45e-07 $layer=LI1_cond $X=1.085 $Y=0.755
+ $X2=0.34 $Y2=0.755
r87 4 31 300 $w=1.7e-07 $l=4.38634e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.695 $Y2=1.855
r88 3 19 300 $w=1.7e-07 $l=4.38634e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.735 $Y2=1.855
r89 2 35 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.235 $X2=2.14 $Y2=0.42
r90 1 25 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.235 $X2=1.18 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_4%A_523_297# 1 2 3 4 13 17 21 23 27 29 35 37
c64 29 0 1.47328e-19 $X=4.735 $Y=1.992
c65 1 0 1.95691e-19 $X=2.615 $Y=1.485
r66 39 40 4.67835 $w=3.78e-07 $l=1.13e-07 $layer=LI1_cond $X=6.805 $Y=1.992
+ $X2=6.805 $Y2=2.105
r67 37 39 10.9785 $w=3.78e-07 $l=3.62e-07 $layer=LI1_cond $X=6.805 $Y=1.63
+ $X2=6.805 $Y2=1.992
r68 32 33 11.7689 $w=3.28e-07 $l=3.37e-07 $layer=LI1_cond $X=4.735 $Y=2
+ $X2=4.735 $Y2=2.337
r69 29 32 0.27938 $w=3.28e-07 $l=8e-09 $layer=LI1_cond $X=4.735 $Y=1.992
+ $X2=4.735 $Y2=2
r70 27 40 8.8128 $w=2.53e-07 $l=1.95e-07 $layer=LI1_cond $X=6.867 $Y=2.3
+ $X2=6.867 $Y2=2.105
r71 24 35 6.68507 $w=2.25e-07 $l=1.55e-07 $layer=LI1_cond $X=5.97 $Y=1.992
+ $X2=5.815 $Y2=1.992
r72 23 39 3.81936 $w=2.25e-07 $l=1.9e-07 $layer=LI1_cond $X=6.615 $Y=1.992
+ $X2=6.805 $Y2=1.992
r73 23 24 33.0367 $w=2.23e-07 $l=6.45e-07 $layer=LI1_cond $X=6.615 $Y=1.992
+ $X2=5.97 $Y2=1.992
r74 19 35 0.218322 $w=3.1e-07 $l=1.13e-07 $layer=LI1_cond $X=5.815 $Y=2.105
+ $X2=5.815 $Y2=1.992
r75 19 21 7.24924 $w=3.08e-07 $l=1.95e-07 $layer=LI1_cond $X=5.815 $Y=2.105
+ $X2=5.815 $Y2=2.3
r76 18 29 2.99809 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.992
+ $X2=4.735 $Y2=1.992
r77 17 35 6.68507 $w=2.25e-07 $l=1.55e-07 $layer=LI1_cond $X=5.66 $Y=1.992
+ $X2=5.815 $Y2=1.992
r78 17 18 38.927 $w=2.23e-07 $l=7.6e-07 $layer=LI1_cond $X=5.66 $Y=1.992 $X2=4.9
+ $Y2=1.992
r79 13 33 2.26808 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=4.57 $Y=2.337
+ $X2=4.735 $Y2=2.337
r80 13 15 82.7047 $w=2.53e-07 $l=1.83e-06 $layer=LI1_cond $X=4.57 $Y=2.337
+ $X2=2.74 $Y2=2.337
r81 4 37 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.685
+ $Y=1.485 $X2=6.83 $Y2=1.63
r82 4 27 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.685
+ $Y=1.485 $X2=6.83 $Y2=2.3
r83 3 21 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=5.725
+ $Y=1.485 $X2=5.875 $Y2=2.3
r84 2 32 300 $w=1.7e-07 $l=6.02557e-07 $layer=licon1_PDIFF $count=2 $X=4.545
+ $Y=1.485 $X2=4.735 $Y2=2
r85 1 15 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.615
+ $Y=1.485 $X2=2.74 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_4%VGND 1 2 3 4 5 6 19 23 25 27 32 37 42 47
+ 54 55 59 66 80 87 93
r104 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r105 87 90 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.825 $Y=0 $X2=4.825
+ $Y2=0.36
r106 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r107 80 83 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.63 $Y=0 $X2=3.63
+ $Y2=0.36
r108 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r109 74 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r110 66 69 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.635 $Y=0
+ $X2=1.635 $Y2=0.36
r111 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r112 59 62 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.675 $Y=0
+ $X2=0.675 $Y2=0.38
r113 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r114 55 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=6.67
+ $Y2=0
r115 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r116 52 93 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.995 $Y=0 $X2=6.805
+ $Y2=0
r117 52 54 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.995 $Y=0
+ $X2=7.13 $Y2=0
r118 51 94 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r119 51 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r120 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r121 48 87 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.01 $Y=0 $X2=4.825
+ $Y2=0
r122 48 50 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.01 $Y=0 $X2=5.29
+ $Y2=0
r123 47 93 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.615 $Y=0 $X2=6.805
+ $Y2=0
r124 47 50 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=6.615 $Y=0
+ $X2=5.29 $Y2=0
r125 46 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r126 46 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r127 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r128 43 80 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.82 $Y=0 $X2=3.63
+ $Y2=0
r129 43 45 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.82 $Y=0 $X2=4.37
+ $Y2=0
r130 42 87 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.64 $Y=0 $X2=4.825
+ $Y2=0
r131 42 45 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.64 $Y=0 $X2=4.37
+ $Y2=0
r132 41 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r133 41 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r134 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r135 38 66 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.635
+ $Y2=0
r136 38 40 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=2.07
+ $Y2=0
r137 37 76 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=2.612 $Y=0
+ $X2=2.612 $Y2=0.36
r138 37 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r139 37 40 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.07
+ $Y2=0
r140 36 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r141 36 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r142 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r143 33 59 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.675
+ $Y2=0
r144 33 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.865 $Y=0
+ $X2=1.15 $Y2=0
r145 32 66 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.635
+ $Y2=0
r146 32 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.15
+ $Y2=0
r147 27 59 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.485 $Y=0 $X2=0.675
+ $Y2=0
r148 27 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.485 $Y=0
+ $X2=0.23 $Y2=0
r149 25 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r150 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r151 21 93 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.805 $Y=0.085
+ $X2=6.805 $Y2=0
r152 21 23 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=6.805 $Y=0.085
+ $X2=6.805 $Y2=0.38
r153 20 37 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.805 $Y=0
+ $X2=2.612 $Y2=0
r154 19 80 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.63
+ $Y2=0
r155 19 20 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.44 $Y=0
+ $X2=2.805 $Y2=0
r156 6 23 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=6.645
+ $Y=0.235 $X2=6.83 $Y2=0.38
r157 5 90 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.235 $X2=4.805 $Y2=0.36
r158 4 83 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.235 $X2=3.655 $Y2=0.36
r159 3 76 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.235 $X2=2.64 $Y2=0.36
r160 2 69 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.47
+ $Y=0.235 $X2=1.66 $Y2=0.36
r161 1 62 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=0.525
+ $Y=0.235 $X2=0.7 $Y2=0.38
.ends

