* File: sky130_fd_sc_hdll__mux2i_4.pex.spice
* Created: Wed Sep  2 08:35:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%A0 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 38 43 47
r62 38 39 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r63 37 38 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.905 $Y2=1.202
r64 36 37 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r65 35 43 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=0.695 $Y2=1.16
r66 34 36 48.5887 $w=3.72e-07 $l=3.75e-07 $layer=POLY_cond $X=1.035 $Y=1.202
+ $X2=1.41 $Y2=1.202
r67 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.035
+ $Y=1.16 $X2=1.035 $Y2=1.16
r68 32 34 9.06989 $w=3.72e-07 $l=7e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.035 $Y2=1.202
r69 31 32 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r70 30 31 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.94 $Y2=1.202
r71 29 30 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r72 26 47 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.155 $Y2=1.16
r73 26 35 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.035 $Y2=1.16
r74 25 43 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.695 $Y2=1.16
r75 22 39 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r76 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r77 19 38 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r78 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r79 16 37 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r80 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r81 13 36 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r82 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r83 10 32 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r84 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r85 7 31 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r86 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
r87 4 30 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r88 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r89 1 29 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r90 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 45 51 54 57 61
r70 45 46 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.81 $Y2=1.202
r71 44 57 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.61 $Y=1.16
+ $X2=3.455 $Y2=1.16
r72 43 45 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=3.61 $Y=1.202
+ $X2=3.785 $Y2=1.202
r73 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.61
+ $Y=1.16 $X2=3.61 $Y2=1.16
r74 41 43 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.61 $Y2=1.202
r75 40 41 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r76 39 40 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.29 $Y2=1.202
r77 38 39 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r78 36 38 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=2.44 $Y=1.202
+ $X2=2.82 $Y2=1.202
r79 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.44
+ $Y=1.16 $X2=2.44 $Y2=1.16
r80 34 36 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.44 $Y2=1.202
r81 33 34 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r82 28 61 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=3.907 $Y=1.16
+ $X2=3.925 $Y2=1.16
r83 28 44 10.372 $w=3.28e-07 $l=2.97e-07 $layer=LI1_cond $X=3.907 $Y=1.16
+ $X2=3.61 $Y2=1.16
r84 27 57 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.45 $Y=1.16
+ $X2=3.455 $Y2=1.16
r85 27 54 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=1.16
+ $X2=2.995 $Y2=1.16
r86 26 54 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=1.16
+ $X2=2.995 $Y2=1.16
r87 26 51 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2.99 $Y=1.16
+ $X2=2.535 $Y2=1.16
r88 25 51 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.53 $Y=1.16
+ $X2=2.535 $Y2=1.16
r89 25 37 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.53 $Y=1.16 $X2=2.44
+ $Y2=1.16
r90 22 46 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r91 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r92 19 45 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r93 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r94 16 41 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r95 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r96 13 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r97 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
r98 10 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r99 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r100 7 38 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r102 4 34 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r103 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r104 1 33 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r105 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%S 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 35 39 43 44 45 46 47 65 71 75 78 81 85
r132 65 66 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.21 $Y2=1.202
r133 64 81 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=6.07 $Y=1.182
+ $X2=5.775 $Y2=1.182
r134 63 65 15.1863 $w=3.65e-07 $l=1.15e-07 $layer=POLY_cond $X=6.07 $Y=1.202
+ $X2=6.185 $Y2=1.202
r135 63 64 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.07
+ $Y=1.16 $X2=6.07 $Y2=1.16
r136 61 63 43.5781 $w=3.65e-07 $l=3.3e-07 $layer=POLY_cond $X=5.74 $Y=1.202
+ $X2=6.07 $Y2=1.202
r137 60 61 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=5.715 $Y=1.202
+ $X2=5.74 $Y2=1.202
r138 59 60 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=5.27 $Y=1.202
+ $X2=5.715 $Y2=1.202
r139 58 59 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=5.245 $Y=1.202
+ $X2=5.27 $Y2=1.202
r140 57 58 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=4.8 $Y=1.202
+ $X2=5.245 $Y2=1.202
r141 56 57 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.8 $Y2=1.202
r142 55 71 8.84433 $w=2.13e-07 $l=1.65e-07 $layer=LI1_cond $X=4.56 $Y=1.182
+ $X2=4.395 $Y2=1.182
r143 54 56 28.3918 $w=3.65e-07 $l=2.15e-07 $layer=POLY_cond $X=4.56 $Y=1.202
+ $X2=4.775 $Y2=1.202
r144 54 55 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.56
+ $Y=1.16 $X2=4.56 $Y2=1.16
r145 47 85 1.07204 $w=2.13e-07 $l=2e-08 $layer=LI1_cond $X=6.21 $Y=1.182
+ $X2=6.23 $Y2=1.182
r146 47 64 7.50428 $w=2.13e-07 $l=1.4e-07 $layer=LI1_cond $X=6.21 $Y=1.182
+ $X2=6.07 $Y2=1.182
r147 46 81 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=5.75 $Y=1.182
+ $X2=5.775 $Y2=1.182
r148 46 78 23.3169 $w=2.13e-07 $l=4.35e-07 $layer=LI1_cond $X=5.75 $Y=1.182
+ $X2=5.315 $Y2=1.182
r149 45 78 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=5.29 $Y=1.182
+ $X2=5.315 $Y2=1.182
r150 45 75 23.3169 $w=2.13e-07 $l=4.35e-07 $layer=LI1_cond $X=5.29 $Y=1.182
+ $X2=4.855 $Y2=1.182
r151 44 75 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=4.83 $Y=1.182
+ $X2=4.855 $Y2=1.182
r152 44 55 14.4725 $w=2.13e-07 $l=2.7e-07 $layer=LI1_cond $X=4.83 $Y=1.182
+ $X2=4.56 $Y2=1.182
r153 43 71 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=4.37 $Y=1.182
+ $X2=4.395 $Y2=1.182
r154 39 85 6.96826 $w=2.13e-07 $l=1.3e-07 $layer=LI1_cond $X=6.36 $Y=1.182
+ $X2=6.23 $Y2=1.182
r155 39 41 21.3989 $w=1.68e-07 $l=3.28e-07 $layer=LI1_cond $X=6.445 $Y=1.182
+ $X2=6.445 $Y2=1.51
r156 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.565
+ $Y=1.16 $X2=8.565 $Y2=1.16
r157 33 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.565 $Y=1.425
+ $X2=8.565 $Y2=1.16
r158 32 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=1.51
+ $X2=6.445 $Y2=1.51
r159 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.48 $Y=1.51
+ $X2=8.565 $Y2=1.425
r160 31 32 127.219 $w=1.68e-07 $l=1.95e-06 $layer=LI1_cond $X=8.48 $Y=1.51
+ $X2=6.53 $Y2=1.51
r161 28 36 38.578 $w=2.95e-07 $l=1.96914e-07 $layer=POLY_cond $X=8.66 $Y=0.995
+ $X2=8.59 $Y2=1.16
r162 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.66 $Y=0.995
+ $X2=8.66 $Y2=0.56
r163 25 36 48.1208 $w=2.95e-07 $l=2.7157e-07 $layer=POLY_cond $X=8.635 $Y=1.41
+ $X2=8.59 $Y2=1.16
r164 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.635 $Y=1.41
+ $X2=8.635 $Y2=1.985
r165 22 66 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.21 $Y=0.995
+ $X2=6.21 $Y2=1.202
r166 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.21 $Y=0.995
+ $X2=6.21 $Y2=0.56
r167 19 65 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r168 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r169 16 61 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=1.202
r170 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=0.56
r171 13 60 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r172 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r173 10 59 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=1.202
r174 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=0.56
r175 7 58 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.202
r176 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r177 4 57 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=1.202
r178 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=0.995 $X2=4.8
+ $Y2=0.56
r179 1 56 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r180 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%A_1311_21# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 37 38 39 42 44 46 50 51 59
c114 19 0 3.63796e-19 $X=7.57 $Y=0.995
r115 59 60 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=8.12 $Y=1.202
+ $X2=8.145 $Y2=1.202
r116 56 57 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.57 $Y=1.202
+ $X2=7.595 $Y2=1.202
r117 55 56 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=7.125 $Y=1.202
+ $X2=7.57 $Y2=1.202
r118 54 55 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.1 $Y=1.202
+ $X2=7.125 $Y2=1.202
r119 53 54 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=6.655 $Y=1.202
+ $X2=7.1 $Y2=1.202
r120 52 53 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.63 $Y=1.202
+ $X2=6.655 $Y2=1.202
r121 48 50 4.18896 $w=2.17e-07 $l=1.03899e-07 $layer=LI1_cond $X=8.957 $Y=0.825
+ $X2=8.915 $Y2=0.74
r122 48 51 61.4753 $w=1.73e-07 $l=9.7e-07 $layer=LI1_cond $X=8.957 $Y=0.825
+ $X2=8.957 $Y2=1.795
r123 44 51 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=8.915 $Y=1.925
+ $X2=8.915 $Y2=1.795
r124 44 46 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=8.915 $Y=1.925
+ $X2=8.915 $Y2=1.96
r125 40 50 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=8.915 $Y=0.655
+ $X2=8.915 $Y2=0.74
r126 40 42 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=8.915 $Y=0.655
+ $X2=8.915 $Y2=0.42
r127 38 50 2.24312 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.785 $Y=0.74
+ $X2=8.915 $Y2=0.74
r128 38 39 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=8.785 $Y=0.74
+ $X2=8.31 $Y2=0.74
r129 36 39 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=8.2 $Y=0.825
+ $X2=8.31 $Y2=0.74
r130 36 37 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=8.2 $Y=0.825
+ $X2=8.2 $Y2=1.075
r131 34 59 14.9811 $w=3.7e-07 $l=1.15e-07 $layer=POLY_cond $X=8.005 $Y=1.202
+ $X2=8.12 $Y2=1.202
r132 34 57 53.4108 $w=3.7e-07 $l=4.1e-07 $layer=POLY_cond $X=8.005 $Y=1.202
+ $X2=7.595 $Y2=1.202
r133 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.005
+ $Y=1.16 $X2=8.005 $Y2=1.16
r134 31 37 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=8.09 $Y=1.16
+ $X2=8.2 $Y2=1.075
r135 31 33 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.09 $Y=1.16
+ $X2=8.005 $Y2=1.16
r136 28 60 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.145 $Y=0.995
+ $X2=8.145 $Y2=1.202
r137 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.145 $Y=0.995
+ $X2=8.145 $Y2=0.56
r138 25 59 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.12 $Y=1.41
+ $X2=8.12 $Y2=1.202
r139 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.12 $Y=1.41
+ $X2=8.12 $Y2=1.985
r140 22 57 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.202
r141 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.985
r142 19 56 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=1.202
r143 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=0.56
r144 16 55 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r145 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r146 13 54 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=1.202
r147 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=0.56
r148 10 53 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r149 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r150 7 52 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.202
r151 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.56
r152 2 46 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.725
+ $Y=1.485 $X2=8.87 $Y2=1.96
r153 1 42 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.235 $X2=8.87 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%Y 1 2 3 4 5 6 7 8 9 10 39 49 51 54 55 56
+ 57 58 65 76
r72 65 76 2.30489 $w=2.23e-07 $l=4.5e-08 $layer=LI1_cond $X=0.207 $Y=2.255
+ $X2=0.207 $Y2=2.21
r73 58 65 3.00067 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.207 $Y=2.34
+ $X2=0.207 $Y2=2.255
r74 58 76 1.02439 $w=2.23e-07 $l=2e-08 $layer=LI1_cond $X=0.207 $Y=2.19
+ $X2=0.207 $Y2=2.21
r75 57 58 16.3903 $w=2.23e-07 $l=3.2e-07 $layer=LI1_cond $X=0.207 $Y=1.87
+ $X2=0.207 $Y2=2.19
r76 56 57 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.53
+ $X2=0.207 $Y2=1.87
r77 55 56 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r78 54 55 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=0.85
+ $X2=0.207 $Y2=1.19
r79 51 54 18.6952 $w=2.23e-07 $l=3.65e-07 $layer=LI1_cond $X=0.207 $Y=0.485
+ $X2=0.207 $Y2=0.85
r80 51 53 3.00067 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.207 $Y=0.485
+ $X2=0.207 $Y2=0.4
r81 47 49 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.08 $Y=2.34
+ $X2=4.02 $Y2=2.34
r82 45 47 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.14 $Y=2.34
+ $X2=3.08 $Y2=2.34
r83 43 45 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.2 $Y=2.34 $X2=2.14
+ $Y2=2.34
r84 41 58 3.98913 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.32 $Y=2.34
+ $X2=0.207 $Y2=2.34
r85 41 43 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.32 $Y=2.34 $X2=1.2
+ $Y2=2.34
r86 37 39 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.08 $Y=0.4 $X2=4.02
+ $Y2=0.4
r87 35 37 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.14 $Y=0.4 $X2=3.08
+ $Y2=0.4
r88 33 35 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.2 $Y=0.4 $X2=2.14
+ $Y2=0.4
r89 31 53 3.98913 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.32 $Y=0.4
+ $X2=0.207 $Y2=0.4
r90 31 33 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.32 $Y=0.4 $X2=1.2
+ $Y2=0.4
r91 10 49 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2.34
r92 9 47 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2.34
r93 8 45 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.34
r94 7 43 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r95 6 58 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r96 5 39 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.4
r97 4 37 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.4
r98 3 35 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.4
r99 2 33 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.4
r100 1 53 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%A_117_297# 1 2 3 4 21
r41 19 21 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.01 $Y=1.66
+ $X2=5.95 $Y2=1.66
r42 17 19 217.904 $w=1.68e-07 $l=3.34e-06 $layer=LI1_cond $X=1.67 $Y=1.66
+ $X2=5.01 $Y2=1.66
r43 14 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.73 $Y=1.66
+ $X2=1.67 $Y2=1.66
r44 4 21 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.66
r45 3 19 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.66
r46 2 17 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r47 1 14 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%A_493_297# 1 2 3 4 13 21 23 25 27 30
r59 25 32 3.40825 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.83 $Y=2.085
+ $X2=7.83 $Y2=1.94
r60 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.83 $Y=2.085
+ $X2=7.83 $Y2=2.3
r61 24 30 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=6.975 $Y=2
+ $X2=6.89 $Y2=1.94
r62 23 32 3.40825 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=7.745 $Y=2
+ $X2=7.83 $Y2=1.94
r63 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.745 $Y=2 $X2=6.975
+ $Y2=2
r64 19 30 1.34256 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.89 $Y=2.085
+ $X2=6.89 $Y2=1.94
r65 19 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.89 $Y=2.085
+ $X2=6.89 $Y2=2.3
r66 15 18 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.61 $Y=2 $X2=3.55
+ $Y2=2
r67 13 30 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=6.805 $Y=2
+ $X2=6.89 $Y2=1.94
r68 13 18 212.358 $w=1.68e-07 $l=3.255e-06 $layer=LI1_cond $X=6.805 $Y=2
+ $X2=3.55 $Y2=2
r69 4 32 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.485 $X2=7.83 $Y2=1.96
r70 4 27 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.485 $X2=7.83 $Y2=2.3
r71 3 30 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.96
r72 3 21 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=2.3
r73 2 18 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2
r74 1 15 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%VPWR 1 2 3 4 5 18 20 22 26 28 29 31 34 38
+ 39 40 57 58 61 68
r117 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r118 68 71 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=6.395 $Y=2.34
+ $X2=6.395 $Y2=2.72
r119 65 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r120 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r121 61 64 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=5.455 $Y=2.34
+ $X2=5.455 $Y2=2.72
r122 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r123 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r124 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r125 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r126 52 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.21 $Y2=2.72
r127 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r128 49 71 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=6.395 $Y2=2.72
r129 49 51 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=7.13 $Y2=2.72
r130 48 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r131 47 48 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r132 43 47 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=4.37 $Y2=2.72
r133 40 48 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=4.37 $Y2=2.72
r134 40 43 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r135 38 54 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.235 $Y=2.72
+ $X2=8.05 $Y2=2.72
r136 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.235 $Y=2.72
+ $X2=8.4 $Y2=2.72
r137 37 57 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.565 $Y=2.72
+ $X2=8.97 $Y2=2.72
r138 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.565 $Y=2.72
+ $X2=8.4 $Y2=2.72
r139 35 54 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=7.525 $Y=2.72
+ $X2=8.05 $Y2=2.72
r140 34 51 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.145 $Y=2.72
+ $X2=7.13 $Y2=2.72
r141 33 35 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.525 $Y2=2.72
r142 33 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.145 $Y2=2.72
r143 31 33 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=7.335 $Y=2.34
+ $X2=7.335 $Y2=2.72
r144 28 47 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.37 $Y2=2.72
r145 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.54 $Y2=2.72
r146 24 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.4 $Y=2.635 $X2=8.4
+ $Y2=2.72
r147 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.4 $Y=2.635
+ $X2=8.4 $Y2=2.34
r148 23 64 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=5.455 $Y2=2.72
r149 22 71 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.205 $Y=2.72
+ $X2=6.395 $Y2=2.72
r150 22 23 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.205 $Y=2.72
+ $X2=5.645 $Y2=2.72
r151 21 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=2.72
+ $X2=4.54 $Y2=2.72
r152 20 64 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.265 $Y=2.72
+ $X2=5.455 $Y2=2.72
r153 20 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.265 $Y=2.72
+ $X2=4.705 $Y2=2.72
r154 16 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.72
r155 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.34
r156 5 26 600 $w=1.7e-07 $l=9.45238e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.485 $X2=8.4 $Y2=2.34
r157 4 31 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=2.34
r158 3 68 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2.34
r159 2 61 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2.34
r160 1 18 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.485 $X2=4.54 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%A_109_47# 1 2 3 4 19 21 24 28 29 35 39 40
+ 45
c94 45 0 1.52763e-19 $X=7.1 $Y=0.825
c95 35 0 1.39973e-19 $X=6.885 $Y=0.85
c96 24 0 7.10587e-20 $X=7.83 $Y=0.675
r97 44 45 11.4037 $w=2.18e-07 $l=2.13e-07 $layer=LI1_cond $X=6.887 $Y=0.825
+ $X2=7.1 $Y2=0.825
r98 39 40 10.6148 $w=2.78e-07 $l=2.15e-07 $layer=LI1_cond $X=1.67 $Y=0.795
+ $X2=1.455 $Y2=0.795
r99 36 44 0.104768 $w=2.18e-07 $l=2e-09 $layer=LI1_cond $X=6.885 $Y=0.825
+ $X2=6.887 $Y2=0.825
r100 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.885 $Y=0.85
+ $X2=6.885 $Y2=0.85
r101 31 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.765 $Y=0.85
+ $X2=1.765 $Y2=0.85
r102 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.91 $Y=0.85
+ $X2=1.765 $Y2=0.85
r103 28 35 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=6.69 $Y=0.85
+ $X2=6.885 $Y2=0.85
r104 28 29 5.91583 $w=1.4e-07 $l=4.78e-06 $layer=MET1_cond $X=6.69 $Y=0.85
+ $X2=1.91 $Y2=0.85
r105 24 26 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.83 $Y=0.675
+ $X2=7.83 $Y2=0.81
r106 21 26 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.745 $Y=0.81
+ $X2=7.83 $Y2=0.81
r107 21 45 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=7.745 $Y=0.81
+ $X2=7.1 $Y2=0.81
r108 17 44 2.10765 $w=1.75e-07 $l=1.1e-07 $layer=LI1_cond $X=6.887 $Y=0.715
+ $X2=6.887 $Y2=0.825
r109 17 19 18.6961 $w=1.73e-07 $l=2.95e-07 $layer=LI1_cond $X=6.887 $Y=0.715
+ $X2=6.887 $Y2=0.42
r110 15 40 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.73 $Y=0.74
+ $X2=1.455 $Y2=0.74
r111 4 24 182 $w=1.7e-07 $l=5.24404e-07 $layer=licon1_NDIFF $count=1 $X=7.645
+ $Y=0.235 $X2=7.83 $Y2=0.675
r112 3 19 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=6.705
+ $Y=0.235 $X2=6.89 $Y2=0.42
r113 2 39 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.74
r114 1 15 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%A_485_47# 1 2 3 4 13 21 23 27 29
r51 25 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.95 $Y=0.655
+ $X2=5.95 $Y2=0.42
r52 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0.74
+ $X2=5.01 $Y2=0.74
r53 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.865 $Y=0.74
+ $X2=5.95 $Y2=0.655
r54 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.865 $Y=0.74
+ $X2=5.095 $Y2=0.74
r55 19 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=0.655
+ $X2=5.01 $Y2=0.74
r56 19 21 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.01 $Y=0.655
+ $X2=5.01 $Y2=0.42
r57 15 18 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.61 $Y=0.74
+ $X2=3.55 $Y2=0.74
r58 13 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.925 $Y=0.74
+ $X2=5.01 $Y2=0.74
r59 13 18 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=4.925 $Y=0.74
+ $X2=3.55 $Y2=0.74
r60 4 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.235 $X2=5.95 $Y2=0.42
r61 3 21 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.42
r62 2 18 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.74
r63 1 15 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_4%VGND 1 2 3 4 5 18 20 22 26 30 34 36 37 39
+ 40 42 43 44 61 62 66 72
r129 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r130 67 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r131 66 69 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=5.455 $Y=0
+ $X2=5.455 $Y2=0.38
r132 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r133 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r134 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r135 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r136 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r137 56 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=6.21
+ $Y2=0
r138 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r139 53 72 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=6.58 $Y=0 $X2=6.392
+ $Y2=0
r140 53 55 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.58 $Y=0 $X2=7.13
+ $Y2=0
r141 52 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r142 51 52 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r143 47 51 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=4.37
+ $Y2=0
r144 44 52 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=4.37
+ $Y2=0
r145 44 47 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r146 42 58 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.235 $Y=0
+ $X2=8.05 $Y2=0
r147 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.235 $Y=0 $X2=8.4
+ $Y2=0
r148 41 61 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.565 $Y=0
+ $X2=8.97 $Y2=0
r149 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.565 $Y=0 $X2=8.4
+ $Y2=0
r150 39 55 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.245 $Y=0
+ $X2=7.13 $Y2=0
r151 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.245 $Y=0 $X2=7.37
+ $Y2=0
r152 38 58 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.495 $Y=0
+ $X2=8.05 $Y2=0
r153 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.495 $Y=0 $X2=7.37
+ $Y2=0
r154 36 51 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.375 $Y=0 $X2=4.37
+ $Y2=0
r155 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.375 $Y=0 $X2=4.54
+ $Y2=0
r156 32 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.4 $Y=0.085 $X2=8.4
+ $Y2=0
r157 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.4 $Y=0.085
+ $X2=8.4 $Y2=0.38
r158 28 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.37 $Y=0.085
+ $X2=7.37 $Y2=0
r159 28 30 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.37 $Y=0.085
+ $X2=7.37 $Y2=0.38
r160 24 72 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=6.392 $Y=0.085
+ $X2=6.392 $Y2=0
r161 24 26 10.4488 $w=3.73e-07 $l=3.4e-07 $layer=LI1_cond $X=6.392 $Y=0.085
+ $X2=6.392 $Y2=0.425
r162 23 66 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.645 $Y=0 $X2=5.455
+ $Y2=0
r163 22 72 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=6.205 $Y=0
+ $X2=6.392 $Y2=0
r164 22 23 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.205 $Y=0
+ $X2=5.645 $Y2=0
r165 21 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=4.54
+ $Y2=0
r166 20 66 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.265 $Y=0 $X2=5.455
+ $Y2=0
r167 20 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.265 $Y=0
+ $X2=4.705 $Y2=0
r168 16 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r169 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.38
r170 5 34 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.235 $X2=8.4 $Y2=0.38
r171 4 30 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.175
+ $Y=0.235 $X2=7.36 $Y2=0.38
r172 3 26 182 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.235 $X2=6.42 $Y2=0.425
r173 2 69 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.235 $X2=5.48 $Y2=0.38
r174 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.415
+ $Y=0.235 $X2=4.54 $Y2=0.38
.ends

