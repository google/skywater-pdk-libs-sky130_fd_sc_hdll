* File: sky130_fd_sc_hdll__mux2_8.pex.spice
* Created: Wed Sep  2 08:34:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%A_79_21# 1 2 3 4 13 15 16 18 19 21 22 24 25
+ 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 58 60 61 70 72
+ 73 74 77 81 83 87 88 89 95 114 116 120
c278 120 0 1.1813e-19 $X=8.26 $Y=0.72
c279 95 0 1.88741e-19 $X=8.235 $Y=0.85
c280 83 0 1.56759e-19 $X=8.15 $Y=0.72
c281 81 0 1.69694e-19 $X=8.81 $Y=1.92
r282 114 115 3.17942 $w=3.79e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.81 $Y2=1.202
r283 111 112 3.17942 $w=3.79e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r284 110 111 56.5937 $w=3.79e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.29 $Y2=1.202
r285 109 110 3.17942 $w=3.79e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r286 108 109 56.5937 $w=3.79e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.82 $Y2=1.202
r287 107 108 3.17942 $w=3.79e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r288 106 107 56.5937 $w=3.79e-07 $l=4.45e-07 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=2.35 $Y2=1.202
r289 105 106 3.17942 $w=3.79e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.202
+ $X2=1.905 $Y2=1.202
r290 104 105 56.5937 $w=3.79e-07 $l=4.45e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.88 $Y2=1.202
r291 103 104 3.17942 $w=3.79e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r292 100 101 3.17942 $w=3.79e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r293 99 100 56.5937 $w=3.79e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.94 $Y2=1.202
r294 98 99 3.17942 $w=3.79e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r295 96 120 6.80989 $w=2.18e-07 $l=1.3e-07 $layer=LI1_cond $X=8.26 $Y=0.85
+ $X2=8.26 $Y2=0.72
r296 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.235 $Y=0.85
+ $X2=8.235 $Y2=0.85
r297 92 116 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.255 $Y=0.85
+ $X2=5.255 $Y2=0.72
r298 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.255 $Y=0.85
+ $X2=5.255 $Y2=0.85
r299 89 91 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.4 $Y=0.85
+ $X2=5.255 $Y2=0.85
r300 88 95 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.09 $Y=0.85
+ $X2=8.235 $Y2=0.85
r301 88 89 3.3292 $w=1.4e-07 $l=2.69e-06 $layer=MET1_cond $X=8.09 $Y=0.85
+ $X2=5.4 $Y2=0.85
r302 83 120 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=8.15 $Y=0.72
+ $X2=8.26 $Y2=0.72
r303 83 85 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.15 $Y=0.72
+ $X2=7.93 $Y2=0.72
r304 79 81 198.332 $w=1.68e-07 $l=3.04e-06 $layer=LI1_cond $X=5.77 $Y=1.92
+ $X2=8.81 $Y2=1.92
r305 77 79 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=3.975 $Y=1.92
+ $X2=5.77 $Y2=1.92
r306 74 76 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=3.975 $Y=0.72
+ $X2=4.94 $Y2=0.72
r307 73 116 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=0.72
+ $X2=5.255 $Y2=0.72
r308 73 76 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.17 $Y=0.72
+ $X2=4.94 $Y2=0.72
r309 72 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.89 $Y=1.835
+ $X2=3.975 $Y2=1.92
r310 71 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.89 $Y=1.245
+ $X2=3.89 $Y2=1.16
r311 71 72 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.89 $Y=1.245
+ $X2=3.89 $Y2=1.835
r312 70 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.89 $Y=1.075
+ $X2=3.89 $Y2=1.16
r313 69 74 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.89 $Y=0.805
+ $X2=3.975 $Y2=0.72
r314 69 70 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.89 $Y=0.805
+ $X2=3.89 $Y2=1.075
r315 68 114 31.1583 $w=3.79e-07 $l=2.45e-07 $layer=POLY_cond $X=3.54 $Y=1.202
+ $X2=3.785 $Y2=1.202
r316 68 112 28.6148 $w=3.79e-07 $l=2.25e-07 $layer=POLY_cond $X=3.54 $Y=1.202
+ $X2=3.315 $Y2=1.202
r317 67 68 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.54
+ $Y=1.16 $X2=3.54 $Y2=1.16
r318 64 103 20.3483 $w=3.79e-07 $l=1.6e-07 $layer=POLY_cond $X=1.25 $Y=1.202
+ $X2=1.41 $Y2=1.202
r319 64 101 36.2454 $w=3.79e-07 $l=2.85e-07 $layer=POLY_cond $X=1.25 $Y=1.202
+ $X2=0.965 $Y2=1.202
r320 63 67 149.401 $w=1.68e-07 $l=2.29e-06 $layer=LI1_cond $X=1.25 $Y=1.16
+ $X2=3.54 $Y2=1.16
r321 63 64 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=1.25
+ $Y=1.16 $X2=1.25 $Y2=1.16
r322 61 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=1.16
+ $X2=3.89 $Y2=1.16
r323 61 67 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.805 $Y=1.16
+ $X2=3.54 $Y2=1.16
r324 58 115 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r325 58 60 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r326 55 114 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r327 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r328 52 112 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r329 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r330 49 111 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r331 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
r332 46 110 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r333 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r334 43 109 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r335 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r336 40 108 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r337 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r338 37 107 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r339 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
r340 34 106 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r341 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r342 31 105 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=1.202
r343 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=0.56
r344 28 104 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r345 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r346 25 103 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r347 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r348 22 101 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r349 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r350 19 100 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r351 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r352 16 99 20.1817 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r353 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r354 13 98 24.5487 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r355 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r356 4 81 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=8.665
+ $Y=1.485 $X2=8.81 $Y2=1.92
r357 3 79 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=5.625
+ $Y=1.485 $X2=5.77 $Y2=1.92
r358 2 85 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=7.745
+ $Y=0.235 $X2=7.93 $Y2=0.72
r359 1 76 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.805
+ $Y=0.235 $X2=4.94 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%S 1 3 4 6 7 9 10 12 13 15 16 18 21 24 25 26
+ 28 31 32 37 43
c148 32 0 1.61039e-19 $X=6.4 $Y=1.53
c149 28 0 1.5381e-19 $X=6.45 $Y=1.16
c150 16 0 1.53048e-19 $X=10.065 $Y=1.41
r151 43 47 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.02 $Y=1.16
+ $X2=10.02 $Y2=1.53
r152 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.15
+ $Y=1.16 $X2=10.15 $Y2=1.16
r153 37 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=1.53
+ $X2=9.89 $Y2=1.53
r154 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.255 $Y=1.53
+ $X2=6.255 $Y2=1.53
r155 32 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.4 $Y=1.53
+ $X2=6.255 $Y2=1.53
r156 31 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.745 $Y=1.53
+ $X2=9.89 $Y2=1.53
r157 31 32 4.13984 $w=1.4e-07 $l=3.345e-06 $layer=MET1_cond $X=9.745 $Y=1.53
+ $X2=6.4 $Y2=1.53
r158 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.16 $X2=6.45 $Y2=1.16
r159 26 35 2.47477 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=6.377 $Y=1.495
+ $X2=6.377 $Y2=1.58
r160 26 28 9.30285 $w=4.13e-07 $l=3.35e-07 $layer=LI1_cond $X=6.377 $Y=1.495
+ $X2=6.377 $Y2=1.16
r161 24 35 6.02678 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=6.17 $Y=1.58
+ $X2=6.377 $Y2=1.58
r162 24 25 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=6.17 $Y=1.58
+ $X2=4.365 $Y2=1.58
r163 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.23
+ $Y=1.16 $X2=4.23 $Y2=1.16
r164 19 25 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.255 $Y=1.495
+ $X2=4.365 $Y2=1.58
r165 19 21 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=4.255 $Y=1.495
+ $X2=4.255 $Y2=1.16
r166 16 42 46.2237 $w=3.35e-07 $l=2.89396e-07 $layer=POLY_cond $X=10.065 $Y=1.41
+ $X2=10.15 $Y2=1.16
r167 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.065 $Y=1.41
+ $X2=10.065 $Y2=1.985
r168 13 42 38.6365 $w=3.35e-07 $l=2.13014e-07 $layer=POLY_cond $X=10.04 $Y=0.995
+ $X2=10.15 $Y2=1.16
r169 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.04 $Y=0.995
+ $X2=10.04 $Y2=0.56
r170 10 29 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=6.5 $Y=0.995
+ $X2=6.475 $Y2=1.16
r171 10 12 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6.5 $Y=0.995
+ $X2=6.5 $Y2=0.555
r172 7 29 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=6.475 $Y=1.41
+ $X2=6.475 $Y2=1.16
r173 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.475 $Y=1.41
+ $X2=6.475 $Y2=1.985
r174 4 22 38.5562 $w=2.99e-07 $l=1.78452e-07 $layer=POLY_cond $X=4.285 $Y=0.995
+ $X2=4.257 $Y2=1.16
r175 4 6 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.285 $Y=0.995
+ $X2=4.285 $Y2=0.555
r176 1 22 47.8775 $w=2.99e-07 $l=2.51496e-07 $layer=POLY_cond $X=4.26 $Y=1.41
+ $X2=4.257 $Y2=1.16
r177 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.26 $Y=1.41
+ $X2=4.26 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%A1 1 3 4 6 7 9 10 12 13 14 19 25 33 36
r96 31 33 4.69045 $w=4.15e-07 $l=3.5e-08 $layer=POLY_cond $X=9.01 $Y=1.202
+ $X2=9.045 $Y2=1.202
r97 31 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.01
+ $Y=1.16 $X2=9.01 $Y2=1.16
r98 28 31 58.2956 $w=4.15e-07 $l=4.35e-07 $layer=POLY_cond $X=8.575 $Y=1.202
+ $X2=9.01 $Y2=1.202
r99 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.79
+ $Y=1.16 $X2=4.79 $Y2=1.16
r100 19 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=1.19
+ $X2=8.97 $Y2=1.19
r101 16 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.775 $Y=1.19
+ $X2=4.775 $Y2=1.19
r102 14 16 0.141131 $w=2.3e-07 $l=1.85e-07 $layer=MET1_cond $X=4.96 $Y=1.19
+ $X2=4.775 $Y2=1.19
r103 13 19 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=8.765 $Y=1.19
+ $X2=8.97 $Y2=1.19
r104 13 14 4.70915 $w=1.4e-07 $l=3.805e-06 $layer=MET1_cond $X=8.765 $Y=1.19
+ $X2=4.96 $Y2=1.19
r105 10 33 22.3416 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.045 $Y=1.41
+ $X2=9.045 $Y2=1.202
r106 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.045 $Y=1.41
+ $X2=9.045 $Y2=1.985
r107 7 28 22.3416 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.575 $Y=1.41
+ $X2=8.575 $Y2=1.202
r108 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.575 $Y=1.41
+ $X2=8.575 $Y2=1.985
r109 4 24 56.9138 $w=3.65e-07 $l=3.6e-07 $layer=POLY_cond $X=5.15 $Y=1.142
+ $X2=4.79 $Y2=1.142
r110 4 6 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=5.15 $Y=0.96 $X2=5.15
+ $Y2=0.555
r111 1 24 9.48563 $w=3.65e-07 $l=6e-08 $layer=POLY_cond $X=4.73 $Y=1.142
+ $X2=4.79 $Y2=1.142
r112 1 3 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.73 $Y=0.96 $X2=4.73
+ $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%A0 1 3 4 6 7 9 10 12 14 17 20 23 24 25 29
+ 35 38 41 43
c120 20 0 3.06871e-19 $X=7.325 $Y=0.73
r121 38 41 0.295498 $w=3.88e-07 $l=1e-08 $layer=LI1_cond $X=6.195 $Y=0.62
+ $X2=6.205 $Y2=0.62
r122 29 43 8.01663 $w=3.88e-07 $l=1.45e-07 $layer=LI1_cond $X=6.245 $Y=0.62
+ $X2=6.39 $Y2=0.62
r123 29 41 1.18199 $w=3.88e-07 $l=4e-08 $layer=LI1_cond $X=6.245 $Y=0.62
+ $X2=6.205 $Y2=0.62
r124 29 38 1.03424 $w=3.88e-07 $l=3.5e-08 $layer=LI1_cond $X=6.16 $Y=0.62
+ $X2=6.195 $Y2=0.62
r125 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.71
+ $Y=1.16 $X2=7.71 $Y2=1.16
r126 25 27 15.443 $w=2.37e-07 $l=3e-07 $layer=LI1_cond $X=7.41 $Y=1.16 $X2=7.71
+ $Y2=1.16
r127 24 29 10.6379 $w=3.88e-07 $l=3.6e-07 $layer=LI1_cond $X=5.8 $Y=0.62
+ $X2=6.16 $Y2=0.62
r128 23 25 2.684 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=0.995
+ $X2=7.41 $Y2=1.16
r129 22 23 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.41 $Y=0.815
+ $X2=7.41 $Y2=0.995
r130 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.325 $Y=0.73
+ $X2=7.41 $Y2=0.815
r131 20 43 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=7.325 $Y=0.73 $X2=6.39
+ $Y2=0.73
r132 18 35 45.5644 $w=4.15e-07 $l=3.4e-07 $layer=POLY_cond $X=5.665 $Y=1.202
+ $X2=6.005 $Y2=1.202
r133 18 32 17.4217 $w=4.15e-07 $l=1.3e-07 $layer=POLY_cond $X=5.665 $Y=1.202
+ $X2=5.535 $Y2=1.202
r134 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.665
+ $Y=1.16 $X2=5.665 $Y2=1.16
r135 15 24 7.70378 $w=2.98e-07 $l=2.43875e-07 $layer=LI1_cond $X=5.69 $Y=0.815
+ $X2=5.8 $Y2=0.62
r136 15 17 18.0724 $w=2.18e-07 $l=3.45e-07 $layer=LI1_cond $X=5.69 $Y=0.815
+ $X2=5.69 $Y2=1.16
r137 12 14 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=8.19 $Y=0.96
+ $X2=8.19 $Y2=0.555
r138 11 28 10.2927 $w=3.65e-07 $l=8.5e-08 $layer=POLY_cond $X=7.745 $Y=1.142
+ $X2=7.66 $Y2=1.142
r139 10 12 33.5422 $w=3.65e-07 $l=2.16273e-07 $layer=POLY_cond $X=8.115 $Y=1.142
+ $X2=8.19 $Y2=0.96
r140 10 11 58.4947 $w=3.65e-07 $l=3.7e-07 $layer=POLY_cond $X=8.115 $Y=1.142
+ $X2=7.745 $Y2=1.142
r141 7 28 23.2495 $w=1.5e-07 $l=1.86933e-07 $layer=POLY_cond $X=7.67 $Y=0.96
+ $X2=7.66 $Y2=1.142
r142 7 9 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=7.67 $Y=0.96 $X2=7.67
+ $Y2=0.555
r143 4 35 22.3416 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.005 $Y=1.41
+ $X2=6.005 $Y2=1.202
r144 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.005 $Y=1.41
+ $X2=6.005 $Y2=1.985
r145 1 32 22.3416 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.535 $Y=1.41
+ $X2=5.535 $Y2=1.202
r146 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.535 $Y=1.41
+ $X2=5.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%A_1369_199# 1 2 7 9 10 12 13 15 16 18 21 24
+ 25 29 33 34 35 36 39 41 43 45
c125 45 0 1.53048e-19 $X=9.525 $Y=1.58
c126 16 0 1.69694e-19 $X=9.515 $Y=1.41
c127 10 0 1.56759e-19 $X=7.035 $Y=0.995
r128 41 47 3.40825 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.3 $Y=2.085
+ $X2=10.3 $Y2=1.94
r129 41 43 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.3 $Y=2.085
+ $X2=10.3 $Y2=2.3
r130 37 39 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=10.3 $Y=0.645
+ $X2=10.3 $Y2=0.46
r131 35 47 3.40825 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=10.215 $Y=2
+ $X2=10.3 $Y2=1.94
r132 35 36 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=10.215 $Y=2
+ $X2=9.635 $Y2=2
r133 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.215 $Y=0.73
+ $X2=10.3 $Y2=0.645
r134 33 34 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=10.215 $Y=0.73
+ $X2=9.635 $Y2=0.73
r135 32 36 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=9.525 $Y=1.915
+ $X2=9.635 $Y2=2
r136 31 45 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=9.525 $Y=1.665
+ $X2=9.525 $Y2=1.58
r137 31 32 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=9.525 $Y=1.665
+ $X2=9.525 $Y2=1.915
r138 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.5
+ $Y=1.16 $X2=9.5 $Y2=1.16
r139 27 45 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=9.525 $Y=1.495
+ $X2=9.525 $Y2=1.58
r140 27 29 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=9.525 $Y=1.495
+ $X2=9.525 $Y2=1.16
r141 26 34 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=9.525 $Y=0.815
+ $X2=9.635 $Y2=0.73
r142 26 29 18.0724 $w=2.18e-07 $l=3.45e-07 $layer=LI1_cond $X=9.525 $Y=0.815
+ $X2=9.525 $Y2=1.16
r143 24 45 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=9.415 $Y=1.58
+ $X2=9.525 $Y2=1.58
r144 24 25 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=9.415 $Y=1.58
+ $X2=7.115 $Y2=1.58
r145 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.98
+ $Y=1.16 $X2=6.98 $Y2=1.16
r146 19 25 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.005 $Y=1.495
+ $X2=7.115 $Y2=1.58
r147 19 21 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=7.005 $Y=1.495
+ $X2=7.005 $Y2=1.16
r148 16 30 48.1208 $w=2.95e-07 $l=2.54951e-07 $layer=POLY_cond $X=9.515 $Y=1.41
+ $X2=9.525 $Y2=1.16
r149 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.515 $Y=1.41
+ $X2=9.515 $Y2=1.985
r150 13 30 38.578 $w=2.95e-07 $l=1.81659e-07 $layer=POLY_cond $X=9.49 $Y=0.995
+ $X2=9.525 $Y2=1.16
r151 13 15 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=9.49 $Y=0.995
+ $X2=9.49 $Y2=0.555
r152 10 22 38.7502 $w=3.47e-07 $l=1.65997e-07 $layer=POLY_cond $X=7.035 $Y=0.995
+ $X2=7.037 $Y2=1.16
r153 10 12 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.035 $Y=0.995
+ $X2=7.035 $Y2=0.555
r154 7 22 45.8462 $w=3.47e-07 $l=2.63154e-07 $layer=POLY_cond $X=7.01 $Y=1.41
+ $X2=7.037 $Y2=1.16
r155 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.01 $Y=1.41
+ $X2=7.01 $Y2=1.985
r156 2 47 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.485 $X2=10.3 $Y2=1.96
r157 2 43 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.485 $X2=10.3 $Y2=2.3
r158 1 39 182 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_NDIFF $count=1 $X=10.115
+ $Y=0.235 $X2=10.3 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 40 43 44
+ 45 47 52 57 62 74 83 84 90 93 96 99 106
r141 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r142 106 109 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=9.855 $Y=2.34
+ $X2=9.855 $Y2=2.72
r143 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r144 99 102 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.995 $Y=2.34
+ $X2=3.995 $Y2=2.72
r145 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r146 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r147 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 84 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=9.89 $Y2=2.72
r149 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r150 81 109 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.045 $Y=2.72
+ $X2=9.855 $Y2=2.72
r151 81 83 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.045 $Y=2.72
+ $X2=10.35 $Y2=2.72
r152 80 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r153 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r154 77 80 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=9.43 $Y2=2.72
r155 76 79 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=7.13 $Y=2.72
+ $X2=9.43 $Y2=2.72
r156 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r157 74 109 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.665 $Y=2.72
+ $X2=9.855 $Y2=2.72
r158 74 79 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.665 $Y=2.72
+ $X2=9.43 $Y2=2.72
r159 73 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r160 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r161 70 73 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.67 $Y2=2.72
r162 70 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r163 69 72 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.67 $Y2=2.72
r164 69 70 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r165 67 102 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=3.995 $Y2=2.72
r166 67 69 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.37 $Y2=2.72
r167 66 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r168 66 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r169 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r170 63 96 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.055 $Y2=2.72
r171 63 65 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.45 $Y2=2.72
r172 62 102 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.995 $Y2=2.72
r173 62 65 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.45 $Y2=2.72
r174 61 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r175 61 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r176 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r177 58 93 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.305 $Y=2.72
+ $X2=2.115 $Y2=2.72
r178 58 60 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.305 $Y=2.72
+ $X2=2.53 $Y2=2.72
r179 57 96 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.055 $Y2=2.72
r180 57 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.53 $Y2=2.72
r181 56 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r182 56 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r183 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r184 53 90 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.175 $Y2=2.72
r185 53 55 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.61 $Y2=2.72
r186 52 93 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.925 $Y=2.72
+ $X2=2.115 $Y2=2.72
r187 52 55 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.925 $Y=2.72
+ $X2=1.61 $Y2=2.72
r188 51 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r189 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r190 48 87 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r191 48 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r192 47 90 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=1.175 $Y2=2.72
r193 47 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=0.69 $Y2=2.72
r194 45 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r195 45 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r196 43 72 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.67 $Y2=2.72
r197 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.76 $Y2=2.72
r198 42 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.845 $Y=2.72
+ $X2=7.13 $Y2=2.72
r199 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=2.72
+ $X2=6.76 $Y2=2.72
r200 38 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=2.635
+ $X2=6.76 $Y2=2.72
r201 38 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.76 $Y=2.635
+ $X2=6.76 $Y2=2.34
r202 34 96 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=2.635
+ $X2=3.055 $Y2=2.72
r203 34 36 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.055 $Y=2.635
+ $X2=3.055 $Y2=2
r204 30 93 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=2.635
+ $X2=2.115 $Y2=2.72
r205 30 32 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.115 $Y=2.635
+ $X2=2.115 $Y2=2
r206 26 90 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=2.635
+ $X2=1.175 $Y2=2.72
r207 26 28 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=1.175 $Y=2.635
+ $X2=1.175 $Y2=2
r208 22 87 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r209 22 24 21.8448 $w=3.33e-07 $l=6.35e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2
r210 7 106 600 $w=1.7e-07 $l=9.60937e-07 $layer=licon1_PDIFF $count=1 $X=9.605
+ $Y=1.485 $X2=9.83 $Y2=2.34
r211 6 40 600 $w=1.7e-07 $l=9.47497e-07 $layer=licon1_PDIFF $count=1 $X=6.565
+ $Y=1.485 $X2=6.76 $Y2=2.34
r212 5 99 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2.34
r213 4 36 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r214 3 32 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r215 2 28 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r216 1 24 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%X 1 2 3 4 5 6 7 8 27 31 33 35 39 43 45 47
+ 51 55 57 59 63 67 70 73 74 75 76 77
r115 71 77 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=0.735 $Y=1.575
+ $X2=0.735 $Y2=1.19
r116 71 72 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=1.575
+ $X2=0.735 $Y2=1.66
r117 69 77 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=0.735 $Y=0.805
+ $X2=0.735 $Y2=1.19
r118 69 70 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.805
+ $X2=0.735 $Y2=0.72
r119 65 67 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.55 $Y=1.745
+ $X2=3.55 $Y2=1.96
r120 61 63 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.55 $Y=0.635
+ $X2=3.55 $Y2=0.46
r121 60 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=1.66
+ $X2=2.61 $Y2=1.66
r122 59 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.465 $Y=1.66
+ $X2=3.55 $Y2=1.745
r123 59 60 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.465 $Y=1.66
+ $X2=2.695 $Y2=1.66
r124 58 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0.72
+ $X2=2.61 $Y2=0.72
r125 57 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.465 $Y=0.72
+ $X2=3.55 $Y2=0.635
r126 57 58 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.465 $Y=0.72
+ $X2=2.695 $Y2=0.72
r127 53 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=1.745
+ $X2=2.61 $Y2=1.66
r128 53 55 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.61 $Y=1.745
+ $X2=2.61 $Y2=1.96
r129 49 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.635
+ $X2=2.61 $Y2=0.72
r130 49 51 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.61 $Y=0.635
+ $X2=2.61 $Y2=0.42
r131 48 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=1.66
+ $X2=1.67 $Y2=1.66
r132 47 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.66
+ $X2=2.61 $Y2=1.66
r133 47 48 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.525 $Y=1.66
+ $X2=1.755 $Y2=1.66
r134 46 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0.72
+ $X2=1.67 $Y2=0.72
r135 45 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0.72
+ $X2=2.61 $Y2=0.72
r136 45 46 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.525 $Y=0.72
+ $X2=1.755 $Y2=0.72
r137 41 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.745
+ $X2=1.67 $Y2=1.66
r138 41 43 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.67 $Y=1.745
+ $X2=1.67 $Y2=1.96
r139 37 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.635
+ $X2=1.67 $Y2=0.72
r140 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.67 $Y=0.635
+ $X2=1.67 $Y2=0.46
r141 36 72 2.53056 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.865 $Y=1.66
+ $X2=0.735 $Y2=1.66
r142 35 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=1.66
+ $X2=1.67 $Y2=1.66
r143 35 36 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.585 $Y=1.66
+ $X2=0.865 $Y2=1.66
r144 34 70 2.53056 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.865 $Y=0.72
+ $X2=0.735 $Y2=0.72
r145 33 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0.72
+ $X2=1.67 $Y2=0.72
r146 33 34 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.585 $Y=0.72
+ $X2=0.865 $Y2=0.72
r147 29 72 3.91525 $w=2.35e-07 $l=9.66954e-08 $layer=LI1_cond $X=0.71 $Y=1.745
+ $X2=0.735 $Y2=1.66
r148 29 31 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=0.71 $Y=1.745
+ $X2=0.71 $Y2=1.96
r149 25 70 3.91525 $w=2.35e-07 $l=9.66954e-08 $layer=LI1_cond $X=0.71 $Y=0.635
+ $X2=0.735 $Y2=0.72
r150 25 27 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=0.71 $Y=0.635
+ $X2=0.71 $Y2=0.42
r151 8 67 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.96
r152 7 55 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.96
r153 6 43 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.96
r154 5 31 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
r155 4 63 182 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.46
r156 3 51 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.42
r157 2 39 182 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.46
r158 1 27 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%A_870_297# 1 2 11
c17 2 0 3.14848e-19 $X=6.095 $Y=1.485
r18 8 11 94.2727 $w=1.68e-07 $l=1.445e-06 $layer=LI1_cond $X=4.795 $Y=2.34
+ $X2=6.24 $Y2=2.34
r19 2 11 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.095
+ $Y=1.485 $X2=6.24 $Y2=2.34
r20 1 8 600 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=4.35
+ $Y=1.485 $X2=4.795 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%A_1420_297# 1 2 11
r17 8 11 132.765 $w=1.68e-07 $l=2.035e-06 $layer=LI1_cond $X=7.245 $Y=2.34
+ $X2=9.28 $Y2=2.34
r18 2 11 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.135
+ $Y=1.485 $X2=9.28 $Y2=2.34
r19 1 8 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=1.485 $X2=7.245 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%VGND 1 2 3 4 5 6 7 22 24 28 30 32 37 42 47
+ 52 57 67 68 75 82 89 96 102 106
r151 106 109 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=9.855 $Y=0
+ $X2=9.855 $Y2=0.38
r152 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r153 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r154 96 99 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.995 $Y=0
+ $X2=3.995 $Y2=0.38
r155 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r156 89 92 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.055 $Y=0
+ $X2=3.055 $Y2=0.38
r157 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r158 82 85 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=2.115 $Y2=0.38
r159 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r160 75 78 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.175 $Y=0
+ $X2=1.175 $Y2=0.38
r161 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r162 68 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=9.89 $Y2=0
r163 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r164 65 106 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.045 $Y=0
+ $X2=9.855 $Y2=0
r165 65 67 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.045 $Y=0
+ $X2=10.35 $Y2=0
r166 64 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r167 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r168 61 64 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=7.13 $Y=0 $X2=9.43
+ $Y2=0
r169 61 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.67 $Y2=0
r170 60 63 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=7.13 $Y=0 $X2=9.43
+ $Y2=0
r171 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r172 58 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.99 $Y=0
+ $X2=6.825 $Y2=0
r173 58 60 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.99 $Y=0 $X2=7.13
+ $Y2=0
r174 57 106 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.855 $Y2=0
r175 57 63 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.43 $Y2=0
r176 56 103 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=6.67 $Y2=0
r177 56 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r178 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r179 53 96 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=3.995
+ $Y2=0
r180 53 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=4.37 $Y2=0
r181 52 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.66 $Y=0
+ $X2=6.825 $Y2=0
r182 52 55 149.401 $w=1.68e-07 $l=2.29e-06 $layer=LI1_cond $X=6.66 $Y=0 $X2=4.37
+ $Y2=0
r183 51 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r184 51 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r185 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r186 48 89 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.055
+ $Y2=0
r187 48 50 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.245 $Y=0
+ $X2=3.45 $Y2=0
r188 47 96 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.995
+ $Y2=0
r189 47 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.805 $Y=0
+ $X2=3.45 $Y2=0
r190 46 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r191 46 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r192 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r193 43 82 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.115
+ $Y2=0
r194 43 45 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.53 $Y2=0
r195 42 89 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=3.055
+ $Y2=0
r196 42 45 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=2.53 $Y2=0
r197 41 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r198 41 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r199 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r200 38 75 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.175
+ $Y2=0
r201 38 40 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r202 37 82 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=2.115
+ $Y2=0
r203 37 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.925 $Y=0
+ $X2=1.61 $Y2=0
r204 36 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r205 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r206 33 71 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r207 33 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r208 32 75 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.175
+ $Y2=0
r209 32 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.69
+ $Y2=0
r210 30 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r211 30 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r212 26 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.825 $Y=0.085
+ $X2=6.825 $Y2=0
r213 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.825 $Y=0.085
+ $X2=6.825 $Y2=0.38
r214 22 71 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r215 22 24 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r216 7 109 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=9.565
+ $Y=0.235 $X2=9.83 $Y2=0.38
r217 6 28 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=6.575
+ $Y=0.235 $X2=6.825 $Y2=0.38
r218 5 99 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.38
r219 4 92 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.38
r220 3 85 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.38
r221 2 78 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.38
r222 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%A_872_47# 1 2 11
r22 8 11 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.52 $Y=0.38 $X2=5.36
+ $Y2=0.38
r23 2 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.225
+ $Y=0.235 $X2=5.36 $Y2=0.38
r24 1 8 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=4.36
+ $Y=0.235 $X2=4.52 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_8%A_1422_47# 1 2 11
r21 8 11 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=7.34 $Y=0.38 $X2=8.4
+ $Y2=0.38
r22 2 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.265
+ $Y=0.235 $X2=8.4 $Y2=0.38
r23 1 8 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=7.11
+ $Y=0.235 $X2=7.34 $Y2=0.38
.ends

