* File: sky130_fd_sc_hdll__nand4bb_1.pxi.spice
* Created: Wed Sep  2 08:39:00 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND4BB_1%B_N N_B_N_M1011_g N_B_N_c_71_n N_B_N_c_72_n
+ N_B_N_M1000_g B_N B_N N_B_N_c_69_n N_B_N_c_70_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_1%B_N
x_PM_SKY130_FD_SC_HDLL__NAND4BB_1%D N_D_c_101_n N_D_M1007_g N_D_c_102_n
+ N_D_M1003_g D PM_SKY130_FD_SC_HDLL__NAND4BB_1%D
x_PM_SKY130_FD_SC_HDLL__NAND4BB_1%C N_C_c_136_n N_C_M1004_g N_C_c_137_n
+ N_C_M1005_g C C PM_SKY130_FD_SC_HDLL__NAND4BB_1%C
x_PM_SKY130_FD_SC_HDLL__NAND4BB_1%A_27_93# N_A_27_93#_M1011_s N_A_27_93#_M1000_s
+ N_A_27_93#_c_170_n N_A_27_93#_M1002_g N_A_27_93#_c_171_n N_A_27_93#_M1009_g
+ N_A_27_93#_c_172_n N_A_27_93#_c_183_n N_A_27_93#_c_193_n N_A_27_93#_c_195_n
+ N_A_27_93#_c_173_n N_A_27_93#_c_174_n N_A_27_93#_c_178_n N_A_27_93#_c_175_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_1%A_27_93#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_1%A_500_21# N_A_500_21#_M1010_d
+ N_A_500_21#_M1008_d N_A_500_21#_c_255_n N_A_500_21#_M1006_g
+ N_A_500_21#_c_260_n N_A_500_21#_M1001_g N_A_500_21#_c_256_n
+ N_A_500_21#_c_262_n N_A_500_21#_c_263_n N_A_500_21#_c_264_n
+ N_A_500_21#_c_257_n N_A_500_21#_c_258_n N_A_500_21#_c_266_n
+ N_A_500_21#_c_259_n PM_SKY130_FD_SC_HDLL__NAND4BB_1%A_500_21#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_1%A_N N_A_N_M1010_g N_A_N_c_326_n N_A_N_c_327_n
+ N_A_N_M1008_g A_N A_N A_N N_A_N_c_325_n PM_SKY130_FD_SC_HDLL__NAND4BB_1%A_N
x_PM_SKY130_FD_SC_HDLL__NAND4BB_1%VPWR N_VPWR_M1000_d N_VPWR_M1005_d
+ N_VPWR_M1001_d N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n
+ VPWR N_VPWR_c_365_n N_VPWR_c_360_n N_VPWR_c_367_n N_VPWR_c_368_n
+ N_VPWR_c_369_n PM_SKY130_FD_SC_HDLL__NAND4BB_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND4BB_1%Y N_Y_M1006_d N_Y_M1003_d N_Y_M1009_d
+ N_Y_c_424_n N_Y_c_453_n N_Y_c_426_n N_Y_c_431_n Y Y Y Y Y N_Y_c_422_n Y
+ PM_SKY130_FD_SC_HDLL__NAND4BB_1%Y
x_PM_SKY130_FD_SC_HDLL__NAND4BB_1%VGND N_VGND_M1011_d N_VGND_M1010_s
+ N_VGND_c_468_n N_VGND_c_469_n VGND N_VGND_c_470_n N_VGND_c_471_n
+ N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_1%VGND
cc_1 VNB B_N 0.00224383f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.105
cc_2 VNB N_B_N_c_69_n 0.0264614f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_3 VNB N_B_N_c_70_n 0.0231421f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=0.995
cc_4 VNB N_D_c_101_n 0.0206618f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_5 VNB N_D_c_102_n 0.0267576f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_6 VNB D 0.00162859f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_7 VNB N_C_c_136_n 0.0172215f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_C_c_137_n 0.0218453f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_9 VNB C 0.00425142f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_10 VNB N_A_27_93#_c_170_n 0.0164519f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_11 VNB N_A_27_93#_c_171_n 0.0217139f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.445
cc_12 VNB N_A_27_93#_c_172_n 0.00692258f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_13 VNB N_A_27_93#_c_173_n 0.00355662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_93#_c_174_n 0.0222415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_93#_c_175_n 0.0187525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_500_21#_c_255_n 0.0200732f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_17 VNB N_A_500_21#_c_256_n 0.00858155f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_18 VNB N_A_500_21#_c_257_n 0.034642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_500_21#_c_258_n 0.0118315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_500_21#_c_259_n 0.0387624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_N_M1010_g 0.0389901f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.675
cc_22 VNB A_N 0.0104844f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.445
cc_23 VNB N_A_N_c_325_n 0.028654f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.325
cc_24 VNB N_VPWR_c_360_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB Y 0.00430886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_422_n 0.00707103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_468_n 0.0100056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_469_n 0.00734388f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_29 VNB N_VGND_c_470_n 0.0580885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_471_n 0.0163091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_472_n 0.232485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_473_n 0.0242936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_474_n 0.00534243f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_B_N_c_71_n 0.0350529f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_35 VPB N_B_N_c_72_n 0.0282632f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_36 VPB B_N 0.00403174f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.105
cc_37 VPB N_B_N_c_69_n 0.00523909f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_38 VPB N_D_c_102_n 0.0298846f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_39 VPB D 2.55023e-19 $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_40 VPB N_C_c_137_n 0.0268996f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_41 VPB C 7.0579e-19 $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_42 VPB N_A_27_93#_c_171_n 0.0254095f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.445
cc_43 VPB N_A_27_93#_c_173_n 5.77489e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_93#_c_178_n 0.0194036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_93#_c_175_n 0.0361352f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_500_21#_c_260_n 0.0190023f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.445
cc_47 VPB N_A_500_21#_c_256_n 0.00769254f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_48 VPB N_A_500_21#_c_262_n 0.0136001f $X=-0.19 $Y=1.305 $X2=0.627 $Y2=1.16
cc_49 VPB N_A_500_21#_c_263_n 0.00245886f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_500_21#_c_264_n 0.0190711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_500_21#_c_257_n 0.0254746f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_500_21#_c_266_n 0.0121661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_500_21#_c_259_n 0.0214201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_N_c_326_n 0.0427239f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_55 VPB N_A_N_c_327_n 0.0313876f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_56 VPB A_N 0.00738658f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.445
cc_57 VPB N_A_N_c_325_n 0.00479329f $X=-0.19 $Y=1.305 $X2=0.562 $Y2=1.325
cc_58 VPB N_VPWR_c_361_n 0.0051226f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_59 VPB N_VPWR_c_362_n 0.00281457f $X=-0.19 $Y=1.305 $X2=0.627 $Y2=1.16
cc_60 VPB N_VPWR_c_363_n 0.0176689f $X=-0.19 $Y=1.305 $X2=0.627 $Y2=1.53
cc_61 VPB N_VPWR_c_364_n 0.00497377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_365_n 0.0170333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_360_n 0.043811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_367_n 0.0244713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_368_n 0.0190428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_369_n 0.0189025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB Y 0.0017729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 N_B_N_c_70_n N_D_c_101_n 0.0148932f $X=0.562 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_69 N_B_N_c_71_n N_D_c_102_n 0.0173606f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_70 N_B_N_c_72_n N_D_c_102_n 0.0105345f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_71 B_N N_D_c_102_n 0.00780538f $X=0.565 $Y=1.105 $X2=0 $Y2=0
cc_72 N_B_N_c_69_n N_D_c_102_n 0.0214792f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_73 B_N D 0.0200067f $X=0.565 $Y=1.105 $X2=0 $Y2=0
cc_74 N_B_N_c_69_n D 2.35237e-19 $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_75 B_N N_A_27_93#_c_172_n 0.0312483f $X=0.565 $Y=1.105 $X2=0 $Y2=0
cc_76 N_B_N_c_69_n N_A_27_93#_c_172_n 0.00478441f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B_N_c_70_n N_A_27_93#_c_172_n 0.0101641f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B_N_c_70_n N_A_27_93#_c_183_n 5.09761e-19 $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_79 N_B_N_c_70_n N_A_27_93#_c_174_n 0.0090214f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B_N_c_72_n N_A_27_93#_c_178_n 0.00745385f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_81 N_B_N_c_72_n N_A_27_93#_c_175_n 5.5452e-19 $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_82 B_N N_A_27_93#_c_175_n 0.0442538f $X=0.565 $Y=1.105 $X2=0 $Y2=0
cc_83 N_B_N_c_70_n N_A_27_93#_c_175_n 0.0276394f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_84 B_N N_VPWR_M1000_d 0.00404667f $X=0.565 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_85 N_B_N_c_71_n N_VPWR_c_361_n 0.00189962f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_86 N_B_N_c_72_n N_VPWR_c_361_n 0.00898196f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_87 B_N N_VPWR_c_361_n 0.0152786f $X=0.565 $Y=1.105 $X2=0 $Y2=0
cc_88 N_B_N_c_69_n N_VPWR_c_361_n 3.3202e-19 $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B_N_c_72_n N_VPWR_c_360_n 0.0133043f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_90 N_B_N_c_72_n N_VPWR_c_367_n 0.0069432f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_91 N_B_N_c_70_n N_VGND_c_468_n 0.00431638f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_92 N_B_N_c_70_n N_VGND_c_472_n 0.00512902f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_93 N_B_N_c_70_n N_VGND_c_473_n 0.00395103f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_94 N_D_c_101_n N_C_c_136_n 0.0229778f $X=1.015 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_95 N_D_c_102_n N_C_c_137_n 0.0427968f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_96 D N_C_c_137_n 7.68782e-19 $X=1.1 $Y=1.105 $X2=0 $Y2=0
cc_97 N_D_c_101_n C 0.00178923f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_98 N_D_c_102_n C 0.00252186f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_99 D C 0.0204004f $X=1.1 $Y=1.105 $X2=0 $Y2=0
cc_100 N_D_c_101_n N_A_27_93#_c_172_n 0.0138756f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_101 N_D_c_102_n N_A_27_93#_c_172_n 0.00349222f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_102 D N_A_27_93#_c_172_n 0.017463f $X=1.1 $Y=1.105 $X2=0 $Y2=0
cc_103 N_D_c_101_n N_A_27_93#_c_183_n 0.00482927f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_104 N_D_c_102_n N_A_27_93#_c_193_n 0.00169961f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_105 D N_A_27_93#_c_193_n 0.00324832f $X=1.1 $Y=1.105 $X2=0 $Y2=0
cc_106 N_D_c_101_n N_A_27_93#_c_195_n 0.00584825f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_107 N_D_c_101_n N_A_27_93#_c_174_n 5.67544e-19 $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_108 N_D_c_102_n N_VPWR_c_361_n 0.013607f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_109 N_D_c_102_n N_VPWR_c_362_n 9.92177e-19 $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_110 N_D_c_102_n N_VPWR_c_363_n 0.0060312f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_111 N_D_c_102_n N_VPWR_c_360_n 0.0103576f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_112 N_D_c_102_n N_Y_c_424_n 0.00351332f $X=1.04 $Y=1.41 $X2=0 $Y2=0
cc_113 D N_Y_c_424_n 0.012395f $X=1.1 $Y=1.105 $X2=0 $Y2=0
cc_114 N_D_c_101_n N_VGND_c_468_n 0.00761434f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_115 N_D_c_101_n N_VGND_c_470_n 0.00421322f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_116 N_D_c_101_n N_VGND_c_472_n 0.00744732f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C_c_136_n N_A_27_93#_c_170_n 0.031128f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_118 C N_A_27_93#_c_170_n 9.20948e-19 $X=1.59 $Y=0.765 $X2=0 $Y2=0
cc_119 N_C_c_137_n N_A_27_93#_c_171_n 0.0451981f $X=1.62 $Y=1.41 $X2=0 $Y2=0
cc_120 C N_A_27_93#_c_171_n 3.66345e-19 $X=1.59 $Y=0.765 $X2=0 $Y2=0
cc_121 N_C_c_136_n N_A_27_93#_c_172_n 0.001278f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_122 C N_A_27_93#_c_172_n 0.00593244f $X=1.59 $Y=0.765 $X2=0 $Y2=0
cc_123 N_C_c_136_n N_A_27_93#_c_183_n 0.00299433f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_124 N_C_c_136_n N_A_27_93#_c_193_n 0.012415f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_125 N_C_c_137_n N_A_27_93#_c_193_n 0.00172794f $X=1.62 $Y=1.41 $X2=0 $Y2=0
cc_126 C N_A_27_93#_c_193_n 0.0127535f $X=1.59 $Y=0.765 $X2=0 $Y2=0
cc_127 N_C_c_136_n N_A_27_93#_c_173_n 4.4173e-19 $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_128 N_C_c_137_n N_A_27_93#_c_173_n 0.00199009f $X=1.62 $Y=1.41 $X2=0 $Y2=0
cc_129 C N_A_27_93#_c_173_n 0.0318251f $X=1.59 $Y=0.765 $X2=0 $Y2=0
cc_130 N_C_c_137_n N_VPWR_c_361_n 0.00103655f $X=1.62 $Y=1.41 $X2=0 $Y2=0
cc_131 N_C_c_137_n N_VPWR_c_362_n 0.0121932f $X=1.62 $Y=1.41 $X2=0 $Y2=0
cc_132 N_C_c_137_n N_VPWR_c_363_n 0.00642146f $X=1.62 $Y=1.41 $X2=0 $Y2=0
cc_133 N_C_c_137_n N_VPWR_c_360_n 0.0110599f $X=1.62 $Y=1.41 $X2=0 $Y2=0
cc_134 N_C_c_137_n N_Y_c_426_n 0.019155f $X=1.62 $Y=1.41 $X2=0 $Y2=0
cc_135 C N_Y_c_426_n 0.0170777f $X=1.59 $Y=0.765 $X2=0 $Y2=0
cc_136 N_C_c_137_n Y 7.85734e-19 $X=1.62 $Y=1.41 $X2=0 $Y2=0
cc_137 N_C_c_136_n N_VGND_c_470_n 0.0037981f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_138 N_C_c_136_n N_VGND_c_472_n 0.00594732f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_139 C A_334_47# 0.00183773f $X=1.59 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_140 N_A_27_93#_c_170_n N_A_500_21#_c_255_n 0.032795f $X=2.095 $Y=0.995 $X2=0
+ $Y2=0
cc_141 N_A_27_93#_c_193_n N_A_500_21#_c_255_n 6.40062e-19 $X=1.99 $Y=0.46 $X2=0
+ $Y2=0
cc_142 N_A_27_93#_c_173_n N_A_500_21#_c_255_n 0.00124105f $X=2.155 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_27_93#_c_171_n N_A_500_21#_c_260_n 0.00888678f $X=2.12 $Y=1.41 $X2=0
+ $Y2=0
cc_144 N_A_27_93#_c_171_n N_A_500_21#_c_259_n 0.0237958f $X=2.12 $Y=1.41 $X2=0
+ $Y2=0
cc_145 N_A_27_93#_c_173_n N_A_500_21#_c_259_n 3.16796e-19 $X=2.155 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_27_93#_c_178_n N_VPWR_c_361_n 0.025525f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_147 N_A_27_93#_c_175_n N_VPWR_c_361_n 0.00809139f $X=0.255 $Y=2.065 $X2=0
+ $Y2=0
cc_148 N_A_27_93#_c_171_n N_VPWR_c_362_n 0.00316312f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_27_93#_M1000_s N_VPWR_c_360_n 0.00217517f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_150 N_A_27_93#_c_171_n N_VPWR_c_360_n 0.0118748f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_27_93#_c_178_n N_VPWR_c_360_n 0.0127747f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_152 N_A_27_93#_c_178_n N_VPWR_c_367_n 0.0214988f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_153 N_A_27_93#_c_171_n N_VPWR_c_368_n 0.00673617f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_27_93#_c_171_n N_Y_c_426_n 0.0144822f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_27_93#_c_173_n N_Y_c_426_n 0.0139622f $X=2.155 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_27_93#_c_171_n N_Y_c_431_n 0.00505905f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_27_93#_c_171_n Y 0.00568733f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_27_93#_c_170_n N_Y_c_422_n 0.00480193f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_27_93#_c_193_n N_Y_c_422_n 0.0168729f $X=1.99 $Y=0.46 $X2=0 $Y2=0
cc_160 N_A_27_93#_c_173_n N_Y_c_422_n 0.0607817f $X=2.155 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_27_93#_c_171_n Y 0.00786995f $X=2.12 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_27_93#_c_173_n Y 0.00279348f $X=2.155 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_27_93#_c_172_n N_VGND_M1011_d 0.00356988f $X=1.05 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_164 N_A_27_93#_c_172_n N_VGND_c_468_n 0.0183225f $X=1.05 $Y=0.81 $X2=0 $Y2=0
cc_165 N_A_27_93#_c_195_n N_VGND_c_468_n 0.014474f $X=1.22 $Y=0.46 $X2=0 $Y2=0
cc_166 N_A_27_93#_c_174_n N_VGND_c_468_n 0.00373046f $X=0.26 $Y=0.61 $X2=0 $Y2=0
cc_167 N_A_27_93#_c_170_n N_VGND_c_470_n 0.0037962f $X=2.095 $Y=0.995 $X2=0
+ $Y2=0
cc_168 N_A_27_93#_c_172_n N_VGND_c_470_n 0.00200003f $X=1.05 $Y=0.81 $X2=0 $Y2=0
cc_169 N_A_27_93#_c_193_n N_VGND_c_470_n 0.0346791f $X=1.99 $Y=0.46 $X2=0 $Y2=0
cc_170 N_A_27_93#_c_195_n N_VGND_c_470_n 0.00572412f $X=1.22 $Y=0.46 $X2=0 $Y2=0
cc_171 N_A_27_93#_c_170_n N_VGND_c_472_n 0.0057355f $X=2.095 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A_27_93#_c_172_n N_VGND_c_472_n 0.0106925f $X=1.05 $Y=0.81 $X2=0 $Y2=0
cc_173 N_A_27_93#_c_193_n N_VGND_c_472_n 0.0343943f $X=1.99 $Y=0.46 $X2=0 $Y2=0
cc_174 N_A_27_93#_c_195_n N_VGND_c_472_n 0.00592206f $X=1.22 $Y=0.46 $X2=0 $Y2=0
cc_175 N_A_27_93#_c_174_n N_VGND_c_472_n 0.0111791f $X=0.26 $Y=0.61 $X2=0 $Y2=0
cc_176 N_A_27_93#_c_172_n N_VGND_c_473_n 0.00273927f $X=1.05 $Y=0.81 $X2=0 $Y2=0
cc_177 N_A_27_93#_c_174_n N_VGND_c_473_n 0.00855792f $X=0.26 $Y=0.61 $X2=0 $Y2=0
cc_178 N_A_27_93#_c_172_n A_218_47# 0.00197881f $X=1.05 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_179 N_A_27_93#_c_183_n A_218_47# 0.00203187f $X=1.135 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_180 N_A_27_93#_c_193_n A_218_47# 0.0105375f $X=1.99 $Y=0.46 $X2=-0.19
+ $Y2=-0.24
cc_181 N_A_27_93#_c_195_n A_218_47# 8.85224e-19 $X=1.22 $Y=0.46 $X2=-0.19
+ $Y2=-0.24
cc_182 N_A_27_93#_c_193_n A_334_47# 0.00974868f $X=1.99 $Y=0.46 $X2=-0.19
+ $Y2=-0.24
cc_183 N_A_27_93#_c_193_n A_434_47# 0.00187059f $X=1.99 $Y=0.46 $X2=-0.19
+ $Y2=-0.24
cc_184 N_A_27_93#_c_173_n A_434_47# 0.00288181f $X=2.155 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_185 N_A_500_21#_c_257_n N_A_N_M1010_g 0.00724859f $X=3.97 $Y=1.835 $X2=0
+ $Y2=0
cc_186 N_A_500_21#_c_258_n N_A_N_M1010_g 0.00634298f $X=3.97 $Y=0.4 $X2=0 $Y2=0
cc_187 N_A_500_21#_c_256_n N_A_N_c_326_n 0.00667543f $X=2.935 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_A_500_21#_c_262_n N_A_N_c_326_n 0.00648827f $X=3.74 $Y=1.92 $X2=0 $Y2=0
cc_189 N_A_500_21#_c_257_n N_A_N_c_326_n 0.00952864f $X=3.97 $Y=1.835 $X2=0
+ $Y2=0
cc_190 N_A_500_21#_c_262_n N_A_N_c_327_n 0.0117093f $X=3.74 $Y=1.92 $X2=0 $Y2=0
cc_191 N_A_500_21#_c_264_n N_A_N_c_327_n 0.00696826f $X=3.825 $Y=2.3 $X2=0 $Y2=0
cc_192 N_A_500_21#_c_255_n A_N 0.00101382f $X=2.575 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_500_21#_c_256_n A_N 0.0507311f $X=2.935 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_500_21#_c_262_n A_N 0.0270371f $X=3.74 $Y=1.92 $X2=0 $Y2=0
cc_195 N_A_500_21#_c_257_n A_N 0.0689268f $X=3.97 $Y=1.835 $X2=0 $Y2=0
cc_196 N_A_500_21#_c_259_n A_N 0.00116266f $X=2.6 $Y=1.202 $X2=0 $Y2=0
cc_197 N_A_500_21#_c_256_n N_A_N_c_325_n 0.00217621f $X=2.935 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A_500_21#_c_262_n N_A_N_c_325_n 8.69584e-19 $X=3.74 $Y=1.92 $X2=0 $Y2=0
cc_199 N_A_500_21#_c_257_n N_A_N_c_325_n 0.00825323f $X=3.97 $Y=1.835 $X2=0
+ $Y2=0
cc_200 N_A_500_21#_c_258_n N_A_N_c_325_n 0.00298101f $X=3.97 $Y=0.4 $X2=0 $Y2=0
cc_201 N_A_500_21#_c_266_n N_A_N_c_325_n 0.00213272f $X=3.897 $Y=1.92 $X2=0
+ $Y2=0
cc_202 N_A_500_21#_c_259_n N_A_N_c_325_n 0.00854921f $X=2.6 $Y=1.202 $X2=0 $Y2=0
cc_203 N_A_500_21#_c_256_n N_VPWR_M1001_d 0.00478544f $X=2.935 $Y=1.16 $X2=0
+ $Y2=0
cc_204 N_A_500_21#_c_263_n N_VPWR_M1001_d 0.00360463f $X=3.125 $Y=1.92 $X2=0
+ $Y2=0
cc_205 N_A_500_21#_c_262_n N_VPWR_c_365_n 0.00310557f $X=3.74 $Y=1.92 $X2=0
+ $Y2=0
cc_206 N_A_500_21#_c_264_n N_VPWR_c_365_n 0.0220212f $X=3.825 $Y=2.3 $X2=0 $Y2=0
cc_207 N_A_500_21#_M1008_d N_VPWR_c_360_n 0.00290256f $X=3.68 $Y=2.065 $X2=0
+ $Y2=0
cc_208 N_A_500_21#_c_260_n N_VPWR_c_360_n 0.00814849f $X=2.6 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_500_21#_c_262_n N_VPWR_c_360_n 0.0065397f $X=3.74 $Y=1.92 $X2=0 $Y2=0
cc_210 N_A_500_21#_c_263_n N_VPWR_c_360_n 0.00120667f $X=3.125 $Y=1.92 $X2=0
+ $Y2=0
cc_211 N_A_500_21#_c_264_n N_VPWR_c_360_n 0.0120431f $X=3.825 $Y=2.3 $X2=0 $Y2=0
cc_212 N_A_500_21#_c_260_n N_VPWR_c_368_n 0.00499348f $X=2.6 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A_500_21#_c_260_n N_VPWR_c_369_n 0.0063669f $X=2.6 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_500_21#_c_262_n N_VPWR_c_369_n 0.0284465f $X=3.74 $Y=1.92 $X2=0 $Y2=0
cc_215 N_A_500_21#_c_263_n N_VPWR_c_369_n 0.0237808f $X=3.125 $Y=1.92 $X2=0
+ $Y2=0
cc_216 N_A_500_21#_c_264_n N_VPWR_c_369_n 0.0194383f $X=3.825 $Y=2.3 $X2=0 $Y2=0
cc_217 N_A_500_21#_c_260_n N_Y_c_431_n 0.012958f $X=2.6 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_500_21#_c_255_n Y 0.00509012f $X=2.575 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_500_21#_c_260_n Y 0.00222052f $X=2.6 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A_500_21#_c_256_n Y 0.0638119f $X=2.935 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_500_21#_c_259_n Y 0.0148681f $X=2.6 $Y=1.202 $X2=0 $Y2=0
cc_222 N_A_500_21#_c_255_n N_Y_c_422_n 0.0132024f $X=2.575 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_500_21#_c_256_n N_Y_c_422_n 0.0128294f $X=2.935 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_500_21#_c_259_n N_Y_c_422_n 0.00796387f $X=2.6 $Y=1.202 $X2=0 $Y2=0
cc_225 N_A_500_21#_c_260_n Y 0.0131494f $X=2.6 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A_500_21#_c_263_n Y 0.0144381f $X=3.125 $Y=1.92 $X2=0 $Y2=0
cc_227 N_A_500_21#_c_255_n N_VGND_c_469_n 0.00216975f $X=2.575 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_500_21#_c_258_n N_VGND_c_469_n 0.0226436f $X=3.97 $Y=0.4 $X2=0 $Y2=0
cc_229 N_A_500_21#_c_255_n N_VGND_c_470_n 0.00357668f $X=2.575 $Y=0.995 $X2=0
+ $Y2=0
cc_230 N_A_500_21#_c_258_n N_VGND_c_471_n 0.0227356f $X=3.97 $Y=0.4 $X2=0 $Y2=0
cc_231 N_A_500_21#_M1010_d N_VGND_c_472_n 0.00329626f $X=3.64 $Y=0.235 $X2=0
+ $Y2=0
cc_232 N_A_500_21#_c_255_n N_VGND_c_472_n 0.00672533f $X=2.575 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_500_21#_c_258_n N_VGND_c_472_n 0.013002f $X=3.97 $Y=0.4 $X2=0 $Y2=0
cc_234 N_A_N_c_327_n N_VPWR_c_365_n 0.00468263f $X=3.59 $Y=1.99 $X2=0 $Y2=0
cc_235 N_A_N_c_327_n N_VPWR_c_360_n 0.00628894f $X=3.59 $Y=1.99 $X2=0 $Y2=0
cc_236 N_A_N_c_327_n N_VPWR_c_369_n 0.0109824f $X=3.59 $Y=1.99 $X2=0 $Y2=0
cc_237 A_N Y 0.00475813f $X=3.46 $Y=0.765 $X2=0 $Y2=0
cc_238 N_A_N_M1010_g N_Y_c_422_n 0.00528968f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_239 A_N N_Y_c_422_n 0.00596729f $X=3.46 $Y=0.765 $X2=0 $Y2=0
cc_240 N_A_N_M1010_g N_VGND_c_469_n 0.0116464f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_241 A_N N_VGND_c_469_n 0.0171518f $X=3.46 $Y=0.765 $X2=0 $Y2=0
cc_242 N_A_N_M1010_g N_VGND_c_471_n 0.00291018f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_243 A_N N_VGND_c_471_n 0.0026424f $X=3.46 $Y=0.765 $X2=0 $Y2=0
cc_244 N_A_N_M1010_g N_VGND_c_472_n 0.00464219f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_245 A_N N_VGND_c_472_n 0.00531656f $X=3.46 $Y=0.765 $X2=0 $Y2=0
cc_246 N_VPWR_c_360_n N_Y_M1003_d 0.00566874f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_247 N_VPWR_c_360_n N_Y_M1009_d 0.00239291f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_248 N_VPWR_c_363_n N_Y_c_453_n 0.0216019f $X=1.695 $Y=2.72 $X2=0 $Y2=0
cc_249 N_VPWR_c_360_n N_Y_c_453_n 0.0126319f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_250 N_VPWR_M1005_d N_Y_c_426_n 0.0089079f $X=1.71 $Y=1.485 $X2=0 $Y2=0
cc_251 N_VPWR_c_362_n N_Y_c_426_n 0.0177842f $X=1.86 $Y=2 $X2=0 $Y2=0
cc_252 N_VPWR_c_360_n N_Y_c_431_n 0.0143952f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_253 N_VPWR_c_368_n N_Y_c_431_n 0.0230589f $X=2.75 $Y=2.49 $X2=0 $Y2=0
cc_254 N_VPWR_c_369_n N_Y_c_431_n 0.0241475f $X=3.52 $Y=2.49 $X2=0 $Y2=0
cc_255 N_VPWR_c_360_n Y 0.00229892f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_256 N_VPWR_c_368_n Y 0.00149185f $X=2.75 $Y=2.49 $X2=0 $Y2=0
cc_257 N_Y_c_422_n N_VGND_c_469_n 0.0234548f $X=2.835 $Y=0.38 $X2=0 $Y2=0
cc_258 N_Y_c_422_n N_VGND_c_470_n 0.036812f $X=2.835 $Y=0.38 $X2=0 $Y2=0
cc_259 N_Y_M1006_d N_VGND_c_472_n 0.00250309f $X=2.65 $Y=0.235 $X2=0 $Y2=0
cc_260 N_Y_c_422_n N_VGND_c_472_n 0.0218303f $X=2.835 $Y=0.38 $X2=0 $Y2=0
cc_261 Y A_434_47# 5.13941e-19 $X=2.535 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_262 N_Y_c_422_n A_434_47# 0.00597507f $X=2.835 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_263 N_VGND_c_472_n A_218_47# 0.00366551f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_264 N_VGND_c_472_n A_334_47# 0.00297453f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_265 N_VGND_c_472_n A_434_47# 0.0086186f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
