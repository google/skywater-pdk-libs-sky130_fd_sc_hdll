* File: sky130_fd_sc_hdll__o21bai_1.spice
* Created: Wed Sep  2 08:44:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21bai_1.pex.spice"
.subckt sky130_fd_sc_hdll__o21bai_1  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1002 N_A_105_352#_M1002_d N_B1_N_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.147 PD=1.37 PS=1.54 NRD=0 NRS=24.276 M=1 R=2.8
+ SA=75000.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_327_47#_M1004_d N_A_105_352#_M1004_g N_Y_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.11375 AS=0.2015 PD=1 PS=1.92 NRD=5.532 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_327_47#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.11375 PD=0.98 PS=1 NRD=0.912 NRS=7.38 M=1 R=4.33333 SA=75000.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_A_327_47#_M1005_d N_A1_M1005_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.10725 PD=1.82 PS=0.98 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_B1_N_M1006_g N_A_105_352#_M1006_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.109644 AS=0.1344 PD=0.84 PS=1.48 NRD=32.8202 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1007 N_Y_M1007_d N_A_105_352#_M1007_g N_VPWR_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.16 AS=0.261056 PD=1.32 PS=2 NRD=6.8753 NRS=13.7703 M=1 R=5.55556
+ SA=90000.5 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1001 A_425_297# N_A2_M1001_g N_Y_M1007_d VPB PHIGHVT L=0.18 W=1 AD=0.14
+ AS=0.16 PD=1.28 PS=1.32 NRD=16.7253 NRS=0.9653 M=1 R=5.55556 SA=90001
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_425_297# VPB PHIGHVT L=0.18 W=1 AD=0.29
+ AS=0.14 PD=2.58 PS=1.28 NRD=0.9653 NRS=16.7253 M=1 R=5.55556 SA=90001.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.778 P=10.41
pX9_noxref noxref_12 Y Y PROBETYPE=1
pX10_noxref noxref_13 A2 A2 PROBETYPE=1
pX11_noxref noxref_14 A1 A1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o21bai_1.pxi.spice"
*
.ends
*
*
