# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a31o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a31o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 1.075000 1.855000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775000 0.735000 2.370000 0.905000 ;
        RECT 0.775000 0.905000 1.255000 1.275000 ;
        RECT 2.185000 0.905000 2.370000 1.075000 ;
        RECT 2.185000 1.075000 2.565000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.525000 1.445000 ;
        RECT 0.145000 1.445000 3.155000 1.615000 ;
        RECT 2.775000 1.075000 3.155000 1.445000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.925000 1.075000 4.455000 1.285000 ;
        RECT 4.215000 0.745000 4.455000 1.075000 ;
    END
  END B1
  PIN VGND
    ANTENNADIFFAREA  1.404000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.760000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.905000 0.655000 6.780000 0.825000 ;
        RECT 4.935000 1.785000 6.780000 1.955000 ;
        RECT 5.045000 1.955000 5.215000 2.465000 ;
        RECT 5.985000 1.955000 6.155000 2.465000 ;
        RECT 6.585000 0.825000 6.780000 1.785000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.175000  1.785000 3.285000 1.955000 ;
      RECT 0.175000  1.955000 0.345000 2.465000 ;
      RECT 0.515000  2.125000 0.895000 2.635000 ;
      RECT 1.115000  1.955000 1.285000 2.465000 ;
      RECT 1.455000  0.395000 2.770000 0.565000 ;
      RECT 1.455000  2.125000 1.835000 2.635000 ;
      RECT 2.055000  1.955000 2.225000 2.465000 ;
      RECT 2.395000  2.125000 2.775000 2.635000 ;
      RECT 2.600000  0.565000 2.770000 0.700000 ;
      RECT 2.600000  0.700000 3.835000 0.805000 ;
      RECT 2.600000  0.805000 3.695000 0.870000 ;
      RECT 2.950000  0.085000 3.285000 0.530000 ;
      RECT 3.115000  1.955000 3.285000 2.295000 ;
      RECT 3.115000  2.295000 4.225000 2.465000 ;
      RECT 3.455000  0.295000 3.835000 0.700000 ;
      RECT 3.455000  0.870000 3.695000 1.455000 ;
      RECT 3.455000  1.455000 4.820000 1.625000 ;
      RECT 3.455000  1.625000 3.835000 2.115000 ;
      RECT 4.055000  1.795000 4.225000 2.295000 ;
      RECT 4.135000  0.085000 4.665000 0.565000 ;
      RECT 4.495000  2.125000 4.825000 2.635000 ;
      RECT 4.650000  0.995000 6.355000 1.325000 ;
      RECT 4.650000  1.325000 4.820000 1.455000 ;
      RECT 5.385000  0.085000 5.765000 0.485000 ;
      RECT 5.385000  2.125000 5.765000 2.635000 ;
      RECT 6.325000  0.085000 6.705000 0.485000 ;
      RECT 6.325000  2.125000 6.705000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31o_4
