* File: sky130_fd_sc_hdll__einvn_8.spice
* Created: Wed Sep  2 08:31:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__einvn_8.pex.spice"
.subckt sky130_fd_sc_hdll__einvn_8  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_TE_B_M1024_g N_A_27_47#_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.2015 PD=1.82 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_235_47#_M1004_d N_A_27_47#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75007.4 A=0.0975 P=1.6 MULT=1
MM1007 N_A_235_47#_M1007_d N_A_27_47#_M1007_g N_VGND_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1008 N_A_235_47#_M1007_d N_A_27_47#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1015 N_A_235_47#_M1015_d N_A_27_47#_M1015_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1018 N_A_235_47#_M1015_d N_A_27_47#_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.1 SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1025 N_A_235_47#_M1025_d N_A_27_47#_M1025_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.6 SB=75005 A=0.0975 P=1.6 MULT=1
MM1028 N_A_235_47#_M1025_d N_A_27_47#_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.108875 PD=0.97 PS=0.985 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1029 N_A_235_47#_M1029_d N_A_27_47#_M1029_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.65 AD=0.10075 AS=0.108875 PD=0.96 PS=0.985 NRD=1.836 NRS=11.076 M=1
+ R=4.33333 SA=75003.5 SB=75004 A=0.0975 P=1.6 MULT=1
MM1009 N_Z_M1009_d N_A_M1009_g N_A_235_47#_M1029_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.10075 PD=0.97 PS=0.96 NRD=8.304 NRS=3.684 M=1 R=4.33333 SA=75004
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1010 N_Z_M1009_d N_A_M1010_g N_A_235_47#_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.5
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1019 N_Z_M1019_d N_A_M1019_g N_A_235_47#_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1020 N_Z_M1019_d N_A_M1020_g N_A_235_47#_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.4
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1021 N_Z_M1021_d N_A_M1021_g N_A_235_47#_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.9
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1022 N_Z_M1021_d N_A_M1022_g N_A_235_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.3
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1030 N_Z_M1030_d N_A_M1030_g N_A_235_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006.8
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1033 N_Z_M1030_d N_A_M1033_g N_A_235_47#_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.182 PD=1.02 PS=1.86 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75007.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_VPWR_M1014_d N_TE_B_M1014_g N_A_27_47#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175206 AS=0.27 PD=1.3866 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.8 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1014_d N_TE_B_M1000_g N_A_222_309#_M1000_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.164694 AS=0.1363 PD=1.3034 PS=1.23 NRD=12.5686 NRS=1.0441 M=1
+ R=5.22222 SA=90000.7 SB=90003.5 A=0.1692 P=2.24 MULT=1
MM1002 N_VPWR_M1002_d N_TE_B_M1002_g N_A_222_309#_M1000_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90001.2 SB=90003 A=0.1692 P=2.24 MULT=1
MM1005 N_VPWR_M1002_d N_TE_B_M1005_g N_A_222_309#_M1005_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90001.6 SB=90002.5 A=0.1692 P=2.24 MULT=1
MM1011 N_VPWR_M1011_d N_TE_B_M1011_g N_A_222_309#_M1005_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90002.1 SB=90002.1 A=0.1692 P=2.24 MULT=1
MM1012 N_VPWR_M1011_d N_TE_B_M1012_g N_A_222_309#_M1012_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90002.6 SB=90001.6 A=0.1692 P=2.24 MULT=1
MM1016 N_VPWR_M1016_d N_TE_B_M1016_g N_A_222_309#_M1012_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90003.1 SB=90001.1 A=0.1692 P=2.24 MULT=1
MM1026 N_VPWR_M1016_d N_TE_B_M1026_g N_A_222_309#_M1026_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90003.5 SB=90000.6 A=0.1692 P=2.24 MULT=1
MM1031 N_VPWR_M1031_d N_TE_B_M1031_g N_A_222_309#_M1026_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.2538 AS=0.1363 PD=2.42 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90004 SB=90000.2 A=0.1692 P=2.24 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g N_A_222_309#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1003 N_Z_M1001_d N_A_M1003_g N_A_222_309#_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1006 N_Z_M1006_d N_A_M1006_g N_A_222_309#_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1013 N_Z_M1006_d N_A_M1013_g N_A_222_309#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1017 N_Z_M1017_d N_A_M1017_g N_A_222_309#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1023 N_Z_M1017_d N_A_M1023_g N_A_222_309#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1027 N_Z_M1027_d N_A_M1027_g N_A_222_309#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1032 N_Z_M1027_d N_A_M1032_g N_A_222_309#_M1032_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX34_noxref VNB VPB NWDIODE A=15.3759 P=22.37
*
.include "sky130_fd_sc_hdll__einvn_8.pxi.spice"
*
.ends
*
*
