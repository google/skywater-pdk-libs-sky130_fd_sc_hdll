* File: sky130_fd_sc_hdll__einvp_4.spice
* Created: Wed Sep  2 08:31:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__einvp_4.pex.spice"
.subckt sky130_fd_sc_hdll__einvp_4  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_TE_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1000 N_A_213_47#_M1000_d N_TE_M1000_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1105 AS=0.104 PD=0.99 PS=0.97 NRD=2.76 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1006 N_A_213_47#_M1000_d N_TE_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1105 AS=0.104 PD=0.99 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1007 N_A_213_47#_M1007_d N_TE_M1007_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_A_213_47#_M1007_d N_TE_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.182 PD=0.97 PS=1.86 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_213_47#_M1001_d N_A_M1001_g N_Z_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1002 N_A_213_47#_M1002_d N_A_M1002_g N_Z_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_213_47#_M1002_d N_A_M1008_g N_Z_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_A_213_47#_M1009_d N_A_M1009_g N_Z_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2145 AS=0.104 PD=1.96 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_TE_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.27 PD=2.54 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A_27_47#_M1003_g N_A_235_309#_M1003_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.2538 PD=1.23 PS=2.42 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90000.2 SB=90003.5 A=0.1692 P=2.24 MULT=1
MM1011 N_VPWR_M1003_d N_A_27_47#_M1011_g N_A_235_309#_M1011_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90000.6 SB=90003.1 A=0.1692 P=2.24 MULT=1
MM1015 N_VPWR_M1015_d N_A_27_47#_M1015_g N_A_235_309#_M1011_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90001.1 SB=90002.6 A=0.1692 P=2.24 MULT=1
MM1016 N_VPWR_M1015_d N_A_27_47#_M1016_g N_A_235_309#_M1016_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.164694 PD=1.23 PS=1.3034 NRD=1.0441 NRS=7.3284 M=1
+ R=5.22222 SA=90001.6 SB=90002.1 A=0.1692 P=2.24 MULT=1
MM1005 N_A_235_309#_M1016_s N_A_M1005_g N_Z_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175206 AS=0.145 PD=1.3866 PS=1.29 NRD=5.8903 NRS=0.9653 M=1 R=5.55556
+ SA=90002 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1012 N_A_235_309#_M1012_d N_A_M1012_g N_Z_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1014 N_A_235_309#_M1012_d N_A_M1014_g N_Z_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.9 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1017 N_A_235_309#_M1017_d N_A_M1017_g N_Z_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.4 SB=90000.2 A=0.18 P=2.36 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.4695 P=15.01
c_44 VNB 0 8.32198e-20 $X=0.15 $Y=-0.085
c_83 VPB 0 1.1096e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__einvp_4.pxi.spice"
*
.ends
*
*
