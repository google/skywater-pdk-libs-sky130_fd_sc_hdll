* File: sky130_fd_sc_hdll__ebufn_4.pex.spice
* Created: Thu Aug 27 19:07:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EBUFN_4%A 1 3 4 6 7 8
c32 1 0 1.8958e-19 $X=0.47 $Y=0.995
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.16 $X2=0.575 $Y2=1.16
r34 8 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.66 $Y=1.53 $X2=0.66
+ $Y2=1.16
r35 7 13 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.66 $Y=0.85 $X2=0.66
+ $Y2=1.16
r36 4 12 46.3664 $w=3.31e-07 $l=2.88097e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.577 $Y2=1.16
r37 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r38 1 12 38.6069 $w=3.31e-07 $l=2.11849e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.577 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_4%TE_B 3 5 7 8 9 10 12 13 15 17 18 20 22 23
+ 25 27 28 29 30 31
c87 31 0 1.8958e-19 $X=1.155 $Y=0.85
r88 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.16 $X2=1.165 $Y2=1.16
r89 34 36 15.0625 $w=3.04e-07 $l=9.5e-08 $layer=POLY_cond $X=1.07 $Y=1.247
+ $X2=1.165 $Y2=1.247
r90 33 34 3.96382 $w=3.04e-07 $l=2.5e-08 $layer=POLY_cond $X=1.045 $Y=1.247
+ $X2=1.07 $Y2=1.247
r91 31 37 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=1.19 $Y=0.85
+ $X2=1.19 $Y2=1.16
r92 25 27 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.47 $Y=1.47
+ $X2=3.47 $Y2=2.015
r93 24 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.09 $Y=1.395 $X2=3
+ $Y2=1.395
r94 23 25 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.38 $Y=1.395
+ $X2=3.47 $Y2=1.47
r95 23 24 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.38 $Y=1.395
+ $X2=3.09 $Y2=1.395
r96 20 30 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3 $Y=1.47 $X2=3
+ $Y2=1.395
r97 20 22 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3 $Y=1.47 $X2=3
+ $Y2=2.015
r98 19 29 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.62 $Y=1.395 $X2=2.53
+ $Y2=1.395
r99 18 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.91 $Y=1.395 $X2=3
+ $Y2=1.395
r100 18 19 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.91 $Y=1.395
+ $X2=2.62 $Y2=1.395
r101 15 29 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.53 $Y=1.47
+ $X2=2.53 $Y2=1.395
r102 15 17 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.53 $Y=1.47
+ $X2=2.53 $Y2=2.015
r103 14 28 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.15 $Y=1.395
+ $X2=2.06 $Y2=1.395
r104 13 29 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.44 $Y=1.395
+ $X2=2.53 $Y2=1.395
r105 13 14 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.44 $Y=1.395
+ $X2=2.15 $Y2=1.395
r106 10 28 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.06 $Y=1.47
+ $X2=2.06 $Y2=1.395
r107 10 12 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.06 $Y=1.47
+ $X2=2.06 $Y2=2.015
r108 9 36 96.4107 $w=3.04e-07 $l=5.9945e-07 $layer=POLY_cond $X=1.695 $Y=1.395
+ $X2=1.165 $Y2=1.247
r109 8 28 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.97 $Y=1.395 $X2=2.06
+ $Y2=1.395
r110 8 9 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=1.97 $Y=1.395
+ $X2=1.695 $Y2=1.395
r111 5 34 15.0262 $w=1.8e-07 $l=1.63e-07 $layer=POLY_cond $X=1.07 $Y=1.41
+ $X2=1.07 $Y2=1.247
r112 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.07 $Y=1.41
+ $X2=1.07 $Y2=1.985
r113 1 33 19.2802 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.045 $Y=1.025
+ $X2=1.045 $Y2=1.247
r114 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.045 $Y=1.025
+ $X2=1.045 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_4%A_224_47# 1 2 7 9 10 11 12 14 15 17 19 20
+ 24 25 26 27 33 36 38 41 48 49 50
c95 50 0 8.82398e-20 $X=3.97 $Y=0.96
r96 49 50 32.0796 $w=3.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.97 $Y=1.035
+ $X2=3.97 $Y2=0.96
r97 42 49 18.2945 $w=3.8e-07 $l=1.25e-07 $layer=POLY_cond $X=3.97 $Y=1.16
+ $X2=3.97 $Y2=1.035
r98 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.945
+ $Y=1.16 $X2=3.945 $Y2=1.16
r99 39 48 1.68792 $w=2.5e-07 $l=1.38e-07 $layer=LI1_cond $X=1.825 $Y=1.15
+ $X2=1.687 $Y2=1.15
r100 39 41 97.7272 $w=2.48e-07 $l=2.12e-06 $layer=LI1_cond $X=1.825 $Y=1.15
+ $X2=3.945 $Y2=1.15
r101 37 48 4.76867 $w=2.75e-07 $l=1.25e-07 $layer=LI1_cond $X=1.687 $Y=1.275
+ $X2=1.687 $Y2=1.15
r102 37 38 13.4102 $w=2.73e-07 $l=3.2e-07 $layer=LI1_cond $X=1.687 $Y=1.275
+ $X2=1.687 $Y2=1.595
r103 36 48 4.76867 $w=2.75e-07 $l=1.25e-07 $layer=LI1_cond $X=1.687 $Y=1.025
+ $X2=1.687 $Y2=1.15
r104 35 36 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=1.687 $Y=0.595
+ $X2=1.687 $Y2=1.025
r105 31 38 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.327 $Y=1.68
+ $X2=1.687 $Y2=1.68
r106 31 33 8.8128 $w=2.53e-07 $l=1.95e-07 $layer=LI1_cond $X=1.327 $Y=1.765
+ $X2=1.327 $Y2=1.96
r107 27 35 6.916 $w=3.4e-07 $l=2.28451e-07 $layer=LI1_cond $X=1.55 $Y=0.425
+ $X2=1.687 $Y2=0.595
r108 27 29 8.30437 $w=3.38e-07 $l=2.45e-07 $layer=LI1_cond $X=1.55 $Y=0.425
+ $X2=1.305 $Y2=0.425
r109 24 50 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.91 $Y=0.56 $X2=3.91
+ $Y2=0.96
r110 21 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.515 $Y=1.035
+ $X2=3.44 $Y2=1.035
r111 20 49 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.78 $Y=1.035
+ $X2=3.97 $Y2=1.035
r112 20 21 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.78 $Y=1.035
+ $X2=3.515 $Y2=1.035
r113 17 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.44 $Y=0.96
+ $X2=3.44 $Y2=1.035
r114 17 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.44 $Y=0.96 $X2=3.44
+ $Y2=0.56
r115 16 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.045 $Y=1.035
+ $X2=2.97 $Y2=1.035
r116 15 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=1.035
+ $X2=3.44 $Y2=1.035
r117 15 16 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.365 $Y=1.035
+ $X2=3.045 $Y2=1.035
r118 12 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.97 $Y=0.96
+ $X2=2.97 $Y2=1.035
r119 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.97 $Y=0.96 $X2=2.97
+ $Y2=0.56
r120 10 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.895 $Y=1.035
+ $X2=2.97 $Y2=1.035
r121 10 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.895 $Y=1.035
+ $X2=2.525 $Y2=1.035
r122 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.45 $Y=0.96
+ $X2=2.525 $Y2=1.035
r123 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.45 $Y=0.96 $X2=2.45
+ $Y2=0.56
r124 2 33 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.16
+ $Y=1.485 $X2=1.305 $Y2=1.96
r125 1 29 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.235 $X2=1.305 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_4%A_27_47# 1 2 9 11 13 16 18 20 23 25 27 28
+ 30 33 35 37 41 50 52 54 56 69 70
r98 70 71 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.885 $Y=1.217
+ $X2=5.91 $Y2=1.217
r99 68 70 16.9511 $w=3.27e-07 $l=1.15e-07 $layer=POLY_cond $X=5.77 $Y=1.217
+ $X2=5.885 $Y2=1.217
r100 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.77
+ $Y=1.16 $X2=5.77 $Y2=1.16
r101 66 68 52.3272 $w=3.27e-07 $l=3.55e-07 $layer=POLY_cond $X=5.415 $Y=1.217
+ $X2=5.77 $Y2=1.217
r102 65 66 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.39 $Y=1.217
+ $X2=5.415 $Y2=1.217
r103 64 65 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=4.945 $Y=1.217
+ $X2=5.39 $Y2=1.217
r104 63 64 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.92 $Y=1.217
+ $X2=4.945 $Y2=1.217
r105 61 63 47.1682 $w=3.27e-07 $l=3.2e-07 $layer=POLY_cond $X=4.6 $Y=1.217
+ $X2=4.92 $Y2=1.217
r106 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.6
+ $Y=1.16 $X2=4.6 $Y2=1.16
r107 59 61 18.4251 $w=3.27e-07 $l=1.25e-07 $layer=POLY_cond $X=4.475 $Y=1.217
+ $X2=4.6 $Y2=1.217
r108 58 59 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.45 $Y=1.217
+ $X2=4.475 $Y2=1.217
r109 55 69 44.9453 $w=2.48e-07 $l=9.75e-07 $layer=LI1_cond $X=4.795 $Y=1.15
+ $X2=5.77 $Y2=1.15
r110 55 62 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=4.795 $Y=1.15
+ $X2=4.6 $Y2=1.15
r111 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.795 $Y=1.19
+ $X2=4.65 $Y2=1.19
r112 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.795 $Y=1.19
+ $X2=4.795 $Y2=1.19
r113 52 56 5.28464 $w=1.4e-07 $l=4.27e-06 $layer=MET1_cond $X=0.38 $Y=1.235
+ $X2=4.65 $Y2=1.235
r114 49 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.235 $Y=1.19
+ $X2=0.38 $Y2=1.19
r115 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.235 $Y=1.19
+ $X2=0.235 $Y2=1.19
r116 45 50 28.1981 $w=2.33e-07 $l=5.75e-07 $layer=LI1_cond $X=0.202 $Y=1.765
+ $X2=0.202 $Y2=1.19
r117 43 50 25.7461 $w=2.33e-07 $l=5.25e-07 $layer=LI1_cond $X=0.202 $Y=0.665
+ $X2=0.202 $Y2=1.19
r118 41 43 9.88221 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.215 $Y=0.445
+ $X2=0.215 $Y2=0.665
r119 35 45 5.89299 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=1.895
+ $X2=0.215 $Y2=1.765
r120 35 37 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.215 $Y=1.895
+ $X2=0.215 $Y2=1.96
r121 31 71 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.91 $Y=1.025
+ $X2=5.91 $Y2=1.217
r122 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.91 $Y=1.025
+ $X2=5.91 $Y2=0.56
r123 28 70 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.885 $Y=1.41
+ $X2=5.885 $Y2=1.217
r124 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.885 $Y=1.41
+ $X2=5.885 $Y2=1.985
r125 25 66 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.415 $Y=1.41
+ $X2=5.415 $Y2=1.217
r126 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.415 $Y=1.41
+ $X2=5.415 $Y2=1.985
r127 21 65 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.39 $Y=1.025
+ $X2=5.39 $Y2=1.217
r128 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.39 $Y=1.025
+ $X2=5.39 $Y2=0.56
r129 18 64 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.945 $Y=1.41
+ $X2=4.945 $Y2=1.217
r130 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.945 $Y=1.41
+ $X2=4.945 $Y2=1.985
r131 14 63 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.92 $Y=1.025
+ $X2=4.92 $Y2=1.217
r132 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.92 $Y=1.025
+ $X2=4.92 $Y2=0.56
r133 11 59 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.475 $Y=1.41
+ $X2=4.475 $Y2=1.217
r134 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.475 $Y=1.41
+ $X2=4.475 $Y2=1.985
r135 7 58 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.45 $Y=1.025
+ $X2=4.45 $Y2=1.217
r136 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.45 $Y=1.025
+ $X2=4.45 $Y2=0.56
r137 2 37 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r138 1 41 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_4%VPWR 1 2 3 12 16 19 22 26 27 28 30 49 50
+ 53
r78 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 49 50 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r80 47 50 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=6.21 $Y2=2.72
r81 46 49 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=6.21 $Y2=2.72
r82 46 47 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 44 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r84 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r85 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r86 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r87 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r88 38 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 37 40 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r90 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r91 35 53 10.8012 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.98 $Y=2.72
+ $X2=0.747 $Y2=2.72
r92 35 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.98 $Y=2.72
+ $X2=1.15 $Y2=2.72
r93 30 53 10.8012 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.747 $Y2=2.72
r94 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 28 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r96 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r97 26 43 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.07 $Y=2.72 $X2=2.99
+ $Y2=2.72
r98 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=2.72
+ $X2=3.235 $Y2=2.72
r99 25 46 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.4 $Y=2.72 $X2=3.45
+ $Y2=2.72
r100 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=2.72
+ $X2=3.235 $Y2=2.72
r101 23 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.46 $Y=2.72
+ $X2=2.99 $Y2=2.72
r102 22 40 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.08 $Y=2.72
+ $X2=2.07 $Y2=2.72
r103 21 23 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.46 $Y2=2.72
r104 21 22 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.08 $Y2=2.72
r105 19 21 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.27 $Y=2.36
+ $X2=2.27 $Y2=2.72
r106 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=2.635
+ $X2=3.235 $Y2=2.72
r107 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.235 $Y=2.635
+ $X2=3.235 $Y2=2.36
r108 10 53 1.88438 $w=4.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=2.635
+ $X2=0.747 $Y2=2.72
r109 10 12 15.8191 $w=4.63e-07 $l=6.15e-07 $layer=LI1_cond $X=0.747 $Y=2.635
+ $X2=0.747 $Y2=2.02
r110 3 16 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.09
+ $Y=1.545 $X2=3.235 $Y2=2.36
r111 2 19 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.15
+ $Y=1.545 $X2=2.295 $Y2=2.36
r112 1 12 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.77 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_4%A_340_309# 1 2 3 4 5 18 22 25 26 30 36
r56 35 36 16.8671 $w=5.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.185 $Y=2.18
+ $X2=3.62 $Y2=2.18
r57 28 30 19.7248 $w=5.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.18 $Y=2.18
+ $X2=6.12 $Y2=2.18
r58 26 35 0.104919 $w=5.68e-07 $l=5e-09 $layer=LI1_cond $X=4.19 $Y=2.18
+ $X2=4.185 $Y2=2.18
r59 26 28 20.774 $w=5.68e-07 $l=9.9e-07 $layer=LI1_cond $X=4.19 $Y=2.18 $X2=5.18
+ $Y2=2.18
r60 25 33 4.99224 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=2 $X2=2.765
+ $Y2=2
r61 25 36 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=2.85 $Y=2 $X2=3.62
+ $Y2=2
r62 20 33 1.63057 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.765 $Y=2.105
+ $X2=2.765 $Y2=2
r63 20 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.765 $Y=2.105
+ $X2=2.765 $Y2=2.3
r64 16 33 60.2606 $w=1.98e-07 $l=9.78e-07 $layer=LI1_cond $X=1.787 $Y=2
+ $X2=2.765 $Y2=2
r65 16 18 9.17251 $w=2.43e-07 $l=1.95e-07 $layer=LI1_cond $X=1.787 $Y=2.105
+ $X2=1.787 $Y2=2.3
r66 5 30 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=5.975
+ $Y=1.485 $X2=6.12 $Y2=2.02
r67 4 28 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=5.035
+ $Y=1.485 $X2=5.18 $Y2=2.02
r68 3 35 150 $w=1.7e-07 $l=8.29156e-07 $layer=licon1_PDIFF $count=4 $X=3.56
+ $Y=1.545 $X2=4.185 $Y2=2.02
r69 2 22 600 $w=1.7e-07 $l=8.24318e-07 $layer=licon1_PDIFF $count=1 $X=2.62
+ $Y=1.545 $X2=2.765 $Y2=2.3
r70 1 18 600 $w=1.7e-07 $l=8.15107e-07 $layer=licon1_PDIFF $count=1 $X=1.7
+ $Y=1.545 $X2=1.825 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_4%Z 1 2 3 4 13 19 20 21 22 23 24 25 26 27 28
+ 41 45 48 51 54 56 62 66 68
c65 13 0 8.82398e-20 $X=6.105 $Y=0.735
r66 64 66 5.14483 $w=2.78e-07 $l=1.25e-07 $layer=LI1_cond $X=5.65 $Y=1.585
+ $X2=5.775 $Y2=1.585
r67 62 64 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.315 $Y=1.585
+ $X2=5.65 $Y2=1.585
r68 54 56 19.962 $w=2.78e-07 $l=4.85e-07 $layer=LI1_cond $X=3.785 $Y=1.585
+ $X2=4.27 $Y2=1.585
r69 27 68 3.48281 $w=2.3e-07 $l=1.2e-07 $layer=LI1_cond $X=6.22 $Y=0.735
+ $X2=6.22 $Y2=0.855
r70 27 28 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.22 $Y=0.895
+ $X2=6.22 $Y2=1.19
r71 27 68 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=6.22 $Y=0.895 $X2=6.22
+ $Y2=0.855
r72 26 41 3.11269 $w=2.8e-07 $l=1.15e-07 $layer=LI1_cond $X=6.22 $Y=1.585
+ $X2=6.105 $Y2=1.585
r73 26 28 9.41096 $w=3.98e-07 $l=2.55e-07 $layer=LI1_cond $X=6.22 $Y=1.445
+ $X2=6.22 $Y2=1.19
r74 25 41 11.936 $w=2.78e-07 $l=2.9e-07 $layer=LI1_cond $X=5.815 $Y=1.585
+ $X2=6.105 $Y2=1.585
r75 25 66 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=5.815 $Y=1.585
+ $X2=5.775 $Y2=1.585
r76 24 62 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=5.305 $Y=1.585
+ $X2=5.315 $Y2=1.585
r77 24 59 24.4894 $w=2.78e-07 $l=5.95e-07 $layer=LI1_cond $X=5.305 $Y=1.585
+ $X2=4.71 $Y2=1.585
r78 23 59 17.4924 $w=2.78e-07 $l=4.25e-07 $layer=LI1_cond $X=4.285 $Y=1.585
+ $X2=4.71 $Y2=1.585
r79 23 56 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=4.285 $Y=1.585
+ $X2=4.27 $Y2=1.585
r80 22 54 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=3.775 $Y=1.585
+ $X2=3.785 $Y2=1.585
r81 22 51 20.7851 $w=2.78e-07 $l=5.05e-07 $layer=LI1_cond $X=3.775 $Y=1.585
+ $X2=3.27 $Y2=1.585
r82 21 51 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=3.265 $Y=1.585
+ $X2=3.27 $Y2=1.585
r83 21 48 20.7851 $w=2.78e-07 $l=5.05e-07 $layer=LI1_cond $X=3.265 $Y=1.585
+ $X2=2.76 $Y2=1.585
r84 20 48 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=2.755 $Y=1.585
+ $X2=2.76 $Y2=1.585
r85 20 45 20.7851 $w=2.78e-07 $l=5.05e-07 $layer=LI1_cond $X=2.755 $Y=1.585
+ $X2=2.25 $Y2=1.585
r86 19 45 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=2.245 $Y=1.585
+ $X2=2.25 $Y2=1.585
r87 15 18 45.1374 $w=2.38e-07 $l=9.4e-07 $layer=LI1_cond $X=4.71 $Y=0.735
+ $X2=5.65 $Y2=0.735
r88 13 27 3.33769 $w=2.4e-07 $l=1.15e-07 $layer=LI1_cond $X=6.105 $Y=0.735
+ $X2=6.22 $Y2=0.735
r89 13 18 21.8484 $w=2.38e-07 $l=4.55e-07 $layer=LI1_cond $X=6.105 $Y=0.735
+ $X2=5.65 $Y2=0.735
r90 4 64 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=1.485 $X2=5.65 $Y2=1.64
r91 3 59 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=4.565
+ $Y=1.485 $X2=4.71 $Y2=1.64
r92 2 18 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=5.465
+ $Y=0.235 $X2=5.65 $Y2=0.76
r93 1 15 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.235 $X2=4.71 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_4%VGND 1 2 3 12 16 18 22 24 26 31 41 42 45
+ 48 51
r79 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r80 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r81 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r82 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r83 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r84 39 42 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.91 $Y=0 $X2=6.21
+ $Y2=0
r85 39 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r86 38 41 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=6.21
+ $Y2=0
r87 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r88 36 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.815 $Y=0 $X2=3.625
+ $Y2=0
r89 36 38 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.815 $Y=0 $X2=3.91
+ $Y2=0
r90 35 49 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r91 35 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r92 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r93 32 45 10.8012 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.747
+ $Y2=0
r94 32 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.15
+ $Y2=0
r95 31 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.685
+ $Y2=0
r96 31 34 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=2.495 $Y=0
+ $X2=1.15 $Y2=0
r97 26 45 10.8012 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.747
+ $Y2=0
r98 26 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r99 24 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r100 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r101 20 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0
r102 20 22 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0.36
r103 19 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.685
+ $Y2=0
r104 18 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.625
+ $Y2=0
r105 18 19 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.435 $Y=0
+ $X2=2.875 $Y2=0
r106 14 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=0.085
+ $X2=2.685 $Y2=0
r107 14 16 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=2.685 $Y=0.085
+ $X2=2.685 $Y2=0.36
r108 10 45 1.88438 $w=4.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=0.085
+ $X2=0.747 $Y2=0
r109 10 12 7.07358 $w=4.63e-07 $l=2.75e-07 $layer=LI1_cond $X=0.747 $Y=0.085
+ $X2=0.747 $Y2=0.36
r110 3 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.65 $Y2=0.36
r111 2 16 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.235 $X2=2.71 $Y2=0.36
r112 1 12 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__EBUFN_4%A_413_47# 1 2 3 4 5 16 19 20 21 24 30 34
+ 36
r62 32 34 54.8708 $w=1.88e-07 $l=9.4e-07 $layer=LI1_cond $X=5.18 $Y=0.35
+ $X2=6.12 $Y2=0.35
r63 30 32 49.9091 $w=1.88e-07 $l=8.55e-07 $layer=LI1_cond $X=4.325 $Y=0.35
+ $X2=5.18 $Y2=0.35
r64 27 29 3.77524 $w=2.88e-07 $l=9.5e-08 $layer=LI1_cond $X=4.18 $Y=0.655
+ $X2=4.18 $Y2=0.56
r65 26 30 7.20849 $w=1.9e-07 $l=1.86548e-07 $layer=LI1_cond $X=4.18 $Y=0.445
+ $X2=4.325 $Y2=0.35
r66 26 29 4.57003 $w=2.88e-07 $l=1.15e-07 $layer=LI1_cond $X=4.18 $Y=0.445
+ $X2=4.18 $Y2=0.56
r67 25 36 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=0.755 $X2=3.18
+ $Y2=0.755
r68 24 27 7.11991 $w=2e-07 $l=1.88481e-07 $layer=LI1_cond $X=4.035 $Y=0.755
+ $X2=4.18 $Y2=0.655
r69 24 25 42.7 $w=1.98e-07 $l=7.7e-07 $layer=LI1_cond $X=4.035 $Y=0.755
+ $X2=3.265 $Y2=0.755
r70 21 36 1.93381 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.18 $Y=0.655 $X2=3.18
+ $Y2=0.755
r71 21 23 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.18 $Y=0.655
+ $X2=3.18 $Y2=0.56
r72 19 36 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.755 $X2=3.18
+ $Y2=0.755
r73 19 20 42.7 $w=1.98e-07 $l=7.7e-07 $layer=LI1_cond $X=3.095 $Y=0.755
+ $X2=2.325 $Y2=0.755
r74 16 20 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.16 $Y=0.655
+ $X2=2.325 $Y2=0.755
r75 16 18 3.51212 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.16 $Y=0.655
+ $X2=2.16 $Y2=0.56
r76 5 34 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.985
+ $Y=0.235 $X2=6.12 $Y2=0.36
r77 4 32 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.995
+ $Y=0.235 $X2=5.18 $Y2=0.36
r78 3 29 182 $w=1.7e-07 $l=4.11096e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.235 $X2=4.18 $Y2=0.56
r79 2 23 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.045
+ $Y=0.235 $X2=3.18 $Y2=0.56
r80 1 18 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.235 $X2=2.19 $Y2=0.56
.ends

