* File: sky130_fd_sc_hdll__nand2b_4.spice
* Created: Thu Aug 27 19:13:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand2b_4.pex.spice"
.subckt sky130_fd_sc_hdll__nand2b_4  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_N_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.2015 PD=1.82 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_225_47#_M1004_d N_A_27_47#_M1004_g N_Y_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1005 N_A_225_47#_M1005_d N_A_27_47#_M1005_g N_Y_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1009 N_A_225_47#_M1005_d N_A_27_47#_M1009_g N_Y_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1014 N_A_225_47#_M1014_d N_A_27_47#_M1014_g N_Y_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.092625 AS=0.104 PD=0.935 PS=0.97 NRD=1.836 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_B_M1000_g N_A_225_47#_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.092625 PD=0.97 PS=0.935 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1000_d N_B_M1001_g N_A_225_47#_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_B_M1007_g N_A_225_47#_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1007_d N_B_M1015_g N_A_225_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.2535 PD=1.02 PS=2.08 NRD=8.304 NRS=19.38 M=1 R=4.33333
+ SA=75003.5 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_A_N_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.27 PD=2.54 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A_27_47#_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.6 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_47#_M1010_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1010_d N_A_27_47#_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1017_d N_A_27_47#_M1017_g N_Y_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1525 AS=0.145 PD=1.305 PS=1.29 NRD=3.9203 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1017_d N_B_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.18 W=1 AD=0.1525
+ AS=0.145 PD=1.305 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_B_M1008_g N_Y_M1002_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.5
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1008_d N_B_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_B_M1016_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1 AD=0.4
+ AS=0.145 PD=2.8 PS=1.29 NRD=22.6353 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.4695 P=15.01
pX19_noxref noxref_10 Y Y PROBETYPE=1
pX20_noxref noxref_11 Y Y PROBETYPE=1
pX21_noxref noxref_12 Y Y PROBETYPE=1
pX22_noxref noxref_13 B B PROBETYPE=1
pX23_noxref noxref_14 N_B_X23_noxref_CONDUCTOR B PROBETYPE=1
pX24_noxref noxref_15 B B PROBETYPE=1
c_44 VNB 0 1.21227e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hdll__nand2b_4.pxi.spice"
*
.ends
*
*
