* File: sky130_fd_sc_hdll__and2_2.spice
* Created: Thu Aug 27 18:56:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and2_2.pex.spice"
.subckt sky130_fd_sc_hdll__and2_2  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1007 A_123_75# N_A_M1007_g N_A_27_75#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1386 PD=0.69 PS=1.5 NRD=22.848 NRS=12.852 M=1 R=2.8 SA=75000.3
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g A_123_75# VNB NSHORT L=0.15 W=0.42
+ AD=0.0960112 AS=0.0567 PD=0.855701 PS=0.69 NRD=48.564 NRS=22.848 M=1 R=2.8
+ SA=75000.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_75#_M1001_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.15925 AS=0.148589 PD=1.14 PS=1.3243 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1001_d N_A_27_75#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.15925 AS=0.221 PD=1.14 PS=1.98 NRD=30.456 NRS=10.152 M=1 R=4.33333
+ SA=75001.5 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_75#_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0609 AS=0.1218 PD=0.71 PS=1.42 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90001.9 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_A_27_75#_M1002_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.102723 AS=0.0609 PD=0.834085 PS=0.71 NRD=59.7895 NRS=2.3443 M=1 R=2.33333
+ SA=90000.7 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1000 N_X_M1000_d N_A_27_75#_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.205 AS=0.244577 PD=1.41 PS=1.98592 NRD=20.685 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1005 N_X_M1000_d N_A_27_75#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.205 AS=0.35 PD=1.41 PS=2.7 NRD=4.9053 NRS=12.7853 M=1 R=5.55556
+ SA=90001.2 SB=90000.3 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hdll__and2_2.pxi.spice"
*
.ends
*
*
