* File: sky130_fd_sc_hdll__a211oi_4.pex.spice
* Created: Wed Sep  2 08:16:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 25 27 28
+ 32 35 48 58
c119 32 0 3.10517e-19 $X=3.76 $Y=1.16
c120 22 0 1.40879e-19 $X=3.785 $Y=1.41
c121 20 0 1.41833e-19 $X=1.46 $Y=0.56
r122 48 49 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.217
+ $X2=1.46 $Y2=1.217
r123 47 58 10.6953 $w=5.88e-07 $l=2.15e-07 $layer=LI1_cond $X=1.32 $Y=1.33
+ $X2=1.535 $Y2=1.33
r124 46 48 16.848 $w=3.29e-07 $l=1.15e-07 $layer=POLY_cond $X=1.32 $Y=1.217
+ $X2=1.435 $Y2=1.217
r125 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.32
+ $Y=1.16 $X2=1.32 $Y2=1.16
r126 44 46 48.3465 $w=3.29e-07 $l=3.3e-07 $layer=POLY_cond $X=0.99 $Y=1.217
+ $X2=1.32 $Y2=1.217
r127 43 44 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.217
+ $X2=0.99 $Y2=1.217
r128 41 43 5.12766 $w=3.29e-07 $l=3.5e-08 $layer=POLY_cond $X=0.93 $Y=1.217
+ $X2=0.965 $Y2=1.217
r129 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.16 $X2=0.93 $Y2=1.16
r130 39 41 60.0669 $w=3.29e-07 $l=4.1e-07 $layer=POLY_cond $X=0.52 $Y=1.217
+ $X2=0.93 $Y2=1.217
r131 38 39 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.217
+ $X2=0.52 $Y2=1.217
r132 35 47 1.88919 $w=7.58e-07 $l=8e-08 $layer=LI1_cond $X=1.24 $Y=1.33 $X2=1.32
+ $Y2=1.33
r133 35 42 4.56132 $w=5.88e-07 $l=2.25e-07 $layer=LI1_cond $X=1.155 $Y=1.33
+ $X2=0.93 $Y2=1.33
r134 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.16 $X2=3.76 $Y2=1.16
r135 30 32 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=3.785 $Y=1.445
+ $X2=3.785 $Y2=1.16
r136 28 30 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=3.595 $Y=1.535
+ $X2=3.785 $Y2=1.445
r137 28 58 126.929 $w=1.78e-07 $l=2.06e-06 $layer=LI1_cond $X=3.595 $Y=1.535
+ $X2=1.535 $Y2=1.535
r138 25 33 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.785 $Y2=1.16
r139 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r140 22 33 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.16
r141 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r142 18 49 21.1507 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.217
r143 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r144 15 48 16.8611 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.217
r145 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r146 11 44 21.1507 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=1.217
r147 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=0.56
r148 8 43 16.8611 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.217
r149 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r150 4 39 21.1507 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=1.217
r151 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=0.56
r152 1 38 16.8611 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.217
r153 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%A1 3 5 7 10 12 14 17 19 21 22 24 27 29 42
+ 43 49
r71 43 44 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.315 $Y=1.217
+ $X2=3.34 $Y2=1.217
r72 42 49 51.1397 $w=2.38e-07 $l=1.065e-06 $layer=LI1_cond $X=3.14 $Y=1.155
+ $X2=2.075 $Y2=1.155
r73 41 43 25.7951 $w=3.27e-07 $l=1.75e-07 $layer=POLY_cond $X=3.14 $Y=1.217
+ $X2=3.315 $Y2=1.217
r74 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.14
+ $Y=1.16 $X2=3.14 $Y2=1.16
r75 39 41 43.4832 $w=3.27e-07 $l=2.95e-07 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=3.14 $Y2=1.217
r76 38 39 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.217
+ $X2=2.845 $Y2=1.217
r77 37 38 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.82 $Y2=1.217
r78 36 37 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r79 34 36 56.0122 $w=3.27e-07 $l=3.8e-07 $layer=POLY_cond $X=1.97 $Y=1.217
+ $X2=2.35 $Y2=1.217
r80 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.97
+ $Y=1.16 $X2=1.97 $Y2=1.16
r81 32 34 9.58104 $w=3.27e-07 $l=6.5e-08 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=1.97 $Y2=1.217
r82 31 32 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.217
+ $X2=1.905 $Y2=1.217
r83 29 49 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=2.07 $Y=1.155
+ $X2=2.075 $Y2=1.155
r84 29 35 4.80185 $w=2.38e-07 $l=1e-07 $layer=LI1_cond $X=2.07 $Y=1.155 $X2=1.97
+ $Y2=1.155
r85 25 44 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.34 $Y=1.025
+ $X2=3.34 $Y2=1.217
r86 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.34 $Y=1.025
+ $X2=3.34 $Y2=0.56
r87 22 43 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r88 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r89 19 39 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r90 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r91 15 38 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=1.217
r92 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=0.56
r93 12 37 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r94 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r95 8 36 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r96 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
r97 5 32 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r98 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r99 1 31 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=1.217
r100 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 27 34 37 38 40 41 43 53 63
c136 63 0 1.7401e-19 $X=4.96 $Y=1.325
c137 38 0 4.54042e-19 $X=4.515 $Y=1.53
c138 37 0 1.74717e-19 $X=7.28 $Y=1.53
c139 19 0 2.07476e-19 $X=7.665 $Y=1.41
c140 13 0 1.85748e-19 $X=5.195 $Y=1.41
c141 4 0 1.17325e-19 $X=4.255 $Y=1.41
r142 53 54 12.9919 $w=3.71e-07 $l=1e-07 $layer=POLY_cond $X=5.195 $Y=1.202
+ $X2=5.295 $Y2=1.202
r143 50 51 11.6927 $w=3.71e-07 $l=9e-08 $layer=POLY_cond $X=4.725 $Y=1.202
+ $X2=4.815 $Y2=1.202
r144 49 63 9.58166 $w=5.78e-07 $l=2.6e-07 $layer=LI1_cond $X=4.7 $Y=1.325
+ $X2=4.96 $Y2=1.325
r145 49 59 6.80527 $w=5.78e-07 $l=3.3e-07 $layer=LI1_cond $X=4.7 $Y=1.325
+ $X2=4.37 $Y2=1.325
r146 48 50 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.202
+ $X2=4.725 $Y2=1.202
r147 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.7
+ $Y=1.16 $X2=4.7 $Y2=1.16
r148 46 48 57.814 $w=3.71e-07 $l=4.45e-07 $layer=POLY_cond $X=4.255 $Y=1.202
+ $X2=4.7 $Y2=1.202
r149 45 46 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.202
+ $X2=4.255 $Y2=1.202
r150 43 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=1.53
+ $X2=4.37 $Y2=1.53
r151 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.425 $Y=1.53
+ $X2=7.425 $Y2=1.53
r152 38 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=1.53
+ $X2=4.37 $Y2=1.53
r153 37 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.28 $Y=1.53
+ $X2=7.425 $Y2=1.53
r154 37 38 3.42202 $w=1.4e-07 $l=2.765e-06 $layer=MET1_cond $X=7.28 $Y=1.53
+ $X2=4.515 $Y2=1.53
r155 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.6
+ $Y=1.16 $X2=7.6 $Y2=1.16
r156 31 41 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=7.405 $Y=1.325
+ $X2=7.405 $Y2=1.53
r157 30 34 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.405 $Y=1.16
+ $X2=7.6 $Y2=1.16
r158 30 31 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=1.16
+ $X2=7.405 $Y2=1.325
r159 28 53 13.6415 $w=3.71e-07 $l=1.05e-07 $layer=POLY_cond $X=5.09 $Y=1.202
+ $X2=5.195 $Y2=1.202
r160 28 51 35.7278 $w=3.71e-07 $l=2.75e-07 $layer=POLY_cond $X=5.09 $Y=1.202
+ $X2=4.815 $Y2=1.202
r161 27 63 6.2424 $w=2.38e-07 $l=1.3e-07 $layer=LI1_cond $X=5.09 $Y=1.155
+ $X2=4.96 $Y2=1.155
r162 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.09
+ $Y=1.16 $X2=5.09 $Y2=1.16
r163 22 35 38.5562 $w=2.99e-07 $l=1.80748e-07 $layer=POLY_cond $X=7.66 $Y=0.995
+ $X2=7.627 $Y2=1.16
r164 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.66 $Y=0.995
+ $X2=7.66 $Y2=0.56
r165 19 35 47.8775 $w=2.99e-07 $l=2.68328e-07 $layer=POLY_cond $X=7.665 $Y=1.41
+ $X2=7.627 $Y2=1.16
r166 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.665 $Y=1.41
+ $X2=7.665 $Y2=1.985
r167 16 54 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.295 $Y=0.995
+ $X2=5.295 $Y2=1.202
r168 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.295 $Y=0.995
+ $X2=5.295 $Y2=0.56
r169 13 53 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.202
r170 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r171 10 51 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=1.202
r172 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=0.56
r173 7 50 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.202
r174 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r175 4 46 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.202
r176 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r177 1 45 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=1.202
r178 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%C1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 27 29 31 43
c88 43 0 1.7401e-19 $X=7.155 $Y=1.202
c89 29 0 2.07476e-19 $X=6.885 $Y=1.16
r90 43 44 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.155 $Y=1.202
+ $X2=7.18 $Y2=1.202
r91 40 41 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=6.655 $Y=1.202
+ $X2=6.71 $Y2=1.202
r92 39 40 54.0622 $w=3.7e-07 $l=4.15e-07 $layer=POLY_cond $X=6.24 $Y=1.202
+ $X2=6.655 $Y2=1.202
r93 38 39 8.46757 $w=3.7e-07 $l=6.5e-08 $layer=POLY_cond $X=6.175 $Y=1.202
+ $X2=6.24 $Y2=1.202
r94 37 38 52.7595 $w=3.7e-07 $l=4.05e-07 $layer=POLY_cond $X=5.77 $Y=1.202
+ $X2=6.175 $Y2=1.202
r95 35 37 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=5.715 $Y=1.202
+ $X2=5.77 $Y2=1.202
r96 33 35 2.60541 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=5.695 $Y=1.202
+ $X2=5.715 $Y2=1.202
r97 31 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.715
+ $Y=1.16 $X2=5.715 $Y2=1.16
r98 30 43 35.173 $w=3.7e-07 $l=2.7e-07 $layer=POLY_cond $X=6.885 $Y=1.202
+ $X2=7.155 $Y2=1.202
r99 30 41 22.7973 $w=3.7e-07 $l=1.75e-07 $layer=POLY_cond $X=6.885 $Y=1.202
+ $X2=6.71 $Y2=1.202
r100 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.885
+ $Y=1.16 $X2=6.885 $Y2=1.16
r101 27 31 55.4613 $w=2.38e-07 $l=1.155e-06 $layer=LI1_cond $X=6.83 $Y=1.155
+ $X2=5.675 $Y2=1.155
r102 27 29 3.26808 $w=2.4e-07 $l=1.1e-07 $layer=LI1_cond $X=6.83 $Y=1.155
+ $X2=6.94 $Y2=1.155
r103 22 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.18 $Y=0.995
+ $X2=7.18 $Y2=1.202
r104 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.18 $Y=0.995
+ $X2=7.18 $Y2=0.56
r105 19 43 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.155 $Y=1.41
+ $X2=7.155 $Y2=1.202
r106 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.155 $Y=1.41
+ $X2=7.155 $Y2=1.985
r107 16 41 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.71 $Y=0.995
+ $X2=6.71 $Y2=1.202
r108 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.71 $Y=0.995
+ $X2=6.71 $Y2=0.56
r109 13 40 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r110 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r111 10 39 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.24 $Y=0.995
+ $X2=6.24 $Y2=1.202
r112 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.24 $Y=0.995
+ $X2=6.24 $Y2=0.56
r113 7 38 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.175 $Y=1.41
+ $X2=6.175 $Y2=1.202
r114 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.175 $Y=1.41
+ $X2=6.175 $Y2=1.985
r115 4 37 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.77 $Y=0.995
+ $X2=5.77 $Y2=1.202
r116 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.77 $Y=0.995
+ $X2=5.77 $Y2=0.56
r117 1 33 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.695 $Y=1.41
+ $X2=5.695 $Y2=1.202
r118 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.695 $Y=1.41
+ $X2=5.695 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%A_27_297# 1 2 3 4 5 6 7 22 24 26 30 32 36
+ 38 42 44 46 47 52 57 59 61
c101 46 0 4.11428e-20 $X=4.02 $Y=2.105
c102 7 0 1.43842e-19 $X=7.755 $Y=1.485
r103 50 52 155.273 $w=2.08e-07 $l=2.94e-06 $layer=LI1_cond $X=4.96 $Y=2.36
+ $X2=7.9 $Y2=2.36
r104 48 65 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=2.36
+ $X2=4.02 $Y2=2.36
r105 48 50 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=4.105 $Y=2.36
+ $X2=4.96 $Y2=2.36
r106 47 65 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.02 $Y=2.255
+ $X2=4.02 $Y2=2.36
r107 46 63 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.02 $Y=2.105
+ $X2=4.02 $Y2=1.95
r108 46 47 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.02 $Y=2.105
+ $X2=4.02 $Y2=2.255
r109 45 61 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=1.95
+ $X2=3.08 $Y2=1.95
r110 44 63 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=1.95
+ $X2=4.02 $Y2=1.95
r111 44 45 28.6252 $w=3.08e-07 $l=7.7e-07 $layer=LI1_cond $X=3.935 $Y=1.95
+ $X2=3.165 $Y2=1.95
r112 40 61 3.57226 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.08 $Y=2.105
+ $X2=3.08 $Y2=1.95
r113 40 42 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.08 $Y=2.105
+ $X2=3.08 $Y2=2.3
r114 39 59 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=1.95
+ $X2=2.14 $Y2=1.95
r115 38 61 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=1.95
+ $X2=3.08 $Y2=1.95
r116 38 39 28.6252 $w=3.08e-07 $l=7.7e-07 $layer=LI1_cond $X=2.995 $Y=1.95
+ $X2=2.225 $Y2=1.95
r117 34 59 3.57226 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.14 $Y=2.105
+ $X2=2.14 $Y2=1.95
r118 34 36 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.14 $Y=2.105
+ $X2=2.14 $Y2=2.3
r119 33 57 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=1.95 $X2=1.2
+ $Y2=1.95
r120 32 59 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.95
+ $X2=2.14 $Y2=1.95
r121 32 33 28.6252 $w=3.08e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=1.95
+ $X2=1.285 $Y2=1.95
r122 28 57 3.44808 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=2.105
+ $X2=1.2 $Y2=1.95
r123 28 30 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.2 $Y=2.105
+ $X2=1.2 $Y2=2.3
r124 27 55 3.17836 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=0.345 $Y=1.94
+ $X2=0.22 $Y2=1.94
r125 26 57 3.14896 $w=3e-07 $l=8.9861e-08 $layer=LI1_cond $X=1.115 $Y=1.94
+ $X2=1.2 $Y2=1.95
r126 26 27 30.5993 $w=2.88e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=1.94
+ $X2=0.345 $Y2=1.94
r127 22 55 3.6869 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=0.22 $Y=2.085
+ $X2=0.22 $Y2=1.94
r128 22 24 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=0.22 $Y=2.085
+ $X2=0.22 $Y2=2.3
r129 7 52 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.755
+ $Y=1.485 $X2=7.9 $Y2=2.34
r130 6 50 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=2.36
r131 5 65 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2.3
r132 5 63 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.96
r133 4 61 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.96
r134 4 42 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2.3
r135 3 59 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.96
r136 3 36 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.3
r137 2 57 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.96
r138 2 30 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.3
r139 1 55 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r140 1 24 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%VPWR 1 2 3 4 13 15 20 25 30 40 41 44 51
+ 58 65
r117 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r118 65 68 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.525 $Y=2.36
+ $X2=3.525 $Y2=2.72
r119 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r120 58 61 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.585 $Y=2.36
+ $X2=2.585 $Y2=2.72
r121 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 51 54 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.645 $Y=2.36
+ $X2=1.645 $Y2=2.72
r123 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 44 47 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=2.34
+ $X2=0.705 $Y2=2.72
r125 40 41 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r126 38 41 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=8.05 $Y2=2.72
r127 38 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r128 37 40 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=8.05 $Y2=2.72
r129 37 38 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r130 35 68 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.525 $Y2=2.72
r131 35 37 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.91 $Y2=2.72
r132 34 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 34 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r134 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r135 31 61 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.585 $Y2=2.72
r136 31 33 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.99 $Y2=2.72
r137 30 68 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=3.525 $Y2=2.72
r138 30 33 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=2.99 $Y2=2.72
r139 29 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r140 29 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r141 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r142 26 54 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=1.645 $Y2=2.72
r143 26 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=2.07 $Y2=2.72
r144 25 61 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.585 $Y2=2.72
r145 25 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.07 $Y2=2.72
r146 24 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r147 24 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r148 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r149 21 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r150 21 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r151 20 54 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.645 $Y2=2.72
r152 20 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r153 15 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r154 15 17 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r155 13 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r156 13 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r157 4 65 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.36
r158 3 58 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.36
r159 2 51 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.36
r160 1 44 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%A_869_297# 1 2 7 13 15
r46 15 17 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=5.295 $Y=1.57
+ $X2=5.295 $Y2=1.935
r47 11 15 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.46 $Y=1.57
+ $X2=5.295 $Y2=1.57
r48 11 13 44.0233 $w=2.48e-07 $l=9.55e-07 $layer=LI1_cond $X=5.46 $Y=1.57
+ $X2=6.415 $Y2=1.57
r49 7 17 1.29116 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.13 $Y=1.935 $X2=5.295
+ $Y2=1.935
r50 7 9 24.5855 $w=2.98e-07 $l=6.4e-07 $layer=LI1_cond $X=5.13 $Y=1.935 $X2=4.49
+ $Y2=1.935
r51 2 13 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=6.265
+ $Y=1.485 $X2=6.415 $Y2=1.61
r52 1 9 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%Y 1 2 3 4 5 6 7 8 25 31 33 37 39 41 49 51
+ 53 59 61 69 71 72 73 77
c136 77 0 1.43842e-19 $X=7.92 $Y=1.495
c137 72 0 1.74717e-19 $X=7.055 $Y=0.74
c138 41 0 1.85748e-19 $X=7.68 $Y=1.975
c139 31 0 1.61114e-19 $X=4.275 $Y=0.78
c140 25 0 1.41833e-19 $X=3.585 $Y=0.77
r141 73 79 2.61642 $w=4.78e-07 $l=1.05e-07 $layer=LI1_cond $X=7.92 $Y=1.87
+ $X2=7.92 $Y2=1.975
r142 73 77 11.9577 $w=4.78e-07 $l=3.75e-07 $layer=LI1_cond $X=7.92 $Y=1.87
+ $X2=7.92 $Y2=1.495
r143 65 66 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=4.46 $Y=0.76
+ $X2=4.46 $Y2=0.78
r144 63 65 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=4.46 $Y=0.74
+ $X2=4.46 $Y2=0.76
r145 61 63 9.96707 $w=3.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.46 $Y=0.42
+ $X2=4.46 $Y2=0.74
r146 57 77 30.2799 $w=2.53e-07 $l=6.7e-07 $layer=LI1_cond $X=8.032 $Y=0.825
+ $X2=8.032 $Y2=1.495
r147 56 72 18.2208 $w=2.08e-07 $l=3.45e-07 $layer=LI1_cond $X=7.4 $Y=0.72
+ $X2=7.055 $Y2=0.72
r148 53 57 6.89985 $w=2.1e-07 $l=1.71651e-07 $layer=LI1_cond $X=7.905 $Y=0.72
+ $X2=8.032 $Y2=0.825
r149 53 56 26.671 $w=2.08e-07 $l=5.05e-07 $layer=LI1_cond $X=7.905 $Y=0.72
+ $X2=7.4 $Y2=0.72
r150 52 71 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=6.535 $Y=0.74
+ $X2=6.45 $Y2=0.74
r151 51 72 6.09095 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.93 $Y=0.74
+ $X2=7.055 $Y2=0.74
r152 51 52 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=6.93 $Y=0.74
+ $X2=6.535 $Y2=0.74
r153 47 71 2.68609 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.45 $Y=0.615
+ $X2=6.45 $Y2=0.74
r154 47 49 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.45 $Y=0.615
+ $X2=6.45 $Y2=0.42
r155 43 46 51.3361 $w=2.18e-07 $l=9.8e-07 $layer=LI1_cond $X=5.935 $Y=1.975
+ $X2=6.915 $Y2=1.975
r156 41 79 5.32182 $w=2.2e-07 $l=2.4e-07 $layer=LI1_cond $X=7.68 $Y=1.975
+ $X2=7.92 $Y2=1.975
r157 41 46 40.0736 $w=2.18e-07 $l=7.65e-07 $layer=LI1_cond $X=7.68 $Y=1.975
+ $X2=6.915 $Y2=1.975
r158 40 69 3.77418 $w=2.45e-07 $l=8.74643e-08 $layer=LI1_cond $X=5.595 $Y=0.745
+ $X2=5.51 $Y2=0.74
r159 39 71 3.77418 $w=2.45e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.365 $Y=0.745
+ $X2=6.45 $Y2=0.74
r160 39 40 36.9742 $w=2.38e-07 $l=7.7e-07 $layer=LI1_cond $X=6.365 $Y=0.745
+ $X2=5.595 $Y2=0.745
r161 35 69 2.68609 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.51 $Y=0.615
+ $X2=5.51 $Y2=0.74
r162 35 37 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.51 $Y=0.615
+ $X2=5.51 $Y2=0.42
r163 34 63 3.03234 $w=2.5e-07 $l=1.85e-07 $layer=LI1_cond $X=4.645 $Y=0.74
+ $X2=4.46 $Y2=0.74
r164 33 69 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=0.74
+ $X2=5.51 $Y2=0.74
r165 33 34 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=5.425 $Y=0.74
+ $X2=4.645 $Y2=0.74
r166 31 66 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.275 $Y=0.78
+ $X2=4.46 $Y2=0.78
r167 31 59 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.275 $Y=0.78
+ $X2=3.68 $Y2=0.78
r168 27 30 54.8708 $w=1.88e-07 $l=9.4e-07 $layer=LI1_cond $X=2.14 $Y=0.77
+ $X2=3.08 $Y2=0.77
r169 25 59 5.69365 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=3.585 $Y=0.77
+ $X2=3.68 $Y2=0.77
r170 25 30 29.4785 $w=1.88e-07 $l=5.05e-07 $layer=LI1_cond $X=3.585 $Y=0.77
+ $X2=3.08 $Y2=0.77
r171 8 46 600 $w=1.7e-07 $l=5.73738e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.915 $Y2=1.98
r172 7 43 600 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.485 $X2=5.935 $Y2=1.98
r173 6 56 182 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_NDIFF $count=1 $X=7.255
+ $Y=0.235 $X2=7.4 $Y2=0.74
r174 5 71 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=6.315
+ $Y=0.235 $X2=6.45 $Y2=0.76
r175 5 49 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.315
+ $Y=0.235 $X2=6.45 $Y2=0.42
r176 4 69 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=5.37
+ $Y=0.235 $X2=5.51 $Y2=0.76
r177 4 37 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.37
+ $Y=0.235 $X2=5.51 $Y2=0.42
r178 3 65 182 $w=1.7e-07 $l=6.19072e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.51 $Y2=0.76
r179 3 61 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.51 $Y2=0.42
r180 2 30 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.76
r181 1 27 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44
+ 47 48 50 51 53 54 56 57 58 60 81 89 92 93
r128 92 95 9.30509 $w=4.72e-07 $l=3.6e-07 $layer=LI1_cond $X=7.972 $Y=0
+ $X2=7.972 $Y2=0.36
r129 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r130 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r131 84 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.05
+ $Y2=0
r132 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r133 81 92 6.79641 $w=1.7e-07 $l=3.07e-07 $layer=LI1_cond $X=7.665 $Y=0
+ $X2=7.972 $Y2=0
r134 81 83 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.665 $Y=0 $X2=7.59
+ $Y2=0
r135 80 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r136 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r137 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r138 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r139 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r140 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r141 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r142 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r143 68 71 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=3.91
+ $Y2=0
r144 68 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r145 67 70 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=3.91
+ $Y2=0
r146 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r147 65 89 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.142 $Y2=0
r148 65 67 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.61 $Y2=0
r149 64 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r150 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r151 61 86 4.49698 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r152 61 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r153 60 89 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1 $Y=0 $X2=1.142
+ $Y2=0
r154 60 63 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.69
+ $Y2=0
r155 58 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r156 58 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r157 56 79 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.67
+ $Y2=0
r158 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.92
+ $Y2=0
r159 55 83 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=7.59 $Y2=0
r160 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.085 $Y=0 $X2=6.92
+ $Y2=0
r161 53 76 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.815 $Y=0 $X2=5.75
+ $Y2=0
r162 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=0 $X2=5.98
+ $Y2=0
r163 52 79 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=6.145 $Y=0
+ $X2=6.67 $Y2=0
r164 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=0 $X2=5.98
+ $Y2=0
r165 50 73 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.865 $Y=0 $X2=4.83
+ $Y2=0
r166 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=0 $X2=5.03
+ $Y2=0
r167 49 76 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.195 $Y=0
+ $X2=5.75 $Y2=0
r168 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.195 $Y=0 $X2=5.03
+ $Y2=0
r169 47 70 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=0 $X2=3.91
+ $Y2=0
r170 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=0 $X2=4.02
+ $Y2=0
r171 46 73 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.105 $Y=0
+ $X2=4.83 $Y2=0
r172 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.02
+ $Y2=0
r173 42 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0
r174 42 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.36
r175 38 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=0.085
+ $X2=5.98 $Y2=0
r176 38 40 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.98 $Y=0.085
+ $X2=5.98 $Y2=0.36
r177 34 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0
r178 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0.36
r179 30 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r180 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.36
r181 26 89 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.142 $Y=0.085
+ $X2=1.142 $Y2=0
r182 26 28 11.1201 $w=2.83e-07 $l=2.75e-07 $layer=LI1_cond $X=1.142 $Y=0.085
+ $X2=1.142 $Y2=0.36
r183 22 86 3.0207 $w=3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.197 $Y2=0
r184 22 24 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.245 $Y2=0.38
r185 7 95 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.735
+ $Y=0.235 $X2=7.88 $Y2=0.36
r186 6 44 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.785
+ $Y=0.235 $X2=6.92 $Y2=0.36
r187 5 40 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.845
+ $Y=0.235 $X2=5.98 $Y2=0.36
r188 4 36 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.235 $X2=5.03 $Y2=0.36
r189 3 32 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.36
r190 2 28 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.36
r191 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_4%A_119_47# 1 2 3 4 13 15 16 21 24
r39 24 26 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=0.72 $Y=0.7 $X2=0.72
+ $Y2=0.78
r40 19 21 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.61 $Y=0.38
+ $X2=3.55 $Y2=0.38
r41 17 29 3.75819 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=1.755 $Y=0.38
+ $X2=1.605 $Y2=0.38
r42 17 19 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=1.755 $Y=0.38
+ $X2=2.61 $Y2=0.38
r43 15 29 3.13183 $w=3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.605 $Y=0.505
+ $X2=1.605 $Y2=0.38
r44 15 16 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=1.605 $Y=0.505
+ $X2=1.605 $Y2=0.695
r45 14 26 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.825 $Y=0.78
+ $X2=0.72 $Y2=0.78
r46 13 16 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.455 $Y=0.78
+ $X2=1.605 $Y2=0.695
r47 13 14 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.455 $Y=0.78
+ $X2=0.825 $Y2=0.78
r48 4 21 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.55 $Y2=0.36
r49 3 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.36
r50 2 29 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.36
r51 1 24 182 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.7
.ends

