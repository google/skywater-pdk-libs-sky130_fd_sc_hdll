* File: sky130_fd_sc_hdll__xor2_2.pxi.spice
* Created: Thu Aug 27 19:29:52 2020
* 
x_PM_SKY130_FD_SC_HDLL__XOR2_2%A N_A_c_104_n N_A_M1002_g N_A_c_113_n N_A_M1001_g
+ N_A_c_114_n N_A_M1013_g N_A_c_105_n N_A_M1015_g N_A_c_115_n N_A_M1018_g
+ N_A_c_106_n N_A_M1003_g N_A_c_107_n N_A_M1007_g N_A_c_116_n N_A_M1019_g
+ N_A_c_117_n N_A_c_108_n N_A_c_109_n N_A_c_110_n N_A_c_137_p N_A_c_119_n
+ N_A_c_120_n A N_A_c_111_n N_A_c_112_n PM_SKY130_FD_SC_HDLL__XOR2_2%A
x_PM_SKY130_FD_SC_HDLL__XOR2_2%B N_B_c_240_n N_B_M1006_g N_B_c_230_n N_B_M1016_g
+ N_B_c_241_n N_B_M1009_g N_B_c_231_n N_B_M1017_g N_B_c_232_n N_B_M1000_g
+ N_B_c_242_n N_B_M1005_g N_B_c_243_n N_B_M1010_g N_B_c_233_n N_B_M1004_g
+ N_B_c_234_n N_B_c_235_n B N_B_c_236_n N_B_c_237_n N_B_c_238_n N_B_c_239_n
+ PM_SKY130_FD_SC_HDLL__XOR2_2%B
x_PM_SKY130_FD_SC_HDLL__XOR2_2%A_112_47# N_A_112_47#_M1002_s N_A_112_47#_M1016_s
+ N_A_112_47#_M1006_s N_A_112_47#_c_346_n N_A_112_47#_M1008_g
+ N_A_112_47#_c_357_n N_A_112_47#_M1011_g N_A_112_47#_c_358_n
+ N_A_112_47#_M1014_g N_A_112_47#_c_347_n N_A_112_47#_M1012_g
+ N_A_112_47#_c_348_n N_A_112_47#_c_349_n N_A_112_47#_c_350_n
+ N_A_112_47#_c_374_n N_A_112_47#_c_360_n N_A_112_47#_c_380_n
+ N_A_112_47#_c_351_n N_A_112_47#_c_384_n N_A_112_47#_c_361_n
+ N_A_112_47#_c_362_n N_A_112_47#_c_363_n N_A_112_47#_c_364_n
+ N_A_112_47#_c_352_n N_A_112_47#_c_353_n N_A_112_47#_c_354_n
+ N_A_112_47#_c_355_n N_A_112_47#_c_397_n N_A_112_47#_c_356_n
+ PM_SKY130_FD_SC_HDLL__XOR2_2%A_112_47#
x_PM_SKY130_FD_SC_HDLL__XOR2_2%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1013_s
+ N_A_27_297#_M1009_d N_A_27_297#_c_519_n N_A_27_297#_c_534_n
+ N_A_27_297#_c_515_n N_A_27_297#_c_511_n N_A_27_297#_c_512_n
+ N_A_27_297#_c_518_n N_A_27_297#_c_542_n PM_SKY130_FD_SC_HDLL__XOR2_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__XOR2_2%VPWR N_VPWR_M1001_d N_VPWR_M1018_s N_VPWR_M1005_s
+ N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_572_n
+ N_VPWR_c_573_n N_VPWR_c_574_n VPWR N_VPWR_c_575_n N_VPWR_c_567_n
+ N_VPWR_c_577_n PM_SKY130_FD_SC_HDLL__XOR2_2%VPWR
x_PM_SKY130_FD_SC_HDLL__XOR2_2%A_510_297# N_A_510_297#_M1018_d
+ N_A_510_297#_M1019_d N_A_510_297#_M1010_d N_A_510_297#_M1011_d
+ N_A_510_297#_M1014_d N_A_510_297#_c_659_n N_A_510_297#_c_657_n
+ N_A_510_297#_c_660_n N_A_510_297#_c_686_n N_A_510_297#_c_670_n
+ N_A_510_297#_c_700_p N_A_510_297#_c_655_n N_A_510_297#_c_673_n
+ N_A_510_297#_c_661_n N_A_510_297#_c_656_n
+ PM_SKY130_FD_SC_HDLL__XOR2_2%A_510_297#
x_PM_SKY130_FD_SC_HDLL__XOR2_2%X N_X_M1000_d N_X_M1008_s N_X_M1011_s N_X_c_707_n
+ N_X_c_702_n N_X_c_703_n N_X_c_704_n N_X_c_705_n N_X_c_706_n N_X_c_709_n X
+ PM_SKY130_FD_SC_HDLL__XOR2_2%X
x_PM_SKY130_FD_SC_HDLL__XOR2_2%VGND N_VGND_M1002_d N_VGND_M1015_d N_VGND_M1017_d
+ N_VGND_M1003_d N_VGND_M1008_d N_VGND_M1012_d N_VGND_c_756_n N_VGND_c_757_n
+ N_VGND_c_758_n N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n
+ N_VGND_c_763_n N_VGND_c_764_n N_VGND_c_765_n N_VGND_c_766_n N_VGND_c_767_n
+ N_VGND_c_768_n N_VGND_c_769_n N_VGND_c_770_n N_VGND_c_771_n VGND
+ N_VGND_c_772_n N_VGND_c_773_n N_VGND_c_774_n PM_SKY130_FD_SC_HDLL__XOR2_2%VGND
x_PM_SKY130_FD_SC_HDLL__XOR2_2%A_510_47# N_A_510_47#_M1003_s N_A_510_47#_M1007_s
+ N_A_510_47#_M1004_s N_A_510_47#_c_858_n N_A_510_47#_c_859_n
+ N_A_510_47#_c_860_n N_A_510_47#_c_868_n N_A_510_47#_c_870_n
+ N_A_510_47#_c_861_n PM_SKY130_FD_SC_HDLL__XOR2_2%A_510_47#
cc_1 VNB N_A_c_104_n 0.0201075f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_2 VNB N_A_c_105_n 0.0173707f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.995
cc_3 VNB N_A_c_106_n 0.0214938f $X=-0.19 $Y=-0.24 $X2=2.935 $Y2=0.995
cc_4 VNB N_A_c_107_n 0.0164529f $X=-0.19 $Y=-0.24 $X2=3.355 $Y2=0.995
cc_5 VNB N_A_c_108_n 0.00102836f $X=-0.19 $Y=-0.24 $X2=1.97 $Y2=1.445
cc_6 VNB N_A_c_109_n 0.00215578f $X=-0.19 $Y=-0.24 $X2=2.08 $Y2=1.175
cc_7 VNB N_A_c_110_n 0.0262632f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.16
cc_8 VNB N_A_c_111_n 0.0401884f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.202
cc_9 VNB N_A_c_112_n 0.0451807f $X=-0.19 $Y=-0.24 $X2=3.355 $Y2=1.202
cc_10 VNB N_B_c_230_n 0.0169508f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.41
cc_11 VNB N_B_c_231_n 0.0220751f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.995
cc_12 VNB N_B_c_232_n 0.0180574f $X=-0.19 $Y=-0.24 $X2=2.91 $Y2=1.41
cc_13 VNB N_B_c_233_n 0.0228549f $X=-0.19 $Y=-0.24 $X2=3.38 $Y2=1.41
cc_14 VNB N_B_c_234_n 0.00325917f $X=-0.19 $Y=-0.24 $X2=0.84 $Y2=1.275
cc_15 VNB N_B_c_235_n 0.00345446f $X=-0.19 $Y=-0.24 $X2=0.84 $Y2=1.445
cc_16 VNB N_B_c_236_n 0.0022807f $X=-0.19 $Y=-0.24 $X2=0.76 $Y2=1.16
cc_17 VNB N_B_c_237_n 0.042456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_c_238_n 0.0049602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B_c_239_n 0.0452299f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.202
cc_20 VNB N_A_112_47#_c_346_n 0.0223892f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.995
cc_21 VNB N_A_112_47#_c_347_n 0.0200686f $X=-0.19 $Y=-0.24 $X2=3.355 $Y2=0.995
cc_22 VNB N_A_112_47#_c_348_n 0.0189611f $X=-0.19 $Y=-0.24 $X2=3.38 $Y2=1.985
cc_23 VNB N_A_112_47#_c_349_n 0.00411695f $X=-0.19 $Y=-0.24 $X2=3.38 $Y2=1.985
cc_24 VNB N_A_112_47#_c_350_n 0.0077223f $X=-0.19 $Y=-0.24 $X2=0.84 $Y2=1.275
cc_25 VNB N_A_112_47#_c_351_n 0.00538563f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.16
cc_26 VNB N_A_112_47#_c_352_n 0.00141513f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.202
cc_27 VNB N_A_112_47#_c_353_n 0.00396224f $X=-0.19 $Y=-0.24 $X2=0.76 $Y2=1.202
cc_28 VNB N_A_112_47#_c_354_n 0.00210839f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.202
cc_29 VNB N_A_112_47#_c_355_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.202
cc_30 VNB N_A_112_47#_c_356_n 0.0448811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_567_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.202
cc_32 VNB N_X_c_702_n 0.0115773f $X=-0.19 $Y=-0.24 $X2=2.935 $Y2=0.995
cc_33 VNB N_X_c_703_n 0.0226893f $X=-0.19 $Y=-0.24 $X2=3.355 $Y2=0.995
cc_34 VNB N_X_c_704_n 0.00232972f $X=-0.19 $Y=-0.24 $X2=3.38 $Y2=1.985
cc_35 VNB N_X_c_705_n 0.016074f $X=-0.19 $Y=-0.24 $X2=0.84 $Y2=1.445
cc_36 VNB N_X_c_706_n 0.00273756f $X=-0.19 $Y=-0.24 $X2=1.97 $Y2=1.275
cc_37 VNB N_VGND_c_756_n 0.0112403f $X=-0.19 $Y=-0.24 $X2=3.355 $Y2=0.995
cc_38 VNB N_VGND_c_757_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=3.355 $Y2=0.56
cc_39 VNB N_VGND_c_758_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=3.38 $Y2=1.985
cc_40 VNB N_VGND_c_759_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=1.97 $Y2=1.275
cc_41 VNB N_VGND_c_760_n 0.0201004f $X=-0.19 $Y=-0.24 $X2=2.08 $Y2=1.175
cc_42 VNB N_VGND_c_761_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_762_n 0.00466605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_763_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=1.53
cc_45 VNB N_VGND_c_764_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.202
cc_46 VNB N_VGND_c_765_n 0.0221187f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.202
cc_47 VNB N_VGND_c_766_n 0.00323927f $X=-0.19 $Y=-0.24 $X2=2.91 $Y2=1.202
cc_48 VNB N_VGND_c_767_n 0.0427069f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.202
cc_49 VNB N_VGND_c_768_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=3.355 $Y2=1.202
cc_50 VNB N_VGND_c_769_n 0.0104908f $X=-0.19 $Y=-0.24 $X2=3.38 $Y2=1.202
cc_51 VNB N_VGND_c_770_n 0.0213436f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.53
cc_52 VNB N_VGND_c_771_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_772_n 0.329657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_773_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_774_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_510_47#_c_858_n 0.00554256f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.56
cc_57 VNB N_A_510_47#_c_859_n 0.00466178f $X=-0.19 $Y=-0.24 $X2=2.91 $Y2=1.985
cc_58 VNB N_A_510_47#_c_860_n 0.00496799f $X=-0.19 $Y=-0.24 $X2=2.91 $Y2=1.985
cc_59 VNB N_A_510_47#_c_861_n 0.00300719f $X=-0.19 $Y=-0.24 $X2=3.38 $Y2=1.41
cc_60 VPB N_A_c_113_n 0.019164f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_61 VPB N_A_c_114_n 0.0158458f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_62 VPB N_A_c_115_n 0.0201091f $X=-0.19 $Y=1.305 $X2=2.91 $Y2=1.41
cc_63 VPB N_A_c_116_n 0.0160057f $X=-0.19 $Y=1.305 $X2=3.38 $Y2=1.41
cc_64 VPB N_A_c_117_n 0.00101245f $X=-0.19 $Y=1.305 $X2=0.84 $Y2=1.445
cc_65 VPB N_A_c_108_n 0.00492902f $X=-0.19 $Y=1.305 $X2=1.97 $Y2=1.445
cc_66 VPB N_A_c_119_n 3.51096e-19 $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.53
cc_67 VPB N_A_c_120_n 0.00447127f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=1.53
cc_68 VPB N_A_c_111_n 0.0210787f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.202
cc_69 VPB N_A_c_112_n 0.0238501f $X=-0.19 $Y=1.305 $X2=3.355 $Y2=1.202
cc_70 VPB N_B_c_240_n 0.0159612f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.995
cc_71 VPB N_B_c_241_n 0.0194034f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_72 VPB N_B_c_242_n 0.0164367f $X=-0.19 $Y=1.305 $X2=2.935 $Y2=0.995
cc_73 VPB N_B_c_243_n 0.0198732f $X=-0.19 $Y=1.305 $X2=3.355 $Y2=0.995
cc_74 VPB N_B_c_235_n 0.00164129f $X=-0.19 $Y=1.305 $X2=0.84 $Y2=1.445
cc_75 VPB N_B_c_237_n 0.0207499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_B_c_239_n 0.0224417f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.202
cc_77 VPB N_A_112_47#_c_357_n 0.0190614f $X=-0.19 $Y=1.305 $X2=2.91 $Y2=1.41
cc_78 VPB N_A_112_47#_c_358_n 0.0191634f $X=-0.19 $Y=1.305 $X2=2.935 $Y2=0.995
cc_79 VPB N_A_112_47#_c_348_n 0.0192451f $X=-0.19 $Y=1.305 $X2=3.38 $Y2=1.985
cc_80 VPB N_A_112_47#_c_360_n 0.00712491f $X=-0.19 $Y=1.305 $X2=1.97 $Y2=1.275
cc_81 VPB N_A_112_47#_c_361_n 0.00463147f $X=-0.19 $Y=1.305 $X2=0.84 $Y2=1.175
cc_82 VPB N_A_112_47#_c_362_n 0.00282909f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=1.53
cc_83 VPB N_A_112_47#_c_363_n 0.0260091f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.445
cc_84 VPB N_A_112_47#_c_364_n 0.0024764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_112_47#_c_352_n 0.0034814f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.202
cc_86 VPB N_A_112_47#_c_356_n 0.0209964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_27_297#_c_511_n 0.0106541f $X=-0.19 $Y=1.305 $X2=2.935 $Y2=0.56
cc_88 VPB N_A_27_297#_c_512_n 0.0078945f $X=-0.19 $Y=1.305 $X2=3.355 $Y2=0.56
cc_89 VPB N_VPWR_c_568_n 0.00516582f $X=-0.19 $Y=1.305 $X2=2.91 $Y2=1.985
cc_90 VPB N_VPWR_c_569_n 0.00516582f $X=-0.19 $Y=1.305 $X2=2.935 $Y2=0.56
cc_91 VPB N_VPWR_c_570_n 0.00547498f $X=-0.19 $Y=1.305 $X2=3.38 $Y2=1.41
cc_92 VPB N_VPWR_c_571_n 0.0539344f $X=-0.19 $Y=1.305 $X2=0.84 $Y2=1.275
cc_93 VPB N_VPWR_c_572_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0.84 $Y2=1.445
cc_94 VPB N_VPWR_c_573_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.97 $Y2=1.445
cc_95 VPB N_VPWR_c_574_n 0.00584025f $X=-0.19 $Y=1.305 $X2=2.08 $Y2=1.175
cc_96 VPB N_VPWR_c_575_n 0.0549976f $X=-0.19 $Y=1.305 $X2=0.76 $Y2=1.202
cc_97 VPB N_VPWR_c_567_n 0.0572496f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.202
cc_98 VPB N_VPWR_c_577_n 0.0240178f $X=-0.19 $Y=1.305 $X2=2.935 $Y2=1.202
cc_99 VPB N_A_510_297#_c_655_n 0.00484902f $X=-0.19 $Y=1.305 $X2=0.76 $Y2=1.16
cc_100 VPB N_A_510_297#_c_656_n 0.0112805f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.202
cc_101 VPB N_X_c_707_n 8.41612e-19 $X=-0.19 $Y=1.305 $X2=2.91 $Y2=1.985
cc_102 VPB N_X_c_703_n 0.0214861f $X=-0.19 $Y=1.305 $X2=3.355 $Y2=0.995
cc_103 VPB N_X_c_709_n 0.00216756f $X=-0.19 $Y=1.305 $X2=2.08 $Y2=1.175
cc_104 N_A_c_114_n N_B_c_240_n 0.0380456f $X=0.98 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_105 N_A_c_108_n N_B_c_240_n 2.00149e-19 $X=1.97 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_106 N_A_c_120_n N_B_c_240_n 0.0117284f $X=1.86 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_107 N_A_c_105_n N_B_c_230_n 0.0213001f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_c_108_n N_B_c_241_n 0.001429f $X=1.97 $Y=1.445 $X2=0 $Y2=0
cc_109 N_A_c_120_n N_B_c_241_n 0.0107114f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_110 N_A_c_107_n N_B_c_232_n 0.0195423f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_c_116_n N_B_c_242_n 0.0229853f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_c_109_n N_B_c_234_n 0.017869f $X=2.08 $Y=1.175 $X2=0 $Y2=0
cc_113 N_A_c_110_n N_B_c_234_n 0.0666593f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_c_120_n N_B_c_234_n 0.00664233f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_115 N_A_c_117_n N_B_c_235_n 0.00133759f $X=0.84 $Y=1.445 $X2=0 $Y2=0
cc_116 N_A_c_108_n N_B_c_235_n 8.95935e-19 $X=1.97 $Y=1.445 $X2=0 $Y2=0
cc_117 N_A_c_109_n N_B_c_235_n 2.40733e-19 $X=2.08 $Y=1.175 $X2=0 $Y2=0
cc_118 N_A_c_137_p N_B_c_235_n 0.00639936f $X=0.84 $Y=1.175 $X2=0 $Y2=0
cc_119 N_A_c_120_n N_B_c_235_n 0.00822845f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_120 N_A_c_111_n N_B_c_235_n 0.00484195f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_121 N_A_c_110_n B 4.35466e-19 $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_c_109_n N_B_c_236_n 0.0139407f $X=2.08 $Y=1.175 $X2=0 $Y2=0
cc_123 N_A_c_137_p N_B_c_236_n 0.0102308f $X=0.84 $Y=1.175 $X2=0 $Y2=0
cc_124 N_A_c_120_n N_B_c_236_n 0.0349962f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_125 N_A_c_111_n N_B_c_236_n 0.00173823f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_126 N_A_c_117_n N_B_c_237_n 6.48439e-19 $X=0.84 $Y=1.445 $X2=0 $Y2=0
cc_127 N_A_c_108_n N_B_c_237_n 0.00737674f $X=1.97 $Y=1.445 $X2=0 $Y2=0
cc_128 N_A_c_109_n N_B_c_237_n 0.0179937f $X=2.08 $Y=1.175 $X2=0 $Y2=0
cc_129 N_A_c_120_n N_B_c_237_n 0.00868529f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_130 N_A_c_111_n N_B_c_237_n 0.0226456f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_131 N_A_c_110_n N_B_c_238_n 0.0138657f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_c_112_n N_B_c_238_n 5.94012e-19 $X=3.355 $Y=1.202 $X2=0 $Y2=0
cc_133 N_A_c_110_n N_B_c_239_n 5.93964e-19 $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_c_112_n N_B_c_239_n 0.0244332f $X=3.355 $Y=1.202 $X2=0 $Y2=0
cc_135 N_A_c_120_n N_A_112_47#_M1006_s 0.00187091f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_136 N_A_c_104_n N_A_112_47#_c_348_n 0.0161028f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_113_n N_A_112_47#_c_348_n 0.0111176f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_117_n N_A_112_47#_c_348_n 0.00613788f $X=0.84 $Y=1.445 $X2=0 $Y2=0
cc_139 N_A_c_137_p N_A_112_47#_c_348_n 0.0111408f $X=0.84 $Y=1.175 $X2=0 $Y2=0
cc_140 N_A_c_119_n N_A_112_47#_c_348_n 0.00667101f $X=0.925 $Y=1.53 $X2=0 $Y2=0
cc_141 N_A_c_104_n N_A_112_47#_c_349_n 0.0138393f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_c_113_n N_A_112_47#_c_374_n 0.0179633f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_114_n N_A_112_47#_c_374_n 0.0121497f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_137_p N_A_112_47#_c_374_n 0.00533999f $X=0.84 $Y=1.175 $X2=0 $Y2=0
cc_145 N_A_c_119_n N_A_112_47#_c_374_n 0.00820484f $X=0.925 $Y=1.53 $X2=0 $Y2=0
cc_146 N_A_c_120_n N_A_112_47#_c_374_n 0.0329609f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_147 N_A_c_111_n N_A_112_47#_c_374_n 0.00303036f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_148 N_A_c_104_n N_A_112_47#_c_380_n 0.0110471f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_c_105_n N_A_112_47#_c_351_n 0.0127174f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_c_137_p N_A_112_47#_c_351_n 0.00105293f $X=0.84 $Y=1.175 $X2=0 $Y2=0
cc_151 N_A_c_120_n N_A_112_47#_c_351_n 0.00802966f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_152 N_A_c_105_n N_A_112_47#_c_384_n 5.82315e-19 $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_110_n N_A_112_47#_c_361_n 0.00468456f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_c_120_n N_A_112_47#_c_361_n 0.0137531f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_155 N_A_c_115_n N_A_112_47#_c_362_n 0.00435467f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_115_n N_A_112_47#_c_363_n 0.0136294f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_116_n N_A_112_47#_c_363_n 0.0117777f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_110_n N_A_112_47#_c_363_n 0.0730853f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_c_112_n N_A_112_47#_c_363_n 0.00929098f $X=3.355 $Y=1.202 $X2=0 $Y2=0
cc_160 N_A_c_110_n N_A_112_47#_c_364_n 0.0127997f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_c_120_n N_A_112_47#_c_364_n 0.0154683f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_162 N_A_c_104_n N_A_112_47#_c_355_n 0.00171616f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_c_137_p N_A_112_47#_c_355_n 0.0295837f $X=0.84 $Y=1.175 $X2=0 $Y2=0
cc_164 N_A_c_111_n N_A_112_47#_c_355_n 0.00486271f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_165 N_A_c_120_n N_A_112_47#_c_397_n 0.0130925f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_166 N_A_c_120_n N_A_27_297#_M1013_s 0.0018286f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_167 N_A_c_120_n N_A_27_297#_M1009_d 0.00158182f $X=1.86 $Y=1.53 $X2=0 $Y2=0
cc_168 N_A_c_113_n N_A_27_297#_c_515_n 0.00299383f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_114_n N_A_27_297#_c_515_n 0.00299383f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_113_n N_A_27_297#_c_511_n 6.73061e-19 $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_114_n N_A_27_297#_c_518_n 5.82762e-19 $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_c_119_n N_VPWR_M1001_d 0.00254399f $X=0.925 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_173 N_A_c_113_n N_VPWR_c_568_n 0.0032479f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_114_n N_VPWR_c_568_n 0.0032479f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_115_n N_VPWR_c_569_n 0.00300743f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_116_n N_VPWR_c_569_n 0.00300743f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_c_114_n N_VPWR_c_571_n 0.00702461f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_c_115_n N_VPWR_c_571_n 0.00702461f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_c_116_n N_VPWR_c_573_n 0.00702461f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_c_113_n N_VPWR_c_567_n 0.00655851f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_c_114_n N_VPWR_c_567_n 0.0056586f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_c_115_n N_VPWR_c_567_n 0.00821692f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_c_116_n N_VPWR_c_567_n 0.00695979f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_c_113_n N_VPWR_c_577_n 0.00702461f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_c_115_n N_A_510_297#_c_657_n 0.0112605f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_c_116_n N_A_510_297#_c_657_n 0.0112175f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_c_104_n N_VGND_c_757_n 0.00438629f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_104_n N_VGND_c_758_n 0.00423334f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_105_n N_VGND_c_758_n 0.00437852f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_105_n N_VGND_c_759_n 0.00276126f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_106_n N_VGND_c_761_n 0.00223901f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_c_109_n N_VGND_c_761_n 2.22494e-19 $X=2.08 $Y=1.175 $X2=0 $Y2=0
cc_193 N_A_c_110_n N_VGND_c_761_n 0.00470501f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_c_106_n N_VGND_c_762_n 0.00268723f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_107_n N_VGND_c_762_n 0.00268723f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_106_n N_VGND_c_765_n 0.00437852f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_107_n N_VGND_c_767_n 0.00421816f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_c_104_n N_VGND_c_772_n 0.00692693f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_c_105_n N_VGND_c_772_n 0.00627444f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_c_106_n N_VGND_c_772_n 0.00721278f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_107_n N_VGND_c_772_n 0.00591527f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_c_106_n N_A_510_47#_c_859_n 0.0106572f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_c_107_n N_A_510_47#_c_859_n 0.0114066f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_c_110_n N_A_510_47#_c_859_n 0.045703f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_c_112_n N_A_510_47#_c_859_n 0.0047738f $X=3.355 $Y=1.202 $X2=0 $Y2=0
cc_206 N_A_c_110_n N_A_510_47#_c_860_n 0.0252819f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_c_112_n N_A_510_47#_c_860_n 0.00137765f $X=3.355 $Y=1.202 $X2=0 $Y2=0
cc_208 N_A_c_106_n N_A_510_47#_c_868_n 4.68304e-19 $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_c_107_n N_A_510_47#_c_868_n 0.00390262f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_c_107_n N_A_510_47#_c_870_n 0.00374052f $X=3.355 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B_c_240_n N_A_112_47#_c_374_n 0.0107885f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_212 N_B_c_230_n N_A_112_47#_c_351_n 0.00879976f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B_c_231_n N_A_112_47#_c_351_n 3.48922e-19 $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B_c_234_n N_A_112_47#_c_351_n 0.00650896f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_215 N_B_c_235_n N_A_112_47#_c_351_n 0.00797709f $X=1.395 $Y=1.19 $X2=0 $Y2=0
cc_216 N_B_c_236_n N_A_112_47#_c_351_n 0.0369526f $X=1.475 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B_c_237_n N_A_112_47#_c_351_n 0.00579101f $X=1.92 $Y=1.202 $X2=0 $Y2=0
cc_218 N_B_c_230_n N_A_112_47#_c_384_n 0.00850899f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B_c_241_n N_A_112_47#_c_361_n 0.0124173f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_220 N_B_c_234_n N_A_112_47#_c_361_n 0.00186462f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_221 N_B_c_241_n N_A_112_47#_c_362_n 0.00547967f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_222 N_B_c_242_n N_A_112_47#_c_363_n 0.0120687f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B_c_243_n N_A_112_47#_c_363_n 0.0142166f $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_224 N_B_c_234_n N_A_112_47#_c_363_n 0.0144347f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_225 B N_A_112_47#_c_363_n 0.00704316f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_226 N_B_c_238_n N_A_112_47#_c_363_n 0.0515453f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_227 N_B_c_239_n N_A_112_47#_c_363_n 0.0092979f $X=4.375 $Y=1.202 $X2=0 $Y2=0
cc_228 N_B_c_241_n N_A_112_47#_c_364_n 0.00113114f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B_c_234_n N_A_112_47#_c_364_n 0.00139134f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_230 N_B_c_243_n N_A_112_47#_c_352_n 7.99457e-19 $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_231 N_B_c_238_n N_A_112_47#_c_352_n 0.00110099f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_232 N_B_c_239_n N_A_112_47#_c_352_n 0.00362886f $X=4.375 $Y=1.202 $X2=0 $Y2=0
cc_233 N_B_c_238_n N_A_112_47#_c_353_n 0.0072319f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_234 N_B_c_239_n N_A_112_47#_c_353_n 0.00107803f $X=4.375 $Y=1.202 $X2=0 $Y2=0
cc_235 N_B_c_240_n N_A_27_297#_c_519_n 0.00976749f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_236 N_B_c_241_n N_A_27_297#_c_519_n 0.0100164f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B_c_240_n N_A_27_297#_c_518_n 0.00375678f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_238 N_B_c_241_n N_A_27_297#_c_518_n 7.48748e-19 $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_239 N_B_c_242_n N_VPWR_c_570_n 0.00513149f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_240 N_B_c_243_n N_VPWR_c_570_n 0.00315692f $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_241 N_B_c_240_n N_VPWR_c_571_n 0.00429453f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_242 N_B_c_241_n N_VPWR_c_571_n 0.00429453f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_243 N_B_c_242_n N_VPWR_c_573_n 0.00702461f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B_c_243_n N_VPWR_c_575_n 0.00702461f $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_245 N_B_c_240_n N_VPWR_c_567_n 0.00596028f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_246 N_B_c_241_n N_VPWR_c_567_n 0.00734734f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_247 N_B_c_242_n N_VPWR_c_567_n 0.0071456f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B_c_243_n N_VPWR_c_567_n 0.00835069f $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_249 N_B_c_241_n N_A_510_297#_c_659_n 0.00372147f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_250 N_B_c_241_n N_A_510_297#_c_660_n 5.81899e-19 $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_251 N_B_c_242_n N_A_510_297#_c_661_n 0.0115086f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B_c_243_n N_A_510_297#_c_661_n 0.0115788f $X=4.375 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B_c_232_n N_X_c_704_n 0.00289058f $X=3.825 $Y=0.995 $X2=0 $Y2=0
cc_254 B N_X_c_704_n 0.00191347f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_255 N_B_c_238_n N_X_c_704_n 0.0368306f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B_c_239_n N_X_c_704_n 0.0061036f $X=4.375 $Y=1.202 $X2=0 $Y2=0
cc_257 N_B_c_233_n N_X_c_705_n 0.0115877f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B_c_230_n N_VGND_c_759_n 0.00359159f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_259 N_B_c_230_n N_VGND_c_760_n 0.00396605f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_260 N_B_c_231_n N_VGND_c_760_n 0.00585385f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_261 N_B_c_231_n N_VGND_c_761_n 0.00438629f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_262 N_B_c_234_n N_VGND_c_761_n 0.00123192f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_263 N_B_c_233_n N_VGND_c_763_n 0.0019578f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_264 N_B_c_232_n N_VGND_c_767_n 0.00357877f $X=3.825 $Y=0.995 $X2=0 $Y2=0
cc_265 N_B_c_233_n N_VGND_c_767_n 0.00357877f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_266 N_B_c_230_n N_VGND_c_772_n 0.00583329f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_267 N_B_c_231_n N_VGND_c_772_n 0.0119902f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_268 N_B_c_232_n N_VGND_c_772_n 0.00578582f $X=3.825 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B_c_233_n N_VGND_c_772_n 0.00692199f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B_c_231_n N_A_510_47#_c_858_n 0.0031408f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_271 N_B_c_232_n N_A_510_47#_c_859_n 9.49477e-19 $X=3.825 $Y=0.995 $X2=0 $Y2=0
cc_272 N_B_c_234_n N_A_510_47#_c_859_n 0.010004f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_273 N_B_c_231_n N_A_510_47#_c_860_n 0.00319308f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_274 N_B_c_234_n N_A_510_47#_c_860_n 0.00254218f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_275 N_B_c_232_n N_A_510_47#_c_861_n 0.013128f $X=3.825 $Y=0.995 $X2=0 $Y2=0
cc_276 N_B_c_233_n N_A_510_47#_c_861_n 0.0104406f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_277 B N_A_510_47#_c_861_n 0.00365912f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_278 N_B_c_238_n N_A_510_47#_c_861_n 0.00308757f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A_112_47#_c_348_n N_A_27_297#_M1001_s 0.00561099f $X=0.205 $Y=1.785
+ $X2=-0.19 $Y2=-0.24
cc_280 N_A_112_47#_c_374_n N_A_27_297#_M1001_s 0.00344657f $X=1.56 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_281 N_A_112_47#_c_360_n N_A_27_297#_M1001_s 0.00252471f $X=0.29 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_282 N_A_112_47#_c_374_n N_A_27_297#_M1013_s 0.00352135f $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_283 N_A_112_47#_c_361_n N_A_27_297#_M1009_d 0.00616915f $X=2.25 $Y=1.87 $X2=0
+ $Y2=0
cc_284 N_A_112_47#_c_362_n N_A_27_297#_M1009_d 0.00232242f $X=2.335 $Y=1.785
+ $X2=0 $Y2=0
cc_285 N_A_112_47#_c_364_n N_A_27_297#_M1009_d 0.00137528f $X=2.42 $Y=1.53 $X2=0
+ $Y2=0
cc_286 N_A_112_47#_M1006_s N_A_27_297#_c_519_n 0.00352392f $X=1.54 $Y=1.485
+ $X2=0 $Y2=0
cc_287 N_A_112_47#_c_374_n N_A_27_297#_c_519_n 0.00597191f $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_288 N_A_112_47#_c_361_n N_A_27_297#_c_519_n 0.00608347f $X=2.25 $Y=1.87 $X2=0
+ $Y2=0
cc_289 N_A_112_47#_c_397_n N_A_27_297#_c_519_n 0.0127274f $X=1.685 $Y=1.87 $X2=0
+ $Y2=0
cc_290 N_A_112_47#_c_361_n N_A_27_297#_c_534_n 0.0151964f $X=2.25 $Y=1.87 $X2=0
+ $Y2=0
cc_291 N_A_112_47#_c_374_n N_A_27_297#_c_515_n 0.0190031f $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_292 N_A_112_47#_c_374_n N_A_27_297#_c_511_n 0.00242129f $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_293 N_A_112_47#_c_360_n N_A_27_297#_c_511_n 0.00499157f $X=0.29 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_112_47#_c_374_n N_A_27_297#_c_512_n 0.004685f $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_295 N_A_112_47#_c_360_n N_A_27_297#_c_512_n 0.0120194f $X=0.29 $Y=1.87 $X2=0
+ $Y2=0
cc_296 N_A_112_47#_c_374_n N_A_27_297#_c_518_n 0.00822939f $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_297 N_A_112_47#_c_397_n N_A_27_297#_c_518_n 0.00140981f $X=1.685 $Y=1.87
+ $X2=0 $Y2=0
cc_298 N_A_112_47#_c_374_n N_A_27_297#_c_542_n 0.0121336f $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_299 N_A_112_47#_c_374_n N_VPWR_M1001_d 0.00394424f $X=1.56 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_300 N_A_112_47#_c_363_n N_VPWR_M1018_s 0.00187547f $X=5.015 $Y=1.53 $X2=0
+ $Y2=0
cc_301 N_A_112_47#_c_363_n N_VPWR_M1005_s 0.00246156f $X=5.015 $Y=1.53 $X2=0
+ $Y2=0
cc_302 N_A_112_47#_c_374_n N_VPWR_c_568_n 0.0124746f $X=1.56 $Y=1.87 $X2=0 $Y2=0
cc_303 N_A_112_47#_c_357_n N_VPWR_c_575_n 0.00429453f $X=5.365 $Y=1.41 $X2=0
+ $Y2=0
cc_304 N_A_112_47#_c_358_n N_VPWR_c_575_n 0.00429453f $X=5.835 $Y=1.41 $X2=0
+ $Y2=0
cc_305 N_A_112_47#_M1006_s N_VPWR_c_567_n 0.00231289f $X=1.54 $Y=1.485 $X2=0
+ $Y2=0
cc_306 N_A_112_47#_c_357_n N_VPWR_c_567_n 0.00734734f $X=5.365 $Y=1.41 $X2=0
+ $Y2=0
cc_307 N_A_112_47#_c_358_n N_VPWR_c_567_n 0.00706378f $X=5.835 $Y=1.41 $X2=0
+ $Y2=0
cc_308 N_A_112_47#_c_374_n N_VPWR_c_567_n 8.00021e-19 $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_309 N_A_112_47#_c_361_n N_VPWR_c_567_n 0.00673268f $X=2.25 $Y=1.87 $X2=0
+ $Y2=0
cc_310 N_A_112_47#_c_363_n N_A_510_297#_M1018_d 0.00321105f $X=5.015 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_311 N_A_112_47#_c_363_n N_A_510_297#_M1019_d 0.00187091f $X=5.015 $Y=1.53
+ $X2=0 $Y2=0
cc_312 N_A_112_47#_c_363_n N_A_510_297#_M1010_d 0.00291237f $X=5.015 $Y=1.53
+ $X2=0 $Y2=0
cc_313 N_A_112_47#_c_363_n N_A_510_297#_M1011_d 0.00463079f $X=5.015 $Y=1.53
+ $X2=0 $Y2=0
cc_314 N_A_112_47#_c_363_n N_A_510_297#_c_657_n 0.0359197f $X=5.015 $Y=1.53
+ $X2=0 $Y2=0
cc_315 N_A_112_47#_c_361_n N_A_510_297#_c_660_n 0.0155001f $X=2.25 $Y=1.87 $X2=0
+ $Y2=0
cc_316 N_A_112_47#_c_363_n N_A_510_297#_c_660_n 0.0135795f $X=5.015 $Y=1.53
+ $X2=0 $Y2=0
cc_317 N_A_112_47#_c_357_n N_A_510_297#_c_670_n 0.0143578f $X=5.365 $Y=1.41
+ $X2=0 $Y2=0
cc_318 N_A_112_47#_c_358_n N_A_510_297#_c_670_n 0.01161f $X=5.835 $Y=1.41 $X2=0
+ $Y2=0
cc_319 N_A_112_47#_c_363_n N_A_510_297#_c_655_n 0.0037422f $X=5.015 $Y=1.53
+ $X2=0 $Y2=0
cc_320 N_A_112_47#_c_363_n N_A_510_297#_c_673_n 0.013815f $X=5.015 $Y=1.53 $X2=0
+ $Y2=0
cc_321 N_A_112_47#_c_363_n N_A_510_297#_c_661_n 0.081218f $X=5.015 $Y=1.53 $X2=0
+ $Y2=0
cc_322 N_A_112_47#_c_363_n N_A_510_297#_c_656_n 0.0150001f $X=5.015 $Y=1.53
+ $X2=0 $Y2=0
cc_323 N_A_112_47#_c_354_n N_A_510_297#_c_656_n 0.00179065f $X=5.56 $Y=1.16
+ $X2=0 $Y2=0
cc_324 N_A_112_47#_c_358_n N_X_c_707_n 0.0183165f $X=5.835 $Y=1.41 $X2=0 $Y2=0
cc_325 N_A_112_47#_c_356_n N_X_c_707_n 0.00107224f $X=5.835 $Y=1.202 $X2=0 $Y2=0
cc_326 N_A_112_47#_c_347_n N_X_c_702_n 0.0140232f $X=5.86 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_112_47#_c_347_n N_X_c_703_n 0.0211434f $X=5.86 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A_112_47#_c_354_n N_X_c_703_n 0.0103529f $X=5.56 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_112_47#_c_346_n N_X_c_705_n 0.0109318f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_112_47#_c_363_n N_X_c_705_n 0.0178076f $X=5.015 $Y=1.53 $X2=0 $Y2=0
cc_331 N_A_112_47#_c_353_n N_X_c_705_n 0.0141442f $X=5.185 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A_112_47#_c_354_n N_X_c_705_n 0.0392005f $X=5.56 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A_112_47#_c_346_n N_X_c_706_n 0.00536716f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_112_47#_c_356_n N_X_c_706_n 0.0047334f $X=5.835 $Y=1.202 $X2=0 $Y2=0
cc_335 N_A_112_47#_c_357_n N_X_c_709_n 8.03792e-19 $X=5.365 $Y=1.41 $X2=0 $Y2=0
cc_336 N_A_112_47#_c_363_n N_X_c_709_n 0.00647942f $X=5.015 $Y=1.53 $X2=0 $Y2=0
cc_337 N_A_112_47#_c_352_n N_X_c_709_n 0.00171573f $X=5.1 $Y=1.445 $X2=0 $Y2=0
cc_338 N_A_112_47#_c_354_n N_X_c_709_n 0.0202439f $X=5.56 $Y=1.16 $X2=0 $Y2=0
cc_339 N_A_112_47#_c_356_n N_X_c_709_n 0.00667431f $X=5.835 $Y=1.202 $X2=0 $Y2=0
cc_340 N_A_112_47#_c_349_n N_VGND_M1002_d 6.44201e-19 $X=0.53 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_341 N_A_112_47#_c_350_n N_VGND_M1002_d 0.00301785f $X=0.29 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_342 N_A_112_47#_c_351_n N_VGND_M1015_d 0.00251047f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_343 N_A_112_47#_c_350_n N_VGND_c_756_n 0.00114168f $X=0.29 $Y=0.815 $X2=0
+ $Y2=0
cc_344 N_A_112_47#_c_349_n N_VGND_c_757_n 0.00491543f $X=0.53 $Y=0.815 $X2=0
+ $Y2=0
cc_345 N_A_112_47#_c_350_n N_VGND_c_757_n 0.00856149f $X=0.29 $Y=0.815 $X2=0
+ $Y2=0
cc_346 N_A_112_47#_c_349_n N_VGND_c_758_n 0.00198695f $X=0.53 $Y=0.815 $X2=0
+ $Y2=0
cc_347 N_A_112_47#_c_380_n N_VGND_c_758_n 0.0231806f $X=0.745 $Y=0.39 $X2=0
+ $Y2=0
cc_348 N_A_112_47#_c_351_n N_VGND_c_758_n 0.00254521f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_349 N_A_112_47#_c_351_n N_VGND_c_759_n 0.0122589f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_350 N_A_112_47#_c_384_n N_VGND_c_759_n 0.0223967f $X=1.685 $Y=0.39 $X2=0
+ $Y2=0
cc_351 N_A_112_47#_c_351_n N_VGND_c_760_n 0.00199443f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_352 N_A_112_47#_c_384_n N_VGND_c_760_n 0.023074f $X=1.685 $Y=0.39 $X2=0 $Y2=0
cc_353 N_A_112_47#_c_346_n N_VGND_c_763_n 0.00438629f $X=5.34 $Y=0.995 $X2=0
+ $Y2=0
cc_354 N_A_112_47#_c_347_n N_VGND_c_764_n 0.00438629f $X=5.86 $Y=0.995 $X2=0
+ $Y2=0
cc_355 N_A_112_47#_c_346_n N_VGND_c_770_n 0.00435595f $X=5.34 $Y=0.995 $X2=0
+ $Y2=0
cc_356 N_A_112_47#_c_347_n N_VGND_c_770_n 0.00437852f $X=5.86 $Y=0.995 $X2=0
+ $Y2=0
cc_357 N_A_112_47#_M1002_s N_VGND_c_772_n 0.00304143f $X=0.56 $Y=0.235 $X2=0
+ $Y2=0
cc_358 N_A_112_47#_M1016_s N_VGND_c_772_n 0.00324782f $X=1.55 $Y=0.235 $X2=0
+ $Y2=0
cc_359 N_A_112_47#_c_346_n N_VGND_c_772_n 0.00746942f $X=5.34 $Y=0.995 $X2=0
+ $Y2=0
cc_360 N_A_112_47#_c_347_n N_VGND_c_772_n 0.00722704f $X=5.86 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A_112_47#_c_349_n N_VGND_c_772_n 0.00412013f $X=0.53 $Y=0.815 $X2=0
+ $Y2=0
cc_362 N_A_112_47#_c_350_n N_VGND_c_772_n 0.0024413f $X=0.29 $Y=0.815 $X2=0
+ $Y2=0
cc_363 N_A_112_47#_c_380_n N_VGND_c_772_n 0.0143352f $X=0.745 $Y=0.39 $X2=0
+ $Y2=0
cc_364 N_A_112_47#_c_351_n N_VGND_c_772_n 0.00977515f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_365 N_A_112_47#_c_384_n N_VGND_c_772_n 0.0141066f $X=1.685 $Y=0.39 $X2=0
+ $Y2=0
cc_366 N_A_112_47#_c_363_n N_A_510_47#_c_859_n 0.0027094f $X=5.015 $Y=1.53 $X2=0
+ $Y2=0
cc_367 N_A_112_47#_c_351_n N_A_510_47#_c_860_n 0.00357823f $X=1.47 $Y=0.815
+ $X2=0 $Y2=0
cc_368 N_A_27_297#_c_515_n N_VPWR_M1001_d 4.93802e-19 $X=1.105 $Y=2.21 $X2=-0.19
+ $Y2=1.305
cc_369 N_A_27_297#_c_515_n N_VPWR_c_568_n 0.013934f $X=1.105 $Y=2.21 $X2=0 $Y2=0
cc_370 N_A_27_297#_c_511_n N_VPWR_c_568_n 3.55827e-19 $X=0.375 $Y=2.21 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_512_n N_VPWR_c_568_n 0.00390479f $X=0.23 $Y=2.21 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_518_n N_VPWR_c_568_n 3.64325e-19 $X=1.25 $Y=2.21 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_542_n N_VPWR_c_568_n 0.00389788f $X=1.25 $Y=2.21 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_c_519_n N_VPWR_c_571_n 0.0386815f $X=2.03 $Y=2.38 $X2=0 $Y2=0
cc_375 N_A_27_297#_c_534_n N_VPWR_c_571_n 0.0154343f $X=2.155 $Y=2.3 $X2=0 $Y2=0
cc_376 N_A_27_297#_c_515_n N_VPWR_c_571_n 0.00106736f $X=1.105 $Y=2.21 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_c_542_n N_VPWR_c_571_n 0.0143977f $X=1.25 $Y=2.21 $X2=0 $Y2=0
cc_378 N_A_27_297#_M1001_s N_VPWR_c_567_n 0.00126254f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_379 N_A_27_297#_M1013_s N_VPWR_c_567_n 0.00125832f $X=1.07 $Y=1.485 $X2=0
+ $Y2=0
cc_380 N_A_27_297#_M1009_d N_VPWR_c_567_n 0.00215913f $X=2.01 $Y=1.485 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_c_519_n N_VPWR_c_567_n 0.0225093f $X=2.03 $Y=2.38 $X2=0 $Y2=0
cc_382 N_A_27_297#_c_534_n N_VPWR_c_567_n 0.00938089f $X=2.155 $Y=2.3 $X2=0
+ $Y2=0
cc_383 N_A_27_297#_c_515_n N_VPWR_c_567_n 0.0607581f $X=1.105 $Y=2.21 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_c_511_n N_VPWR_c_567_n 0.0285979f $X=0.375 $Y=2.21 $X2=0
+ $Y2=0
cc_385 N_A_27_297#_c_512_n N_VPWR_c_567_n 0.00254937f $X=0.23 $Y=2.21 $X2=0
+ $Y2=0
cc_386 N_A_27_297#_c_518_n N_VPWR_c_567_n 0.0281768f $X=1.25 $Y=2.21 $X2=0 $Y2=0
cc_387 N_A_27_297#_c_542_n N_VPWR_c_567_n 0.00227213f $X=1.25 $Y=2.21 $X2=0
+ $Y2=0
cc_388 N_A_27_297#_c_515_n N_VPWR_c_577_n 0.00107419f $X=1.105 $Y=2.21 $X2=0
+ $Y2=0
cc_389 N_A_27_297#_c_511_n N_VPWR_c_577_n 3.6232e-19 $X=0.375 $Y=2.21 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_c_512_n N_VPWR_c_577_n 0.0175488f $X=0.23 $Y=2.21 $X2=0 $Y2=0
cc_391 N_A_27_297#_c_534_n N_A_510_297#_c_655_n 0.0230175f $X=2.155 $Y=2.3 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_567_n N_A_510_297#_M1018_d 0.00227295f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_393 N_VPWR_c_567_n N_A_510_297#_M1019_d 0.00250817f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_567_n N_A_510_297#_M1010_d 0.00228122f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_567_n N_A_510_297#_M1011_d 0.00217543f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_567_n N_A_510_297#_M1014_d 0.00303346f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_397 N_VPWR_M1018_s N_A_510_297#_c_657_n 0.00348982f $X=3 $Y=1.485 $X2=0 $Y2=0
cc_398 N_VPWR_c_569_n N_A_510_297#_c_657_n 0.0132478f $X=3.145 $Y=2.3 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_567_n N_A_510_297#_c_657_n 0.0141814f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_573_n N_A_510_297#_c_686_n 0.0149311f $X=3.96 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_567_n N_A_510_297#_c_686_n 0.00955092f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_575_n N_A_510_297#_c_670_n 0.0162749f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_567_n N_A_510_297#_c_670_n 0.00962421f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_571_n N_A_510_297#_c_655_n 0.0204786f $X=3.02 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_567_n N_A_510_297#_c_655_n 0.0119856f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_M1005_s N_A_510_297#_c_661_n 0.00460956f $X=3.94 $Y=1.485 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_570_n N_A_510_297#_c_661_n 0.0173877f $X=4.14 $Y=2.3 $X2=0 $Y2=0
cc_408 N_VPWR_c_567_n N_A_510_297#_c_661_n 0.014419f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_c_575_n N_A_510_297#_c_656_n 0.0902831f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_567_n N_A_510_297#_c_656_n 0.0535524f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_567_n N_X_M1011_s 0.00232895f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_412 N_A_510_297#_c_670_n N_X_M1011_s 0.00352392f $X=5.945 $Y=2.38 $X2=0 $Y2=0
cc_413 N_A_510_297#_c_670_n N_X_c_707_n 0.003919f $X=5.945 $Y=2.38 $X2=0 $Y2=0
cc_414 N_A_510_297#_M1014_d N_X_c_703_n 0.00411256f $X=5.925 $Y=1.485 $X2=0
+ $Y2=0
cc_415 N_A_510_297#_c_700_p N_X_c_703_n 0.0188231f $X=6.07 $Y=1.96 $X2=0 $Y2=0
cc_416 N_A_510_297#_c_670_n N_X_c_709_n 0.0134553f $X=5.945 $Y=2.38 $X2=0 $Y2=0
cc_417 N_X_c_705_n N_VGND_M1008_d 0.00315681f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_418 N_X_c_702_n N_VGND_M1012_d 0.00326372f $X=5.985 $Y=0.815 $X2=0 $Y2=0
cc_419 N_X_c_705_n N_VGND_c_763_n 0.0127273f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_420 N_X_c_702_n N_VGND_c_764_n 0.0140097f $X=5.985 $Y=0.815 $X2=0 $Y2=0
cc_421 N_X_c_705_n N_VGND_c_767_n 0.00401766f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_422 N_X_c_702_n N_VGND_c_769_n 0.00327334f $X=5.985 $Y=0.815 $X2=0 $Y2=0
cc_423 N_X_c_702_n N_VGND_c_770_n 0.00254521f $X=5.985 $Y=0.815 $X2=0 $Y2=0
cc_424 N_X_c_705_n N_VGND_c_770_n 0.00198695f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_425 N_X_c_706_n N_VGND_c_770_n 0.00589303f $X=5.765 $Y=0.775 $X2=0 $Y2=0
cc_426 N_X_M1000_d N_VGND_c_772_n 0.00342404f $X=3.9 $Y=0.235 $X2=0 $Y2=0
cc_427 N_X_M1008_s N_VGND_c_772_n 0.00439795f $X=5.415 $Y=0.235 $X2=0 $Y2=0
cc_428 N_X_c_702_n N_VGND_c_772_n 0.0112583f $X=5.985 $Y=0.815 $X2=0 $Y2=0
cc_429 N_X_c_705_n N_VGND_c_772_n 0.0126305f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_430 N_X_c_706_n N_VGND_c_772_n 0.0107037f $X=5.765 $Y=0.775 $X2=0 $Y2=0
cc_431 N_X_c_705_n N_A_510_47#_M1004_s 0.00319929f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_432 N_X_c_704_n N_A_510_47#_c_859_n 0.00627715f $X=4.305 $Y=0.775 $X2=0 $Y2=0
cc_433 N_X_M1000_d N_A_510_47#_c_861_n 0.00693401f $X=3.9 $Y=0.235 $X2=0 $Y2=0
cc_434 N_X_c_704_n N_A_510_47#_c_861_n 0.0211337f $X=4.305 $Y=0.775 $X2=0 $Y2=0
cc_435 N_X_c_705_n N_A_510_47#_c_861_n 0.0198081f $X=5.385 $Y=0.775 $X2=0 $Y2=0
cc_436 N_VGND_c_772_n N_A_510_47#_M1003_s 0.00258952f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_437 N_VGND_c_772_n N_A_510_47#_M1007_s 0.00256961f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_438 N_VGND_c_772_n N_A_510_47#_M1004_s 0.00209344f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_c_761_n N_A_510_47#_c_858_n 0.0168055f $X=2.155 $Y=0.39 $X2=0
+ $Y2=0
cc_440 N_VGND_c_765_n N_A_510_47#_c_858_n 0.0217962f $X=3.06 $Y=0 $X2=0 $Y2=0
cc_441 N_VGND_c_772_n N_A_510_47#_c_858_n 0.0126169f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_442 N_VGND_M1003_d N_A_510_47#_c_859_n 0.00162089f $X=3.01 $Y=0.235 $X2=0
+ $Y2=0
cc_443 N_VGND_c_762_n N_A_510_47#_c_859_n 0.0118745f $X=3.145 $Y=0.39 $X2=0
+ $Y2=0
cc_444 N_VGND_c_765_n N_A_510_47#_c_859_n 0.00254521f $X=3.06 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_c_767_n N_A_510_47#_c_859_n 0.00198695f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_772_n N_A_510_47#_c_859_n 0.0094839f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_447 N_VGND_c_767_n N_A_510_47#_c_870_n 0.0187477f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_448 N_VGND_c_772_n N_A_510_47#_c_870_n 0.0114026f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_449 N_VGND_c_763_n N_A_510_47#_c_861_n 0.0131818f $X=5.13 $Y=0.39 $X2=0 $Y2=0
cc_450 N_VGND_c_767_n N_A_510_47#_c_861_n 0.0626452f $X=5.045 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_772_n N_A_510_47#_c_861_n 0.0390083f $X=6.21 $Y=0 $X2=0 $Y2=0
