* File: sky130_fd_sc_hdll__o21ai_1.spice
* Created: Thu Aug 27 19:19:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21ai_1.pex.spice"
.subckt sky130_fd_sc_hdll__o21ai_1  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A1_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.2015 PD=1.04 PS=1.92 NRD=10.152 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1004 N_A_27_47#_M1004_d N_A2_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12675 PD=0.92 PS=1.04 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75000.8 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_27_47#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.38025 AS=0.08775 PD=2.47 PS=0.92 NRD=35.076 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1002 A_117_297# N_A1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.27 PD=1.23 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_A2_M1001_g A_117_297# VPB PHIGHVT L=0.18 W=1 AD=0.218824
+ AS=0.115 PD=1.67059 PS=1.23 NRD=18.715 NRS=11.8003 M=1 R=5.55556 SA=90000.6
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_Y_M1001_d VPB PHIGHVT L=0.18 W=0.7
+ AD=0.3815 AS=0.153176 PD=2.49 PS=1.16941 NRD=42.1974 NRS=12.6474 M=1 R=3.88889
+ SA=90001.2 SB=90000.5 A=0.126 P=1.76 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hdll__o21ai_1.pxi.spice"
*
.ends
*
*
