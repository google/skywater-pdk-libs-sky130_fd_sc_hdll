* File: sky130_fd_sc_hdll__or2_2.spice
* Created: Thu Aug 27 19:23:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or2_2.pex.spice"
.subckt sky130_fd_sc_hdll__or2_2  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1006 N_A_39_297#_M1006_d N_B_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1302 PD=0.69 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_39_297#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0920467 AS=0.0567 PD=0.828224 PS=0.69 NRD=35.712 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1003_d N_A_39_297#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.142453 AS=0.12025 PD=1.28178 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_39_297#_M1005_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 A_129_297# N_B_M1002_g N_A_39_297#_M1002_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0483 AS=0.1134 PD=0.65 PS=1.38 NRD=28.1316 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_129_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0963338 AS=0.0483 PD=0.81338 PS=0.65 NRD=81.7747 NRS=28.1316 M=1
+ R=2.33333 SA=90000.6 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1001 N_X_M1001_d N_A_39_297#_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.229366 PD=1.29 PS=1.93662 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1007 N_X_M1001_d N_A_39_297#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
c_179 A_129_297# 0 1.05688e-19 $X=0.645 $Y=1.485
*
.include "sky130_fd_sc_hdll__or2_2.pxi.spice"
*
.ends
*
*
