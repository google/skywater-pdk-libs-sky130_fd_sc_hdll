* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__muxb16to1_2 D[15] D[14] D[13] D[12] D[11] D[10] D[9] D[8]
+ D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] S[15] S[14] S[13] S[12] S[11] S[10] S[9]
+ S[8] S[7] S[6] S[5] S[4] S[3] S[2] S[1] S[0] VGND VNB VPB VPWR Z
X0 a_27_591# D[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_3421_915# D[13] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_2603_47# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_3891_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_4709_915# S[15] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X6 a_2112_333# a_1989_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X7 VGND S[13] a_3277_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X8 a_1566_793# S[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_3891_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X10 VPWR D[5] a_3400_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 Z a_4142_793# a_3891_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X12 a_27_911# D[8] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND D[15] a_4709_915# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Z a_278_265# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X15 VGND S[11] a_1989_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X16 Z S[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X17 a_4688_591# D[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND D[13] a_3421_915# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Z S[15] a_4709_915# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X20 a_845_69# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X21 a_4142_793# S[14] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X22 VPWR D[3] a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_1315_911# D[10] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR S[9] a_701_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 Z a_701_937# a_824_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X26 a_3400_591# D[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_3891_591# D[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 VPWR D[12] a_2603_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_1315_911# S[10] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X30 a_27_911# S[8] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X31 a_27_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 VGND D[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 Z a_4142_265# a_3891_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X34 a_824_591# a_701_937# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X35 VGND D[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VGND D[5] a_3421_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VGND S[15] a_4565_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X38 a_27_591# a_278_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X39 a_2112_591# D[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 a_278_793# S[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 a_2603_591# D[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X42 VPWR D[9] a_824_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X43 VPWR D[10] a_1315_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 VGND S[5] a_3277_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X45 a_1566_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 VGND S[7] a_4565_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X47 Z S[10] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X48 VPWR S[15] a_4565_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X49 a_4688_333# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X50 Z a_4565_937# a_4688_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X51 VGND D[6] a_3891_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X52 Z a_701_47# a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X53 a_824_591# D[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X54 a_1315_591# D[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X55 a_2603_911# D[12] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 a_845_69# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X57 a_2133_69# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X58 a_3421_69# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X59 a_3891_911# S[14] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 a_824_333# a_701_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X61 VPWR S[1] a_701_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 a_2603_911# S[12] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X63 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X64 a_3891_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X65 a_3400_333# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X66 a_3891_591# a_4142_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X67 Z a_3277_937# a_3400_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X68 VPWR S[13] a_3277_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X69 a_2854_265# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X70 Z S[4] a_2603_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X71 a_27_297# a_278_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X72 a_4142_793# S[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X73 a_4142_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X74 VPWR D[4] a_2603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X75 VGND D[14] a_3891_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X76 a_27_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X77 VGND S[1] a_701_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X78 VGND D[12] a_2603_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X79 Z S[9] a_845_915# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X80 Z a_4565_47# a_4688_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X81 VPWR D[8] a_27_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X82 Z S[14] a_3891_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X83 a_2112_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X84 a_278_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X85 VGND D[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X86 a_2603_297# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X87 a_2854_793# S[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X88 VPWR D[1] a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X89 Z S[12] a_2603_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X90 VPWR D[2] a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X91 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X92 a_2603_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X93 a_3891_911# D[14] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X94 Z S[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X95 VPWR S[7] a_4565_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X96 a_27_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X97 Z S[5] a_3421_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X98 VPWR D[15] a_4688_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X99 a_845_915# D[9] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X100 Z S[7] a_4709_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X101 a_3891_297# a_4142_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X102 Z a_3277_47# a_3400_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X103 a_2133_915# S[11] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X104 a_824_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X105 a_1315_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X106 Z a_2854_793# a_2603_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X107 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X108 a_4709_69# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X109 a_4709_915# D[15] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X110 VGND S[9] a_701_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X111 VPWR S[5] a_3277_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X112 VPWR S[11] a_1989_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X113 a_4142_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X114 VPWR D[14] a_3891_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X115 a_2603_591# a_2854_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X116 a_4688_591# a_4565_937# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X117 VGND D[9] a_845_915# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X118 a_2133_69# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X119 Z a_1566_793# a_1315_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X120 a_3421_69# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X121 Z S[11] a_2133_915# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X122 a_4709_69# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X123 VGND D[7] a_4709_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X124 Z S[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X125 VPWR D[0] a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X126 a_2854_265# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X127 a_1315_591# a_1566_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X128 a_3400_591# a_3277_937# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X129 Z a_2854_265# a_2603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X130 a_2133_915# D[11] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X131 a_3421_915# S[13] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X132 Z a_1989_937# a_2112_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X133 VGND S[3] a_1989_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X134 VPWR D[7] a_4688_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X135 VGND D[10] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X136 VPWR D[13] a_3400_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X137 VGND D[8] a_27_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X138 a_845_915# S[9] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X139 a_278_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X140 a_2603_297# a_2854_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X141 a_4688_333# a_4565_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X142 a_2112_591# a_1989_937# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X143 VGND D[4] a_2603_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X144 Z a_1566_265# a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X145 Z S[8] a_27_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X146 VGND D[11] a_2133_915# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X147 VPWR D[6] a_3891_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X148 Z a_278_793# a_27_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X149 Z S[13] a_3421_915# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X150 VPWR D[11] a_2112_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X151 VPWR S[3] a_1989_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X152 Z S[6] a_3891_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X153 a_1315_297# a_1566_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X154 a_1566_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X155 a_3400_333# a_3277_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X156 a_2854_793# S[12] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X157 Z a_1989_47# a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X158 a_1566_793# S[10] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X159 a_278_793# S[8] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
.ends
