* File: sky130_fd_sc_hdll__or2_8.pex.spice
* Created: Thu Aug 27 19:23:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR2_8%A 1 3 4 6 7 9 10 12 13 19 20 25
c39 10 0 1.11304e-19 $X=0.985 $Y=1.41
r40 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r41 19 25 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=0.92 $Y=1.175
+ $X2=0.695 $Y2=1.175
r42 18 20 5.07368 $w=3.8e-07 $l=4e-08 $layer=POLY_cond $X=0.92 $Y=1.202 $X2=0.96
+ $Y2=1.202
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.92
+ $Y=1.16 $X2=0.92 $Y2=1.16
r44 16 18 48.2 $w=3.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.54 $Y=1.202 $X2=0.92
+ $Y2=1.202
r45 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r46 13 25 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.175
+ $X2=0.695 $Y2=1.175
r47 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r48 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r49 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r50 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=0.56
r51 4 16 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r52 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r53 1 15 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r54 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_8%B 1 3 4 6 7 9 10 12 13 19 20 25
r55 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.9 $Y=1.202
+ $X2=1.925 $Y2=1.202
r56 19 25 13.5864 $w=1.98e-07 $l=2.45e-07 $layer=LI1_cond $X=1.86 $Y=1.175
+ $X2=1.615 $Y2=1.175
r57 18 20 5.07368 $w=3.8e-07 $l=4e-08 $layer=POLY_cond $X=1.86 $Y=1.202 $X2=1.9
+ $Y2=1.202
r58 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.86
+ $Y=1.16 $X2=1.86 $Y2=1.16
r59 16 18 48.2 $w=3.8e-07 $l=3.8e-07 $layer=POLY_cond $X=1.48 $Y=1.202 $X2=1.86
+ $Y2=1.202
r60 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.48 $Y2=1.202
r61 13 25 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=1.175
+ $X2=1.615 $Y2=1.175
r62 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r63 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r64 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.9 $Y=0.995 $X2=1.9
+ $Y2=1.202
r65 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.9 $Y=0.995 $X2=1.9
+ $Y2=0.56
r66 4 16 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=1.202
r67 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.48 $Y=0.995 $X2=1.48
+ $Y2=0.56
r68 1 15 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r69 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_8%A_123_47# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 60 62 63
+ 66 70 72 75 77 83 86 88 89 106
c218 88 0 1.11304e-19 $X=1.69 $Y=1.62
r219 106 107 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.18 $Y=1.202
+ $X2=6.205 $Y2=1.202
r220 105 106 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=5.76 $Y=1.202
+ $X2=6.18 $Y2=1.202
r221 104 105 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.735 $Y=1.202
+ $X2=5.76 $Y2=1.202
r222 101 102 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.24 $Y=1.202
+ $X2=5.265 $Y2=1.202
r223 100 101 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=4.82 $Y=1.202
+ $X2=5.24 $Y2=1.202
r224 99 100 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.795 $Y=1.202
+ $X2=4.82 $Y2=1.202
r225 98 99 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=4.325 $Y=1.202
+ $X2=4.795 $Y2=1.202
r226 97 98 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.3 $Y=1.202
+ $X2=4.325 $Y2=1.202
r227 96 97 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=3.88 $Y=1.202
+ $X2=4.3 $Y2=1.202
r228 95 96 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.855 $Y=1.202
+ $X2=3.88 $Y2=1.202
r229 94 95 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=3.385 $Y=1.202
+ $X2=3.855 $Y2=1.202
r230 93 94 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.36 $Y=1.202
+ $X2=3.385 $Y2=1.202
r231 90 91 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.915 $Y=1.202
+ $X2=2.94 $Y2=1.202
r232 84 104 49.1168 $w=3.68e-07 $l=3.75e-07 $layer=POLY_cond $X=5.36 $Y=1.202
+ $X2=5.735 $Y2=1.202
r233 84 102 12.4429 $w=3.68e-07 $l=9.5e-08 $layer=POLY_cond $X=5.36 $Y=1.202
+ $X2=5.265 $Y2=1.202
r234 83 84 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=5.36
+ $Y=1.16 $X2=5.36 $Y2=1.16
r235 81 93 49.7717 $w=3.68e-07 $l=3.8e-07 $layer=POLY_cond $X=2.98 $Y=1.202
+ $X2=3.36 $Y2=1.202
r236 81 91 5.23913 $w=3.68e-07 $l=4e-08 $layer=POLY_cond $X=2.98 $Y=1.202
+ $X2=2.94 $Y2=1.202
r237 80 83 131.982 $w=1.98e-07 $l=2.38e-06 $layer=LI1_cond $X=2.98 $Y=1.175
+ $X2=5.36 $Y2=1.175
r238 80 81 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=2.98
+ $Y=1.16 $X2=2.98 $Y2=1.16
r239 78 89 0.966048 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=2.375 $Y=1.175
+ $X2=2.285 $Y2=1.175
r240 78 80 33.55 $w=1.98e-07 $l=6.05e-07 $layer=LI1_cond $X=2.375 $Y=1.175
+ $X2=2.98 $Y2=1.175
r241 76 89 5.63431 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=2.285 $Y=1.275
+ $X2=2.285 $Y2=1.175
r242 76 77 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=2.285 $Y=1.275
+ $X2=2.285 $Y2=1.445
r243 75 89 5.63431 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=2.285 $Y=1.075
+ $X2=2.285 $Y2=1.175
r244 74 75 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=2.285 $Y=0.905
+ $X2=2.285 $Y2=1.075
r245 73 88 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=1.555
+ $X2=1.69 $Y2=1.555
r246 72 77 6.90553 $w=2.2e-07 $l=1.48324e-07 $layer=LI1_cond $X=2.195 $Y=1.555
+ $X2=2.285 $Y2=1.445
r247 72 73 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.195 $Y=1.555
+ $X2=1.855 $Y2=1.555
r248 71 86 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.855 $Y=0.82
+ $X2=1.69 $Y2=0.815
r249 70 74 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.195 $Y=0.82
+ $X2=2.285 $Y2=0.905
r250 70 71 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.195 $Y=0.82
+ $X2=1.855 $Y2=0.82
r251 64 86 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=0.725
+ $X2=1.69 $Y2=0.815
r252 64 66 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.69 $Y=0.725
+ $X2=1.69 $Y2=0.39
r253 62 86 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=0.815
+ $X2=1.69 $Y2=0.815
r254 62 63 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=1.525 $Y=0.815
+ $X2=0.915 $Y2=0.815
r255 58 63 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.75 $Y=0.725
+ $X2=0.915 $Y2=0.815
r256 58 60 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.75 $Y=0.725
+ $X2=0.75 $Y2=0.39
r257 55 107 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.205 $Y=1.41
+ $X2=6.205 $Y2=1.202
r258 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.205 $Y=1.41
+ $X2=6.205 $Y2=1.985
r259 52 106 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.18 $Y=0.995
+ $X2=6.18 $Y2=1.202
r260 52 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.18 $Y=0.995
+ $X2=6.18 $Y2=0.56
r261 49 105 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.76 $Y=0.995
+ $X2=5.76 $Y2=1.202
r262 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.76 $Y=0.995
+ $X2=5.76 $Y2=0.56
r263 46 104 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.735 $Y=1.41
+ $X2=5.735 $Y2=1.202
r264 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.735 $Y=1.41
+ $X2=5.735 $Y2=1.985
r265 43 102 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.202
r266 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.985
r267 40 101 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=1.202
r268 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=0.56
r269 37 100 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=1.202
r270 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=0.56
r271 34 99 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.202
r272 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.985
r273 31 98 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.325 $Y=1.41
+ $X2=4.325 $Y2=1.202
r274 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.325 $Y=1.41
+ $X2=4.325 $Y2=1.985
r275 28 97 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.3 $Y=0.995
+ $X2=4.3 $Y2=1.202
r276 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.3 $Y=0.995
+ $X2=4.3 $Y2=0.56
r277 25 96 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.88 $Y=0.995
+ $X2=3.88 $Y2=1.202
r278 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.88 $Y=0.995
+ $X2=3.88 $Y2=0.56
r279 22 95 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.855 $Y=1.41
+ $X2=3.855 $Y2=1.202
r280 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.855 $Y=1.41
+ $X2=3.855 $Y2=1.985
r281 19 94 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.385 $Y2=1.202
r282 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.385 $Y2=1.985
r283 16 93 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=1.202
r284 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=0.56
r285 13 91 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.94 $Y=0.995
+ $X2=2.94 $Y2=1.202
r286 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.94 $Y=0.995
+ $X2=2.94 $Y2=0.56
r287 10 90 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.915 $Y=1.41
+ $X2=2.915 $Y2=1.202
r288 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.915 $Y=1.41
+ $X2=2.915 $Y2=1.985
r289 3 88 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.62
r290 2 66 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.39
r291 1 60 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_8%A_27_297# 1 2 3 10 12 14 16 17 18 22
r34 20 22 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=2.175 $Y=2.295
+ $X2=2.175 $Y2=2
r35 19 29 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.355 $Y=2.38
+ $X2=1.22 $Y2=2.38
r36 18 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.025 $Y=2.38
+ $X2=2.175 $Y2=2.295
r37 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=2.38
+ $X2=1.355 $Y2=2.38
r38 17 29 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.295
+ $X2=1.22 $Y2=2.38
r39 16 27 3.04322 $w=2.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.56
r40 16 17 26.8903 $w=2.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=2.295
r41 15 25 4.39997 $w=2.1e-07 $l=1.63e-07 $layer=LI1_cond $X=0.415 $Y=1.56
+ $X2=0.252 $Y2=1.56
r42 14 27 3.91272 $w=2.1e-07 $l=1.35e-07 $layer=LI1_cond $X=1.085 $Y=1.56
+ $X2=1.22 $Y2=1.56
r43 14 15 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.085 $Y=1.56
+ $X2=0.415 $Y2=1.56
r44 10 25 2.83434 $w=3.25e-07 $l=1.05e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=1.56
r45 10 12 22.517 $w=3.23e-07 $l=6.35e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=2.3
r46 3 22 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2
r47 2 29 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r48 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r49 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r50 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_8%VPWR 1 2 3 4 5 6 21 25 31 35 39 43 46 47 49
+ 50 52 53 55 56 58 59 60 62 87 88 91
r91 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r92 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r93 85 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r94 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r95 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r96 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r97 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r98 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r99 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r100 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r101 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r102 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r103 70 73 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r104 70 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r105 69 72 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r106 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r107 67 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=0.75 $Y2=2.72
r108 67 69 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r109 62 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=2.72
+ $X2=0.75 $Y2=2.72
r110 62 64 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.585 $Y=2.72
+ $X2=0.23 $Y2=2.72
r111 60 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r112 60 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r113 58 84 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.305 $Y=2.72
+ $X2=6.21 $Y2=2.72
r114 58 59 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.305 $Y=2.72
+ $X2=6.44 $Y2=2.72
r115 57 87 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=6.67 $Y2=2.72
r116 57 59 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=6.44 $Y2=2.72
r117 55 81 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.365 $Y=2.72
+ $X2=5.29 $Y2=2.72
r118 55 56 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.365 $Y=2.72
+ $X2=5.5 $Y2=2.72
r119 54 84 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=6.21 $Y2=2.72
r120 54 56 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=5.5 $Y2=2.72
r121 52 78 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.37 $Y2=2.72
r122 52 53 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.56 $Y2=2.72
r123 51 81 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.695 $Y=2.72
+ $X2=5.29 $Y2=2.72
r124 51 53 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.695 $Y=2.72
+ $X2=4.56 $Y2=2.72
r125 49 75 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.45 $Y2=2.72
r126 49 50 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.485 $Y=2.72
+ $X2=3.62 $Y2=2.72
r127 48 78 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=4.37 $Y2=2.72
r128 48 50 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.62 $Y2=2.72
r129 46 72 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.53 $Y2=2.72
r130 46 47 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.68 $Y2=2.72
r131 45 75 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=3.45 $Y2=2.72
r132 45 47 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=2.68 $Y2=2.72
r133 41 59 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=2.635
+ $X2=6.44 $Y2=2.72
r134 41 43 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.44 $Y=2.635
+ $X2=6.44 $Y2=2
r135 37 56 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=2.635
+ $X2=5.5 $Y2=2.72
r136 37 39 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.5 $Y=2.635
+ $X2=5.5 $Y2=2
r137 33 53 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=2.635
+ $X2=4.56 $Y2=2.72
r138 33 35 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.56 $Y=2.635
+ $X2=4.56 $Y2=2
r139 29 50 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.72
r140 29 31 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2
r141 25 28 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.68 $Y=1.66
+ $X2=2.68 $Y2=2.34
r142 23 47 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=2.635
+ $X2=2.68 $Y2=2.72
r143 23 28 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.68 $Y=2.635
+ $X2=2.68 $Y2=2.34
r144 19 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r145 19 21 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2
r146 6 43 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.295
+ $Y=1.485 $X2=6.44 $Y2=2
r147 5 39 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.355
+ $Y=1.485 $X2=5.5 $Y2=2
r148 4 35 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.415
+ $Y=1.485 $X2=4.56 $Y2=2
r149 3 31 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.475
+ $Y=1.485 $X2=3.62 $Y2=2
r150 2 28 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=1.485 $X2=2.68 $Y2=2.34
r151 2 25 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=1.485 $X2=2.68 $Y2=1.66
r152 1 21 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_8%X 1 2 3 4 5 6 7 8 27 29 31 33 34 35 39 43 45
+ 47 51 55 57 59 63 67 72 73 75 76 79 81 82
r134 80 82 8.21116 $w=3.98e-07 $l=2.85e-07 $layer=LI1_cond $X=6.135 $Y=0.905
+ $X2=6.135 $Y2=1.19
r135 80 81 3.0006 $w=3.35e-07 $l=1.1225e-07 $layer=LI1_cond $X=6.135 $Y=0.905
+ $X2=6.085 $Y2=0.815
r136 77 82 8.78738 $w=3.98e-07 $l=3.05e-07 $layer=LI1_cond $X=6.135 $Y=1.495
+ $X2=6.135 $Y2=1.19
r137 77 79 2.63236 $w=3.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=6.135 $Y=1.495
+ $X2=6.07 $Y2=1.58
r138 65 81 3.0006 $w=3.35e-07 $l=1.53542e-07 $layer=LI1_cond $X=5.97 $Y=0.725
+ $X2=6.085 $Y2=0.815
r139 65 67 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.97 $Y=0.725
+ $X2=5.97 $Y2=0.42
r140 61 79 2.63236 $w=3.65e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.97 $Y=1.665
+ $X2=6.07 $Y2=1.58
r141 61 63 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.97 $Y=1.665
+ $X2=5.97 $Y2=2.34
r142 60 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.195 $Y=1.58
+ $X2=5.03 $Y2=1.58
r143 59 79 4.19346 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=5.805 $Y=1.58
+ $X2=6.07 $Y2=1.58
r144 59 60 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.805 $Y=1.58
+ $X2=5.195 $Y2=1.58
r145 58 76 7.13466 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=5.165 $Y=0.815
+ $X2=5.03 $Y2=0.815
r146 57 81 3.64962 $w=1.8e-07 $l=2.5e-07 $layer=LI1_cond $X=5.835 $Y=0.815
+ $X2=6.085 $Y2=0.815
r147 57 58 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=5.835 $Y=0.815
+ $X2=5.165 $Y2=0.815
r148 53 76 0.067832 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=5.03 $Y=0.725
+ $X2=5.03 $Y2=0.815
r149 53 55 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.03 $Y=0.725
+ $X2=5.03 $Y2=0.42
r150 49 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=1.665
+ $X2=5.03 $Y2=1.58
r151 49 51 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.03 $Y=1.665
+ $X2=5.03 $Y2=2.34
r152 48 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=1.58
+ $X2=4.09 $Y2=1.58
r153 47 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=1.58
+ $X2=5.03 $Y2=1.58
r154 47 48 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.865 $Y=1.58
+ $X2=4.255 $Y2=1.58
r155 46 73 7.13466 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=4.225 $Y=0.815
+ $X2=4.09 $Y2=0.815
r156 45 76 7.13466 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=4.895 $Y=0.815
+ $X2=5.03 $Y2=0.815
r157 45 46 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.895 $Y=0.815
+ $X2=4.225 $Y2=0.815
r158 41 73 0.067832 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=4.09 $Y=0.725
+ $X2=4.09 $Y2=0.815
r159 41 43 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.09 $Y=0.725
+ $X2=4.09 $Y2=0.42
r160 37 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=1.665
+ $X2=4.09 $Y2=1.58
r161 37 39 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.09 $Y=1.665
+ $X2=4.09 $Y2=2.34
r162 36 70 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=1.58
+ $X2=3.15 $Y2=1.58
r163 35 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=1.58
+ $X2=4.09 $Y2=1.58
r164 35 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.925 $Y=1.58
+ $X2=3.315 $Y2=1.58
r165 33 73 7.13466 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=3.955 $Y=0.815
+ $X2=4.09 $Y2=0.815
r166 33 34 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.955 $Y=0.815
+ $X2=3.285 $Y2=0.815
r167 29 70 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=1.665
+ $X2=3.15 $Y2=1.58
r168 29 31 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.15 $Y=1.665
+ $X2=3.15 $Y2=2.34
r169 25 34 7.38573 $w=1.8e-07 $l=1.89737e-07 $layer=LI1_cond $X=3.135 $Y=0.725
+ $X2=3.285 $Y2=0.815
r170 25 27 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=3.135 $Y=0.725
+ $X2=3.135 $Y2=0.42
r171 8 79 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.825
+ $Y=1.485 $X2=5.97 $Y2=1.66
r172 8 63 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.825
+ $Y=1.485 $X2=5.97 $Y2=2.34
r173 7 75 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.885
+ $Y=1.485 $X2=5.03 $Y2=1.66
r174 7 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.885
+ $Y=1.485 $X2=5.03 $Y2=2.34
r175 6 72 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.485 $X2=4.09 $Y2=1.66
r176 6 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.485 $X2=4.09 $Y2=2.34
r177 5 70 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=1.485 $X2=3.15 $Y2=1.66
r178 5 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=1.485 $X2=3.15 $Y2=2.34
r179 4 67 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=5.835
+ $Y=0.235 $X2=5.97 $Y2=0.42
r180 3 55 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.895
+ $Y=0.235 $X2=5.03 $Y2=0.42
r181 2 43 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.955
+ $Y=0.235 $X2=4.09 $Y2=0.42
r182 1 27 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.015
+ $Y=0.235 $X2=3.15 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_8%VGND 1 2 3 4 5 6 7 22 24 26 30 36 40 44 48
+ 52 55 56 58 59 61 62 64 65 66 82 83 89 94 103
r112 102 103 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=0.235
+ $X2=2.815 $Y2=0.235
r113 100 102 0.934436 $w=6.38e-07 $l=5e-08 $layer=LI1_cond $X=2.68 $Y=0.235
+ $X2=2.73 $Y2=0.235
r114 98 100 2.80331 $w=6.38e-07 $l=1.5e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.68 $Y2=0.235
r115 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r116 96 98 7.84926 $w=6.38e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=0.235
+ $X2=2.53 $Y2=0.235
r117 93 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r118 92 96 0.747549 $w=6.38e-07 $l=4e-08 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.11 $Y2=0.235
r119 92 94 8.17421 $w=6.38e-07 $l=4.5e-08 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.025 $Y2=0.235
r120 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r121 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r122 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r123 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r124 80 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r125 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r126 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r127 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r128 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r129 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r130 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r131 71 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r132 70 103 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=2.815 $Y2=0
r133 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r134 66 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r135 66 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r136 64 79 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.21
+ $Y2=0
r137 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.44
+ $Y2=0
r138 63 82 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=0 $X2=6.67
+ $Y2=0
r139 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=0 $X2=6.44
+ $Y2=0
r140 61 76 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.29
+ $Y2=0
r141 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.5
+ $Y2=0
r142 60 79 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.665 $Y=0
+ $X2=6.21 $Y2=0
r143 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=5.5
+ $Y2=0
r144 58 73 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.37
+ $Y2=0
r145 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.56
+ $Y2=0
r146 57 76 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.725 $Y=0 $X2=5.29
+ $Y2=0
r147 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=0 $X2=4.56
+ $Y2=0
r148 55 70 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.45
+ $Y2=0
r149 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.62
+ $Y2=0
r150 54 73 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.785 $Y=0
+ $X2=4.37 $Y2=0
r151 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.62
+ $Y2=0
r152 50 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0
r153 50 52 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0.42
r154 46 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=0.085 $X2=5.5
+ $Y2=0
r155 46 48 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.5 $Y=0.085
+ $X2=5.5 $Y2=0.42
r156 42 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0
r157 42 44 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0.42
r158 38 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0
r159 38 40 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0.42
r160 34 100 5.8233 $w=2.7e-07 $l=3.2e-07 $layer=LI1_cond $X=2.68 $Y=0.555
+ $X2=2.68 $Y2=0.235
r161 34 36 7.89637 $w=2.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.68 $Y=0.555
+ $X2=2.68 $Y2=0.74
r162 33 89 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.22
+ $Y2=0
r163 33 94 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=2.025 $Y2=0
r164 28 89 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r165 28 30 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r166 27 86 4.13993 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=0
+ $X2=0.207 $Y2=0
r167 26 89 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.085 $Y=0 $X2=1.22
+ $Y2=0
r168 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.085 $Y=0
+ $X2=0.415 $Y2=0
r169 22 86 3.14476 $w=2.7e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.207 $Y2=0
r170 22 24 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.39
r171 7 52 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=6.255
+ $Y=0.235 $X2=6.44 $Y2=0.42
r172 6 48 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=5.315
+ $Y=0.235 $X2=5.5 $Y2=0.42
r173 5 44 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.235 $X2=4.56 $Y2=0.42
r174 4 40 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=3.435
+ $Y=0.235 $X2=3.62 $Y2=0.42
r175 3 102 182 $w=1.7e-07 $l=8.24318e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.73 $Y2=0.38
r176 3 96 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.11 $Y2=0.39
r177 3 36 182 $w=1.7e-07 $l=9.75346e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.73 $Y2=0.74
r178 2 30 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
r179 1 24 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

