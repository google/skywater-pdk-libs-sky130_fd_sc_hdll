* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor2_1 A B VGND VNB VPB VPWR Y
M1000 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=6.1e+11p pd=3.22e+06u as=2.9e+11p ps=2.58e+06u
M1001 VGND A Y VNB nshort w=650000u l=150000u
+  ad=5.915e+11p pd=4.42e+06u as=1.755e+11p ps=1.84e+06u
M1002 a_117_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
