* File: sky130_fd_sc_hdll__and3_4.pxi.spice
* Created: Thu Aug 27 18:58:10 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND3_4%A N_A_c_61_n N_A_M1013_g N_A_c_62_n N_A_M1002_g A
+ A A A A N_A_c_63_n N_A_c_64_n PM_SKY130_FD_SC_HDLL__AND3_4%A
x_PM_SKY130_FD_SC_HDLL__AND3_4%B N_B_c_92_n N_B_M1001_g N_B_c_93_n N_B_M1006_g B
+ B PM_SKY130_FD_SC_HDLL__AND3_4%B
x_PM_SKY130_FD_SC_HDLL__AND3_4%C N_C_c_123_n N_C_M1007_g N_C_c_124_n N_C_M1009_g
+ C N_C_c_125_n C PM_SKY130_FD_SC_HDLL__AND3_4%C
x_PM_SKY130_FD_SC_HDLL__AND3_4%A_85_297# N_A_85_297#_M1002_s N_A_85_297#_M1013_s
+ N_A_85_297#_M1001_d N_A_85_297#_c_162_n N_A_85_297#_M1003_g
+ N_A_85_297#_c_170_n N_A_85_297#_M1000_g N_A_85_297#_c_163_n
+ N_A_85_297#_M1008_g N_A_85_297#_c_171_n N_A_85_297#_M1004_g
+ N_A_85_297#_c_164_n N_A_85_297#_M1011_g N_A_85_297#_c_172_n
+ N_A_85_297#_M1005_g N_A_85_297#_c_173_n N_A_85_297#_M1010_g
+ N_A_85_297#_c_165_n N_A_85_297#_M1012_g N_A_85_297#_c_178_n
+ N_A_85_297#_c_179_n N_A_85_297#_c_181_n N_A_85_297#_c_184_n
+ N_A_85_297#_c_194_n N_A_85_297#_c_195_n N_A_85_297#_c_207_n
+ N_A_85_297#_c_209_n N_A_85_297#_c_196_n N_A_85_297#_c_166_n
+ N_A_85_297#_c_174_n N_A_85_297#_c_175_n N_A_85_297#_c_167_n
+ N_A_85_297#_c_217_n N_A_85_297#_c_168_n N_A_85_297#_c_169_n
+ PM_SKY130_FD_SC_HDLL__AND3_4%A_85_297#
x_PM_SKY130_FD_SC_HDLL__AND3_4%VPWR N_VPWR_M1013_d N_VPWR_M1009_d N_VPWR_M1004_s
+ N_VPWR_M1010_s N_VPWR_c_306_n N_VPWR_c_307_n N_VPWR_c_308_n N_VPWR_c_309_n
+ N_VPWR_c_310_n N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_313_n VPWR
+ N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_305_n
+ PM_SKY130_FD_SC_HDLL__AND3_4%VPWR
x_PM_SKY130_FD_SC_HDLL__AND3_4%X N_X_M1003_d N_X_M1011_d N_X_M1000_d N_X_M1005_d
+ N_X_c_399_n N_X_c_373_n N_X_c_376_n N_X_c_380_n N_X_c_413_p N_X_c_403_n
+ N_X_c_382_n N_X_c_371_n N_X_c_386_n N_X_c_390_n N_X_c_392_n X N_X_c_369_n X
+ PM_SKY130_FD_SC_HDLL__AND3_4%X
x_PM_SKY130_FD_SC_HDLL__AND3_4%VGND N_VGND_M1007_d N_VGND_M1008_s N_VGND_M1012_s
+ N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n VGND N_VGND_c_439_n
+ N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n
+ PM_SKY130_FD_SC_HDLL__AND3_4%VGND
cc_1 VNB N_A_c_61_n 0.0287135f $X=-0.19 $Y=-0.24 $X2=0.825 $Y2=1.41
cc_2 VNB N_A_c_62_n 0.023905f $X=-0.19 $Y=-0.24 $X2=0.85 $Y2=0.995
cc_3 VNB N_A_c_63_n 0.00747357f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=1.16
cc_4 VNB N_A_c_64_n 0.0238471f $X=-0.19 $Y=-0.24 $X2=0.222 $Y2=1.34
cc_5 VNB N_B_c_92_n 0.0290583f $X=-0.19 $Y=-0.24 $X2=0.825 $Y2=1.41
cc_6 VNB N_B_c_93_n 0.0175624f $X=-0.19 $Y=-0.24 $X2=0.85 $Y2=0.995
cc_7 VNB B 0.00402692f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_C_c_123_n 0.0174857f $X=-0.19 $Y=-0.24 $X2=0.825 $Y2=1.41
cc_9 VNB N_C_c_124_n 0.0243152f $X=-0.19 $Y=-0.24 $X2=0.85 $Y2=0.995
cc_10 VNB N_C_c_125_n 0.00239997f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.105
cc_11 VNB N_A_85_297#_c_162_n 0.0177885f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=2.125
cc_12 VNB N_A_85_297#_c_163_n 0.016944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_85_297#_c_164_n 0.0173868f $X=-0.19 $Y=-0.24 $X2=0.222 $Y2=1.87
cc_14 VNB N_A_85_297#_c_165_n 0.0191674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_85_297#_c_166_n 0.00132882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_85_297#_c_167_n 0.0212305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_85_297#_c_168_n 0.00171227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_85_297#_c_169_n 0.0785344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_305_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_369_n 0.0127049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB X 0.0247125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_436_n 0.00504984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_437_n 0.00537481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_438_n 0.0167438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_439_n 0.0532936f $X=-0.19 $Y=-0.24 $X2=0.222 $Y2=2.21
cc_26 VNB N_VGND_c_440_n 0.012727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_441_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_442_n 0.0262989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_443_n 0.255248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VPB N_A_c_61_n 0.032369f $X=-0.19 $Y=1.305 $X2=0.825 $Y2=1.41
cc_31 VPB A 0.0529602f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_32 VPB N_A_c_63_n 0.00882125f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=1.16
cc_33 VPB N_A_c_64_n 0.00170379f $X=-0.19 $Y=1.305 $X2=0.222 $Y2=1.34
cc_34 VPB N_B_c_92_n 0.0317184f $X=-0.19 $Y=1.305 $X2=0.825 $Y2=1.41
cc_35 VPB B 0.00362357f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_36 VPB N_C_c_124_n 0.0275791f $X=-0.19 $Y=1.305 $X2=0.85 $Y2=0.995
cc_37 VPB N_C_c_125_n 0.00226523f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.105
cc_38 VPB N_A_85_297#_c_170_n 0.0166972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_85_297#_c_171_n 0.0160009f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=1.16
cc_40 VPB N_A_85_297#_c_172_n 0.0162834f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.167
cc_41 VPB N_A_85_297#_c_173_n 0.0182115f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=1.167
cc_42 VPB N_A_85_297#_c_174_n 0.00127583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_85_297#_c_175_n 0.00920717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_85_297#_c_168_n 4.55278e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_85_297#_c_169_n 0.0493244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_306_n 9.99961e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_307_n 0.0183766f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=1.16
cc_48 VPB N_VPWR_c_308_n 0.00449519f $X=-0.19 $Y=1.305 $X2=0.222 $Y2=1.53
cc_49 VPB N_VPWR_c_309_n 3.32571e-19 $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.167
cc_50 VPB N_VPWR_c_310_n 0.016009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_311_n 0.024116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_312_n 0.0168506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_313_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_314_n 0.0263363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_315_n 0.0145309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_316_n 0.00725393f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_317_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_305_n 0.0566397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_X_c_371_n 0.0166083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB X 0.0121821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 N_A_c_61_n N_B_c_92_n 0.0534161f $X=0.825 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_62 N_A_c_63_n N_B_c_92_n 3.13472e-19 $X=0.74 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_63 N_A_c_62_n N_B_c_93_n 0.0189374f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_64 N_A_c_62_n B 0.00791509f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_65 N_A_c_63_n B 0.0286461f $X=0.74 $Y=1.16 $X2=0 $Y2=0
cc_66 A N_A_85_297#_c_178_n 0.0442161f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_67 N_A_c_61_n N_A_85_297#_c_179_n 0.0203469f $X=0.825 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A_c_63_n N_A_85_297#_c_179_n 0.00938697f $X=0.74 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_c_61_n N_A_85_297#_c_181_n 5.43884e-19 $X=0.825 $Y=1.41 $X2=0 $Y2=0
cc_70 A N_A_85_297#_c_181_n 0.0142904f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_71 N_A_c_63_n N_A_85_297#_c_181_n 0.0121352f $X=0.74 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_c_62_n N_A_85_297#_c_184_n 0.0107266f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A_c_63_n N_A_85_297#_c_184_n 0.00205352f $X=0.74 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_c_61_n N_A_85_297#_c_167_n 0.0038788f $X=0.825 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_c_62_n N_A_85_297#_c_167_n 0.00814623f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A_c_63_n N_A_85_297#_c_167_n 0.0230914f $X=0.74 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_c_61_n N_VPWR_c_306_n 0.0222473f $X=0.825 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_c_61_n N_VPWR_c_314_n 0.00622633f $X=0.825 $Y=1.41 $X2=0 $Y2=0
cc_79 A N_VPWR_c_314_n 0.00834355f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_80 N_A_c_61_n N_VPWR_c_305_n 0.0116835f $X=0.825 $Y=1.41 $X2=0 $Y2=0
cc_81 A N_VPWR_c_305_n 0.00762833f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_82 N_A_c_62_n N_VGND_c_439_n 0.00357842f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_c_62_n N_VGND_c_443_n 0.00705378f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_84 N_B_c_93_n N_C_c_123_n 0.0381493f $X=1.495 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_85 N_B_c_92_n N_C_c_124_n 0.0636513f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B_c_92_n N_C_c_125_n 0.0108441f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_87 B N_C_c_125_n 0.0255313f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_88 N_B_c_92_n N_A_85_297#_c_179_n 0.0235498f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_89 B N_A_85_297#_c_179_n 0.0188821f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_90 N_B_c_92_n N_A_85_297#_c_184_n 0.00199278f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B_c_93_n N_A_85_297#_c_184_n 0.0147991f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_92 B N_A_85_297#_c_184_n 0.0144726f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_93 N_B_c_92_n N_A_85_297#_c_194_n 0.00561728f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_c_93_n N_A_85_297#_c_195_n 0.00389251f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B_c_93_n N_A_85_297#_c_196_n 0.0044884f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_96 B N_A_85_297#_c_196_n 0.00351608f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_97 N_B_c_93_n N_A_85_297#_c_167_n 0.0013259f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_98 B N_A_85_297#_c_167_n 0.00350553f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_99 N_B_c_92_n N_VPWR_c_306_n 0.0203884f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B_c_92_n N_VPWR_c_307_n 0.00642146f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B_c_92_n N_VPWR_c_305_n 0.0107572f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_102 B A_185_47# 0.0085886f $X=1.115 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_103 N_B_c_93_n N_VGND_c_439_n 0.00357877f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_104 N_B_c_93_n N_VGND_c_443_n 0.00563206f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_105 N_C_c_123_n N_A_85_297#_c_162_n 0.0161742f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_106 N_C_c_124_n N_A_85_297#_c_170_n 0.0168868f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_107 N_C_c_125_n N_A_85_297#_c_179_n 0.003649f $X=1.915 $Y=1.16 $X2=0 $Y2=0
cc_108 N_C_c_123_n N_A_85_297#_c_184_n 0.00461919f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_109 N_C_c_125_n N_A_85_297#_c_184_n 0.00254262f $X=1.915 $Y=1.16 $X2=0 $Y2=0
cc_110 N_C_c_124_n N_A_85_297#_c_194_n 0.00587833f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_111 N_C_c_123_n N_A_85_297#_c_195_n 0.00455101f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_112 N_C_c_124_n N_A_85_297#_c_207_n 0.0193873f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_113 N_C_c_125_n N_A_85_297#_c_207_n 0.0111973f $X=1.915 $Y=1.16 $X2=0 $Y2=0
cc_114 N_C_c_123_n N_A_85_297#_c_209_n 0.00888113f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_115 N_C_c_124_n N_A_85_297#_c_209_n 0.00482144f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_116 N_C_c_125_n N_A_85_297#_c_209_n 0.0131446f $X=1.915 $Y=1.16 $X2=0 $Y2=0
cc_117 N_C_c_123_n N_A_85_297#_c_196_n 0.00254166f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_118 N_C_c_125_n N_A_85_297#_c_196_n 0.0123549f $X=1.915 $Y=1.16 $X2=0 $Y2=0
cc_119 N_C_c_123_n N_A_85_297#_c_166_n 0.00382474f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_120 N_C_c_125_n N_A_85_297#_c_166_n 0.00186941f $X=1.915 $Y=1.16 $X2=0 $Y2=0
cc_121 N_C_c_124_n N_A_85_297#_c_174_n 0.00501441f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_122 N_C_c_124_n N_A_85_297#_c_217_n 5.16671e-19 $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_123 N_C_c_125_n N_A_85_297#_c_217_n 0.0115646f $X=1.915 $Y=1.16 $X2=0 $Y2=0
cc_124 N_C_c_124_n N_A_85_297#_c_168_n 0.00334719f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_125 N_C_c_125_n N_A_85_297#_c_168_n 0.0266044f $X=1.915 $Y=1.16 $X2=0 $Y2=0
cc_126 N_C_c_124_n N_A_85_297#_c_169_n 0.0151169f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_127 N_C_c_125_n N_A_85_297#_c_169_n 2.85928e-19 $X=1.915 $Y=1.16 $X2=0 $Y2=0
cc_128 N_C_c_124_n N_VPWR_c_306_n 6.1829e-19 $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_129 N_C_c_124_n N_VPWR_c_307_n 0.00702461f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_130 N_C_c_124_n N_VPWR_c_308_n 0.0018504f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_131 N_C_c_124_n N_VPWR_c_305_n 0.0126716f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_132 N_C_c_123_n N_VGND_c_436_n 0.004993f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_133 N_C_c_123_n N_VGND_c_439_n 0.00402779f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_134 N_C_c_123_n N_VGND_c_443_n 0.00599272f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_85_297#_c_179_n N_VPWR_M1013_d 0.0106296f $X=1.62 $Y=1.665 $X2=-0.19
+ $Y2=-0.24
cc_136 N_A_85_297#_c_207_n N_VPWR_M1009_d 0.00759183f $X=2.22 $Y=1.665 $X2=0
+ $Y2=0
cc_137 N_A_85_297#_c_174_n N_VPWR_M1009_d 0.00114268f $X=2.325 $Y=1.58 $X2=0
+ $Y2=0
cc_138 N_A_85_297#_c_179_n N_VPWR_c_306_n 0.0291564f $X=1.62 $Y=1.665 $X2=0
+ $Y2=0
cc_139 N_A_85_297#_c_194_n N_VPWR_c_306_n 0.0327169f $X=1.71 $Y=1.96 $X2=0 $Y2=0
cc_140 N_A_85_297#_c_194_n N_VPWR_c_307_n 0.0125171f $X=1.71 $Y=1.96 $X2=0 $Y2=0
cc_141 N_A_85_297#_c_170_n N_VPWR_c_308_n 0.00176848f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_85_297#_c_207_n N_VPWR_c_308_n 0.0209938f $X=2.22 $Y=1.665 $X2=0
+ $Y2=0
cc_143 N_A_85_297#_c_170_n N_VPWR_c_309_n 6.3373e-19 $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_144 N_A_85_297#_c_171_n N_VPWR_c_309_n 0.0137193f $X=2.985 $Y=1.41 $X2=0
+ $Y2=0
cc_145 N_A_85_297#_c_172_n N_VPWR_c_309_n 0.0102323f $X=3.465 $Y=1.41 $X2=0
+ $Y2=0
cc_146 N_A_85_297#_c_173_n N_VPWR_c_309_n 5.80987e-19 $X=3.945 $Y=1.41 $X2=0
+ $Y2=0
cc_147 N_A_85_297#_c_172_n N_VPWR_c_311_n 6.18489e-19 $X=3.465 $Y=1.41 $X2=0
+ $Y2=0
cc_148 N_A_85_297#_c_173_n N_VPWR_c_311_n 0.0146077f $X=3.945 $Y=1.41 $X2=0
+ $Y2=0
cc_149 N_A_85_297#_c_170_n N_VPWR_c_312_n 0.00702461f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_150 N_A_85_297#_c_171_n N_VPWR_c_312_n 0.00447018f $X=2.985 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_A_85_297#_c_178_n N_VPWR_c_314_n 0.0124822f $X=0.59 $Y=1.96 $X2=0 $Y2=0
cc_152 N_A_85_297#_c_172_n N_VPWR_c_315_n 0.00642146f $X=3.465 $Y=1.41 $X2=0
+ $Y2=0
cc_153 N_A_85_297#_c_173_n N_VPWR_c_315_n 0.00447018f $X=3.945 $Y=1.41 $X2=0
+ $Y2=0
cc_154 N_A_85_297#_M1013_s N_VPWR_c_305_n 0.00705085f $X=0.425 $Y=1.485 $X2=0
+ $Y2=0
cc_155 N_A_85_297#_M1001_d N_VPWR_c_305_n 0.00655879f $X=1.56 $Y=1.485 $X2=0
+ $Y2=0
cc_156 N_A_85_297#_c_170_n N_VPWR_c_305_n 0.0126606f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_157 N_A_85_297#_c_171_n N_VPWR_c_305_n 0.00766229f $X=2.985 $Y=1.41 $X2=0
+ $Y2=0
cc_158 N_A_85_297#_c_172_n N_VPWR_c_305_n 0.0107337f $X=3.465 $Y=1.41 $X2=0
+ $Y2=0
cc_159 N_A_85_297#_c_173_n N_VPWR_c_305_n 0.00766229f $X=3.945 $Y=1.41 $X2=0
+ $Y2=0
cc_160 N_A_85_297#_c_178_n N_VPWR_c_305_n 0.00684987f $X=0.59 $Y=1.96 $X2=0
+ $Y2=0
cc_161 N_A_85_297#_c_194_n N_VPWR_c_305_n 0.00685509f $X=1.71 $Y=1.96 $X2=0
+ $Y2=0
cc_162 N_A_85_297#_c_163_n N_X_c_373_n 0.0115023f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_85_297#_c_164_n N_X_c_373_n 0.0114248f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_85_297#_c_169_n N_X_c_373_n 0.00359098f $X=3.945 $Y=1.202 $X2=0 $Y2=0
cc_165 N_A_85_297#_c_171_n N_X_c_376_n 0.0175805f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_85_297#_c_172_n N_X_c_376_n 0.0168709f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_85_297#_c_175_n N_X_c_376_n 0.0480846f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_85_297#_c_169_n N_X_c_376_n 0.00161384f $X=3.945 $Y=1.202 $X2=0 $Y2=0
cc_169 N_A_85_297#_c_175_n N_X_c_380_n 0.0156439f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_85_297#_c_169_n N_X_c_380_n 0.00136562f $X=3.945 $Y=1.202 $X2=0 $Y2=0
cc_171 N_A_85_297#_c_165_n N_X_c_382_n 0.0174044f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_85_297#_c_175_n N_X_c_382_n 0.00554628f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_85_297#_c_173_n N_X_c_371_n 0.021688f $X=3.945 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_85_297#_c_175_n N_X_c_371_n 0.0056208f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_85_297#_c_209_n N_X_c_386_n 0.0135923f $X=2.22 $Y=0.71 $X2=0 $Y2=0
cc_176 N_A_85_297#_c_166_n N_X_c_386_n 0.0025314f $X=2.325 $Y=1.02 $X2=0 $Y2=0
cc_177 N_A_85_297#_c_175_n N_X_c_386_n 0.0620053f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_85_297#_c_169_n N_X_c_386_n 0.00339319f $X=3.945 $Y=1.202 $X2=0 $Y2=0
cc_179 N_A_85_297#_c_175_n N_X_c_390_n 0.0151856f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_85_297#_c_169_n N_X_c_390_n 0.00452326f $X=3.945 $Y=1.202 $X2=0 $Y2=0
cc_181 N_A_85_297#_c_175_n N_X_c_392_n 0.0156439f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_85_297#_c_169_n N_X_c_392_n 0.00136936f $X=3.945 $Y=1.202 $X2=0 $Y2=0
cc_183 N_A_85_297#_c_173_n X 0.00457136f $X=3.945 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_85_297#_c_165_n X 0.0180079f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_85_297#_c_175_n X 0.0177921f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_85_297#_c_184_n A_185_47# 0.0115399f $X=1.635 $Y=0.35 $X2=-0.19
+ $Y2=-0.24
cc_187 N_A_85_297#_c_184_n A_314_47# 0.00105457f $X=1.635 $Y=0.35 $X2=-0.19
+ $Y2=-0.24
cc_188 N_A_85_297#_c_195_n A_314_47# 0.00187568f $X=1.73 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_189 N_A_85_297#_c_196_n A_314_47# 0.00333255f $X=1.825 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_190 N_A_85_297#_c_209_n N_VGND_M1007_d 0.0111271f $X=2.22 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_191 N_A_85_297#_c_166_n N_VGND_M1007_d 0.00103313f $X=2.325 $Y=1.02 $X2=-0.19
+ $Y2=-0.24
cc_192 N_A_85_297#_c_162_n N_VGND_c_436_n 0.00192556f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_193 N_A_85_297#_c_184_n N_VGND_c_436_n 0.0123921f $X=1.635 $Y=0.35 $X2=0
+ $Y2=0
cc_194 N_A_85_297#_c_209_n N_VGND_c_436_n 0.0232062f $X=2.22 $Y=0.71 $X2=0 $Y2=0
cc_195 N_A_85_297#_c_162_n N_VGND_c_437_n 0.00108514f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_85_297#_c_163_n N_VGND_c_437_n 0.00842193f $X=2.96 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_85_297#_c_164_n N_VGND_c_437_n 0.00685144f $X=3.44 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_85_297#_c_165_n N_VGND_c_437_n 4.66497e-19 $X=3.97 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_85_297#_c_162_n N_VGND_c_438_n 0.00558147f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_85_297#_c_163_n N_VGND_c_438_n 0.0035176f $X=2.96 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_85_297#_c_209_n N_VGND_c_438_n 6.66898e-19 $X=2.22 $Y=0.71 $X2=0
+ $Y2=0
cc_202 N_A_85_297#_c_184_n N_VGND_c_439_n 0.0589979f $X=1.635 $Y=0.35 $X2=0
+ $Y2=0
cc_203 N_A_85_297#_c_209_n N_VGND_c_439_n 0.00363772f $X=2.22 $Y=0.71 $X2=0
+ $Y2=0
cc_204 N_A_85_297#_c_167_n N_VGND_c_439_n 0.0211961f $X=0.635 $Y=0.38 $X2=0
+ $Y2=0
cc_205 N_A_85_297#_c_164_n N_VGND_c_440_n 0.0035176f $X=3.44 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_85_297#_c_165_n N_VGND_c_440_n 0.00210367f $X=3.97 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_85_297#_c_164_n N_VGND_c_442_n 5.14844e-19 $X=3.44 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_85_297#_c_165_n N_VGND_c_442_n 0.0103132f $X=3.97 $Y=0.995 $X2=0
+ $Y2=0
cc_209 N_A_85_297#_M1002_s N_VGND_c_443_n 0.0024621f $X=0.47 $Y=0.235 $X2=0
+ $Y2=0
cc_210 N_A_85_297#_c_162_n N_VGND_c_443_n 0.0103473f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_85_297#_c_163_n N_VGND_c_443_n 0.00424616f $X=2.96 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_A_85_297#_c_164_n N_VGND_c_443_n 0.00431085f $X=3.44 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_85_297#_c_165_n N_VGND_c_443_n 0.00294796f $X=3.97 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A_85_297#_c_184_n N_VGND_c_443_n 0.0369861f $X=1.635 $Y=0.35 $X2=0
+ $Y2=0
cc_215 N_A_85_297#_c_209_n N_VGND_c_443_n 0.00898191f $X=2.22 $Y=0.71 $X2=0
+ $Y2=0
cc_216 N_A_85_297#_c_167_n N_VGND_c_443_n 0.0126448f $X=0.635 $Y=0.38 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_305_n N_X_M1000_d 0.00621163f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_c_305_n N_X_M1005_d 0.00621163f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_c_312_n N_X_c_399_n 0.0131506f $X=3.01 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_c_305_n N_X_c_399_n 0.00722976f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_221 N_VPWR_M1004_s N_X_c_376_n 0.00364629f $X=3.075 $Y=1.485 $X2=0 $Y2=0
cc_222 N_VPWR_c_309_n N_X_c_376_n 0.0209288f $X=3.225 $Y=2.02 $X2=0 $Y2=0
cc_223 N_VPWR_c_315_n N_X_c_403_n 0.0131506f $X=3.97 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_c_305_n N_X_c_403_n 0.00722976f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_M1010_s N_X_c_371_n 0.00866677f $X=4.035 $Y=1.485 $X2=0 $Y2=0
cc_226 N_VPWR_c_311_n N_X_c_371_n 0.0272529f $X=4.185 $Y=2.02 $X2=0 $Y2=0
cc_227 N_VPWR_M1010_s X 9.17578e-19 $X=4.035 $Y=1.485 $X2=0 $Y2=0
cc_228 N_X_c_373_n N_VGND_M1008_s 0.00421224f $X=3.61 $Y=0.73 $X2=0 $Y2=0
cc_229 N_X_c_382_n N_VGND_M1012_s 0.00533494f $X=4.21 $Y=0.73 $X2=0 $Y2=0
cc_230 N_X_c_369_n N_VGND_M1012_s 0.00260919f $X=4.35 $Y=0.845 $X2=0 $Y2=0
cc_231 X N_VGND_M1012_s 7.05546e-19 $X=4.345 $Y=0.85 $X2=0 $Y2=0
cc_232 N_X_c_373_n N_VGND_c_437_n 0.0200941f $X=3.61 $Y=0.73 $X2=0 $Y2=0
cc_233 N_X_c_413_p N_VGND_c_437_n 0.0117256f $X=3.705 $Y=0.42 $X2=0 $Y2=0
cc_234 N_X_c_373_n N_VGND_c_438_n 0.00264153f $X=3.61 $Y=0.73 $X2=0 $Y2=0
cc_235 N_X_c_386_n N_VGND_c_438_n 0.00449666f $X=2.84 $Y=0.68 $X2=0 $Y2=0
cc_236 N_X_c_373_n N_VGND_c_440_n 0.00346656f $X=3.61 $Y=0.73 $X2=0 $Y2=0
cc_237 N_X_c_413_p N_VGND_c_440_n 0.0130838f $X=3.705 $Y=0.42 $X2=0 $Y2=0
cc_238 N_X_c_382_n N_VGND_c_440_n 0.00258244f $X=4.21 $Y=0.73 $X2=0 $Y2=0
cc_239 N_X_c_413_p N_VGND_c_442_n 0.014372f $X=3.705 $Y=0.42 $X2=0 $Y2=0
cc_240 N_X_c_382_n N_VGND_c_442_n 0.013705f $X=4.21 $Y=0.73 $X2=0 $Y2=0
cc_241 N_X_c_369_n N_VGND_c_442_n 0.0147598f $X=4.35 $Y=0.845 $X2=0 $Y2=0
cc_242 N_X_M1003_d N_VGND_c_443_n 0.00648119f $X=2.555 $Y=0.235 $X2=0 $Y2=0
cc_243 N_X_M1011_d N_VGND_c_443_n 0.00368069f $X=3.515 $Y=0.235 $X2=0 $Y2=0
cc_244 N_X_c_373_n N_VGND_c_443_n 0.0118634f $X=3.61 $Y=0.73 $X2=0 $Y2=0
cc_245 N_X_c_413_p N_VGND_c_443_n 0.00721345f $X=3.705 $Y=0.42 $X2=0 $Y2=0
cc_246 N_X_c_382_n N_VGND_c_443_n 0.00561718f $X=4.21 $Y=0.73 $X2=0 $Y2=0
cc_247 N_X_c_386_n N_VGND_c_443_n 0.00604783f $X=2.84 $Y=0.68 $X2=0 $Y2=0
cc_248 N_X_c_369_n N_VGND_c_443_n 0.00500503f $X=4.35 $Y=0.845 $X2=0 $Y2=0
cc_249 A_185_47# N_VGND_c_443_n 0.00399797f $X=0.925 $Y=0.235 $X2=0 $Y2=0
cc_250 A_314_47# N_VGND_c_443_n 0.00168634f $X=1.57 $Y=0.235 $X2=0.68 $Y2=1.665
