* File: sky130_fd_sc_hdll__dlrtp_1.pxi.spice
* Created: Wed Sep  2 08:29:32 2020
* 
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%GATE N_GATE_c_138_n N_GATE_c_139_n
+ N_GATE_M1001_g N_GATE_c_133_n N_GATE_M1014_g N_GATE_c_134_n GATE GATE
+ N_GATE_c_136_n N_GATE_c_137_n PM_SKY130_FD_SC_HDLL__DLRTP_1%GATE
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%A_27_363# N_A_27_363#_M1014_s
+ N_A_27_363#_M1001_s N_A_27_363#_M1002_g N_A_27_363#_c_185_n
+ N_A_27_363#_M1016_g N_A_27_363#_c_186_n N_A_27_363#_c_187_n
+ N_A_27_363#_M1017_g N_A_27_363#_c_176_n N_A_27_363#_M1005_g
+ N_A_27_363#_c_189_n N_A_27_363#_c_321_p N_A_27_363#_c_178_n
+ N_A_27_363#_c_179_n N_A_27_363#_c_190_n N_A_27_363#_c_191_n
+ N_A_27_363#_c_180_n N_A_27_363#_c_181_n N_A_27_363#_c_193_n
+ N_A_27_363#_c_194_n N_A_27_363#_c_195_n N_A_27_363#_c_241_p
+ N_A_27_363#_c_182_n N_A_27_363#_c_183_n N_A_27_363#_c_184_n
+ PM_SKY130_FD_SC_HDLL__DLRTP_1%A_27_363#
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%D N_D_c_334_n N_D_c_335_n N_D_M1008_g
+ N_D_M1007_g N_D_c_331_n N_D_c_332_n D PM_SKY130_FD_SC_HDLL__DLRTP_1%D
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%A_319_369# N_A_319_369#_M1007_s
+ N_A_319_369#_M1008_s N_A_319_369#_c_373_n N_A_319_369#_c_379_n
+ N_A_319_369#_M1004_g N_A_319_369#_M1018_g N_A_319_369#_c_380_n
+ N_A_319_369#_c_374_n N_A_319_369#_c_382_n N_A_319_369#_c_375_n
+ N_A_319_369#_c_376_n N_A_319_369#_c_377_n
+ PM_SKY130_FD_SC_HDLL__DLRTP_1%A_319_369#
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%A_203_47# N_A_203_47#_M1002_d
+ N_A_203_47#_M1016_d N_A_203_47#_M1010_g N_A_203_47#_c_456_n
+ N_A_203_47#_M1015_g N_A_203_47#_c_452_n N_A_203_47#_c_453_n
+ N_A_203_47#_c_459_n N_A_203_47#_c_454_n N_A_203_47#_c_455_n
+ N_A_203_47#_c_460_n N_A_203_47#_c_461_n N_A_203_47#_c_462_n
+ N_A_203_47#_c_533_p N_A_203_47#_c_463_n
+ PM_SKY130_FD_SC_HDLL__DLRTP_1%A_203_47#
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%A_750_21# N_A_750_21#_M1013_s
+ N_A_750_21#_M1019_d N_A_750_21#_M1000_g N_A_750_21#_c_570_n
+ N_A_750_21#_M1003_g N_A_750_21#_c_571_n N_A_750_21#_M1011_g
+ N_A_750_21#_c_572_n N_A_750_21#_M1006_g N_A_750_21#_c_579_n
+ N_A_750_21#_c_573_n N_A_750_21#_c_574_n N_A_750_21#_c_594_p
+ N_A_750_21#_c_619_p N_A_750_21#_c_581_n N_A_750_21#_c_575_n
+ N_A_750_21#_c_591_p N_A_750_21#_c_576_n
+ PM_SKY130_FD_SC_HDLL__DLRTP_1%A_750_21#
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%A_604_47# N_A_604_47#_M1010_d
+ N_A_604_47#_M1017_d N_A_604_47#_c_669_n N_A_604_47#_c_677_n
+ N_A_604_47#_M1019_g N_A_604_47#_M1013_g N_A_604_47#_c_671_n
+ N_A_604_47#_c_682_n N_A_604_47#_c_683_n N_A_604_47#_c_672_n
+ N_A_604_47#_c_679_n N_A_604_47#_c_673_n N_A_604_47#_c_674_n
+ N_A_604_47#_c_675_n PM_SKY130_FD_SC_HDLL__DLRTP_1%A_604_47#
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%RESET_B N_RESET_B_c_762_n N_RESET_B_M1009_g
+ N_RESET_B_c_763_n N_RESET_B_M1012_g RESET_B
+ PM_SKY130_FD_SC_HDLL__DLRTP_1%RESET_B
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%VPWR N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_M1003_d N_VPWR_M1012_d N_VPWR_c_795_n N_VPWR_c_796_n N_VPWR_c_797_n
+ N_VPWR_c_853_n N_VPWR_c_798_n N_VPWR_c_799_n VPWR N_VPWR_c_800_n
+ N_VPWR_c_801_n N_VPWR_c_802_n N_VPWR_c_803_n N_VPWR_c_794_n N_VPWR_c_805_n
+ N_VPWR_c_806_n N_VPWR_c_807_n PM_SKY130_FD_SC_HDLL__DLRTP_1%VPWR
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%Q N_Q_M1011_d N_Q_M1006_d N_Q_c_891_n
+ N_Q_c_893_n N_Q_c_894_n N_Q_c_895_n Q PM_SKY130_FD_SC_HDLL__DLRTP_1%Q
x_PM_SKY130_FD_SC_HDLL__DLRTP_1%VGND N_VGND_M1014_d N_VGND_M1007_d
+ N_VGND_M1000_d N_VGND_M1009_d N_VGND_c_914_n N_VGND_c_915_n N_VGND_c_916_n
+ N_VGND_c_917_n N_VGND_c_918_n N_VGND_c_919_n N_VGND_c_974_n VGND
+ N_VGND_c_920_n N_VGND_c_921_n N_VGND_c_922_n N_VGND_c_923_n N_VGND_c_924_n
+ N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n
+ PM_SKY130_FD_SC_HDLL__DLRTP_1%VGND
cc_1 VNB N_GATE_c_133_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_2 VNB N_GATE_c_134_n 0.0254358f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_3 VNB GATE 0.0176317f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_GATE_c_136_n 0.0192744f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.235
cc_5 VNB N_GATE_c_137_n 0.0161691f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.07
cc_6 VNB N_A_27_363#_M1002_g 0.0390164f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_7 VNB N_A_27_363#_c_176_n 0.0132521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_363#_M1005_g 0.0385424f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.235
cc_9 VNB N_A_27_363#_c_178_n 0.00122303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_363#_c_179_n 0.00595335f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_363#_c_180_n 0.00288001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_363#_c_181_n 0.00401055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_363#_c_182_n 0.0215048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_363#_c_183_n 0.00964173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_363#_c_184_n 0.00774225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1007_g 0.0323122f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_17 VNB N_D_c_331_n 0.0294428f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_18 VNB N_D_c_332_n 0.0116306f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=0.805
cc_19 VNB D 0.0122424f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_319_369#_c_373_n 0.0137191f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_21 VNB N_A_319_369#_c_374_n 0.00197693f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_22 VNB N_A_319_369#_c_375_n 0.0140494f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_23 VNB N_A_319_369#_c_376_n 0.0231274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_319_369#_c_377_n 0.0172162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_203_47#_M1010_g 0.0200544f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_26 VNB N_A_203_47#_c_452_n 0.0143934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_203_47#_c_453_n 0.00362448f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_28 VNB N_A_203_47#_c_454_n 0.0267668f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.235
cc_29 VNB N_A_203_47#_c_455_n 0.00955011f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.07
cc_30 VNB N_A_750_21#_M1000_g 0.0440056f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_31 VNB N_A_750_21#_c_570_n 0.00267512f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=0.805
cc_32 VNB N_A_750_21#_c_571_n 0.0214386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_750_21#_c_572_n 0.0241266f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_34 VNB N_A_750_21#_c_573_n 0.00461115f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_35 VNB N_A_750_21#_c_574_n 0.00473847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_750_21#_c_575_n 0.00314085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_750_21#_c_576_n 0.0045085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_604_47#_c_669_n 0.0116996f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_39 VNB N_A_604_47#_M1013_g 0.0273327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_604_47#_c_671_n 0.00540275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_604_47#_c_672_n 0.00311441f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_42 VNB N_A_604_47#_c_673_n 0.0089303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_604_47#_c_674_n 0.00336267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_604_47#_c_675_n 0.0289378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_c_762_n 0.0169297f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=0.88
cc_46 VNB N_RESET_B_c_763_n 0.0197191f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.59
cc_47 VNB RESET_B 0.0100492f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_48 VNB N_VPWR_c_794_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_Q_c_891_n 0.0348014f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_50 VNB Q 0.0215011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_914_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.665
cc_52 VNB N_VGND_c_915_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_53 VNB N_VGND_c_916_n 0.00703343f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.235
cc_54 VNB N_VGND_c_917_n 0.00525786f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_55 VNB N_VGND_c_918_n 0.0323621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_919_n 0.00528586f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_57 VNB N_VGND_c_920_n 0.0167943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_921_n 0.0299753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_922_n 0.03956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_923_n 0.0236451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_924_n 0.347955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_925_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_926_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_927_n 0.00507956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VPB N_GATE_c_138_n 0.0140771f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.59
cc_66 VPB N_GATE_c_139_n 0.0453152f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_67 VPB GATE 0.0133135f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_68 VPB N_GATE_c_136_n 0.00895075f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.235
cc_69 VPB N_A_27_363#_c_185_n 0.0315264f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_70 VPB N_A_27_363#_c_186_n 0.0136262f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_71 VPB N_A_27_363#_c_187_n 0.0232482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_363#_c_176_n 0.0170551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_363#_c_189_n 0.0141256f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_74 VPB N_A_27_363#_c_190_n 2.97507e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_363#_c_191_n 0.0311637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_363#_c_180_n 0.00156054f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_363#_c_193_n 0.018179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_363#_c_194_n 0.00382566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_363#_c_195_n 0.00508133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_363#_c_182_n 0.01105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_363#_c_183_n 0.0231911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_363#_c_184_n 0.00381159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_D_c_334_n 0.0219771f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.07
cc_84 VPB N_D_c_335_n 0.0271128f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.4
cc_85 VPB N_D_c_331_n 0.0118988f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_86 VPB N_D_c_332_n 6.82386e-19 $X=-0.19 $Y=1.305 $X2=0.33 $Y2=0.805
cc_87 VPB D 0.00308729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_319_369#_c_373_n 0.0175584f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_89 VPB N_A_319_369#_c_379_n 0.0233198f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_90 VPB N_A_319_369#_c_380_n 0.00818123f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_91 VPB N_A_319_369#_c_374_n 0.00137236f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_92 VPB N_A_319_369#_c_382_n 0.00599855f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.235
cc_93 VPB N_A_203_47#_c_456_n 0.0478596f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=0.805
cc_94 VPB N_A_203_47#_c_452_n 0.00835207f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_203_47#_c_453_n 0.00298141f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_96 VPB N_A_203_47#_c_459_n 0.00412793f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_97 VPB N_A_203_47#_c_460_n 0.00977716f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_98 VPB N_A_203_47#_c_461_n 9.68792e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_203_47#_c_462_n 0.00684047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_203_47#_c_463_n 0.00859475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_750_21#_c_570_n 0.0882876f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=0.805
cc_102 VPB N_A_750_21#_c_572_n 0.0294676f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_103 VPB N_A_750_21#_c_579_n 0.0031059f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_104 VPB N_A_750_21#_c_574_n 0.00223949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_750_21#_c_581_n 0.00166281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_750_21#_c_576_n 0.00149364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_604_47#_c_669_n 0.00770302f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_108 VPB N_A_604_47#_c_677_n 0.0198076f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_109 VPB N_A_604_47#_c_671_n 0.00700495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_604_47#_c_679_n 0.0052925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_604_47#_c_674_n 0.00167692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_604_47#_c_675_n 0.00663603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_RESET_B_c_763_n 0.0246089f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.59
cc_114 VPB RESET_B 0.00222063f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_115 VPB N_VPWR_c_795_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.665
cc_116 VPB N_VPWR_c_796_n 0.0083008f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_117 VPB N_VPWR_c_797_n 0.00264814f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.235
cc_118 VPB N_VPWR_c_798_n 0.0187301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_799_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_120 VPB N_VPWR_c_800_n 0.0157721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_801_n 0.0302711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_802_n 0.0481942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_803_n 0.0226788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_794_n 0.0546256f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_805_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_806_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_807_n 0.0183527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_Q_c_893_n 0.0110377f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.665
cc_129 VPB N_Q_c_894_n 0.0251921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_Q_c_895_n 0.00902941f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_131 VPB Q 0.00962814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 N_GATE_c_133_n N_A_27_363#_M1002_g 0.0188581f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_133 N_GATE_c_137_n N_A_27_363#_M1002_g 0.00431579f $X=0.3 $Y=1.07 $X2=0 $Y2=0
cc_134 N_GATE_c_139_n N_A_27_363#_c_185_n 0.0246962f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_135 N_GATE_c_136_n N_A_27_363#_c_189_n 0.00509098f $X=0.3 $Y=1.235 $X2=0
+ $Y2=0
cc_136 N_GATE_c_133_n N_A_27_363#_c_178_n 0.00683119f $X=0.52 $Y=0.73 $X2=0
+ $Y2=0
cc_137 N_GATE_c_134_n N_A_27_363#_c_178_n 0.00844637f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_138 GATE N_A_27_363#_c_178_n 0.00279004f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_139 N_GATE_c_134_n N_A_27_363#_c_179_n 0.0084549f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_140 GATE N_A_27_363#_c_179_n 0.0134132f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_141 N_GATE_c_139_n N_A_27_363#_c_190_n 0.0149414f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_142 GATE N_A_27_363#_c_190_n 0.00295527f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_143 N_GATE_c_139_n N_A_27_363#_c_191_n 0.005546f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_144 GATE N_A_27_363#_c_191_n 0.0280207f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_145 N_GATE_c_136_n N_A_27_363#_c_191_n 2.83366e-19 $X=0.3 $Y=1.235 $X2=0
+ $Y2=0
cc_146 N_GATE_c_136_n N_A_27_363#_c_180_n 0.00208392f $X=0.3 $Y=1.235 $X2=0
+ $Y2=0
cc_147 N_GATE_c_134_n N_A_27_363#_c_181_n 0.00194152f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_148 GATE N_A_27_363#_c_181_n 0.0470252f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_149 N_GATE_c_137_n N_A_27_363#_c_181_n 0.00208392f $X=0.3 $Y=1.07 $X2=0 $Y2=0
cc_150 N_GATE_c_138_n N_A_27_363#_c_194_n 0.00359932f $X=0.33 $Y=1.59 $X2=0
+ $Y2=0
cc_151 N_GATE_c_139_n N_A_27_363#_c_194_n 0.0019946f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_152 N_GATE_c_134_n N_A_27_363#_c_194_n 7.30071e-19 $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_153 GATE N_A_27_363#_c_194_n 0.00696823f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_154 N_GATE_c_138_n N_A_27_363#_c_195_n 0.00208392f $X=0.33 $Y=1.59 $X2=0
+ $Y2=0
cc_155 N_GATE_c_139_n N_A_27_363#_c_195_n 0.00455102f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_156 GATE N_A_27_363#_c_182_n 3.1077e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_157 N_GATE_c_136_n N_A_27_363#_c_182_n 0.0166463f $X=0.3 $Y=1.235 $X2=0 $Y2=0
cc_158 N_GATE_c_139_n N_VPWR_c_795_n 0.00923594f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_159 N_GATE_c_139_n N_VPWR_c_800_n 0.0044329f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_160 N_GATE_c_139_n N_VPWR_c_794_n 0.00608656f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_161 N_GATE_c_133_n N_VGND_c_914_n 0.00913236f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_162 N_GATE_c_133_n N_VGND_c_920_n 0.00339367f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_163 N_GATE_c_134_n N_VGND_c_920_n 5.87962e-19 $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_164 N_GATE_c_133_n N_VGND_c_924_n 0.00502432f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_165 N_A_27_363#_c_193_n N_D_c_334_n 0.0041274f $X=2.665 $Y=1.53 $X2=0 $Y2=0
cc_166 N_A_27_363#_c_184_n N_D_c_334_n 3.09224e-19 $X=2.87 $Y=1.44 $X2=0 $Y2=0
cc_167 N_A_27_363#_M1002_g N_D_c_331_n 0.00692544f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_27_363#_c_193_n N_D_c_331_n 0.00222839f $X=2.665 $Y=1.53 $X2=0 $Y2=0
cc_169 N_A_27_363#_c_184_n N_D_c_332_n 2.52874e-19 $X=2.87 $Y=1.44 $X2=0 $Y2=0
cc_170 N_A_27_363#_c_193_n D 0.0112094f $X=2.665 $Y=1.53 $X2=0 $Y2=0
cc_171 N_A_27_363#_c_186_n N_A_319_369#_c_373_n 0.00540817f $X=2.95 $Y=1.89
+ $X2=0 $Y2=0
cc_172 N_A_27_363#_c_193_n N_A_319_369#_c_373_n 0.00352657f $X=2.665 $Y=1.53
+ $X2=0 $Y2=0
cc_173 N_A_27_363#_c_183_n N_A_319_369#_c_373_n 0.0253968f $X=2.892 $Y=1.32
+ $X2=0 $Y2=0
cc_174 N_A_27_363#_c_184_n N_A_319_369#_c_373_n 0.0118476f $X=2.87 $Y=1.44 $X2=0
+ $Y2=0
cc_175 N_A_27_363#_c_186_n N_A_319_369#_c_379_n 0.00877513f $X=2.95 $Y=1.89
+ $X2=0 $Y2=0
cc_176 N_A_27_363#_c_187_n N_A_319_369#_c_379_n 0.0230867f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_177 N_A_27_363#_c_184_n N_A_319_369#_c_379_n 0.0018263f $X=2.87 $Y=1.44 $X2=0
+ $Y2=0
cc_178 N_A_27_363#_c_193_n N_A_319_369#_c_380_n 4.87587e-19 $X=2.665 $Y=1.53
+ $X2=0 $Y2=0
cc_179 N_A_27_363#_c_184_n N_A_319_369#_c_380_n 5.53168e-19 $X=2.87 $Y=1.44
+ $X2=0 $Y2=0
cc_180 N_A_27_363#_c_193_n N_A_319_369#_c_374_n 0.0111584f $X=2.665 $Y=1.53
+ $X2=0 $Y2=0
cc_181 N_A_27_363#_c_241_p N_A_319_369#_c_374_n 2.15582e-19 $X=2.81 $Y=1.53
+ $X2=0 $Y2=0
cc_182 N_A_27_363#_c_184_n N_A_319_369#_c_374_n 0.0101463f $X=2.87 $Y=1.44 $X2=0
+ $Y2=0
cc_183 N_A_27_363#_c_193_n N_A_319_369#_c_382_n 0.0178505f $X=2.665 $Y=1.53
+ $X2=0 $Y2=0
cc_184 N_A_27_363#_c_241_p N_A_319_369#_c_382_n 2.48695e-19 $X=2.81 $Y=1.53
+ $X2=0 $Y2=0
cc_185 N_A_27_363#_c_184_n N_A_319_369#_c_382_n 0.0065905f $X=2.87 $Y=1.44 $X2=0
+ $Y2=0
cc_186 N_A_27_363#_c_193_n N_A_319_369#_c_375_n 0.0126321f $X=2.665 $Y=1.53
+ $X2=0 $Y2=0
cc_187 N_A_27_363#_c_184_n N_A_319_369#_c_375_n 0.00654622f $X=2.87 $Y=1.44
+ $X2=0 $Y2=0
cc_188 N_A_27_363#_M1005_g N_A_203_47#_M1010_g 0.00922459f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_189 N_A_27_363#_c_186_n N_A_203_47#_c_456_n 0.0053733f $X=2.95 $Y=1.89 $X2=0
+ $Y2=0
cc_190 N_A_27_363#_c_187_n N_A_203_47#_c_456_n 0.0112656f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_191 N_A_27_363#_c_176_n N_A_203_47#_c_456_n 0.018099f $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_192 N_A_27_363#_c_183_n N_A_203_47#_c_456_n 0.016719f $X=2.892 $Y=1.32 $X2=0
+ $Y2=0
cc_193 N_A_27_363#_M1002_g N_A_203_47#_c_452_n 0.0177545f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_A_27_363#_c_185_n N_A_203_47#_c_452_n 0.00400552f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_195 N_A_27_363#_c_178_n N_A_203_47#_c_452_n 0.00911803f $X=0.605 $Y=0.72
+ $X2=0 $Y2=0
cc_196 N_A_27_363#_c_180_n N_A_203_47#_c_452_n 0.024482f $X=0.81 $Y=1.235 $X2=0
+ $Y2=0
cc_197 N_A_27_363#_c_181_n N_A_203_47#_c_452_n 0.0136901f $X=0.75 $Y=1.07 $X2=0
+ $Y2=0
cc_198 N_A_27_363#_c_193_n N_A_203_47#_c_452_n 0.0189902f $X=2.665 $Y=1.53 $X2=0
+ $Y2=0
cc_199 N_A_27_363#_c_194_n N_A_203_47#_c_452_n 0.00256031f $X=0.835 $Y=1.53
+ $X2=0 $Y2=0
cc_200 N_A_27_363#_c_195_n N_A_203_47#_c_452_n 0.0173414f $X=0.69 $Y=1.53 $X2=0
+ $Y2=0
cc_201 N_A_27_363#_c_176_n N_A_203_47#_c_453_n 0.012296f $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_202 N_A_27_363#_M1005_g N_A_203_47#_c_453_n 0.00335377f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_203 N_A_27_363#_c_241_p N_A_203_47#_c_453_n 0.00446852f $X=2.81 $Y=1.53 $X2=0
+ $Y2=0
cc_204 N_A_27_363#_c_183_n N_A_203_47#_c_453_n 0.00411158f $X=2.892 $Y=1.32
+ $X2=0 $Y2=0
cc_205 N_A_27_363#_c_184_n N_A_203_47#_c_453_n 0.0212936f $X=2.87 $Y=1.44 $X2=0
+ $Y2=0
cc_206 N_A_27_363#_c_185_n N_A_203_47#_c_459_n 0.00241063f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_207 N_A_27_363#_c_190_n N_A_203_47#_c_459_n 0.00552354f $X=0.605 $Y=1.88
+ $X2=0 $Y2=0
cc_208 N_A_27_363#_c_193_n N_A_203_47#_c_459_n 0.0035784f $X=2.665 $Y=1.53 $X2=0
+ $Y2=0
cc_209 N_A_27_363#_M1005_g N_A_203_47#_c_454_n 0.0121069f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_210 N_A_27_363#_c_183_n N_A_203_47#_c_454_n 0.0211774f $X=2.892 $Y=1.32 $X2=0
+ $Y2=0
cc_211 N_A_27_363#_c_176_n N_A_203_47#_c_455_n 8.98998e-19 $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_212 N_A_27_363#_M1005_g N_A_203_47#_c_455_n 0.00357812f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_213 N_A_27_363#_c_241_p N_A_203_47#_c_455_n 9.8074e-19 $X=2.81 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_27_363#_c_183_n N_A_203_47#_c_455_n 0.00551002f $X=2.892 $Y=1.32
+ $X2=0 $Y2=0
cc_215 N_A_27_363#_c_184_n N_A_203_47#_c_455_n 0.0132372f $X=2.87 $Y=1.44 $X2=0
+ $Y2=0
cc_216 N_A_27_363#_c_186_n N_A_203_47#_c_460_n 0.005923f $X=2.95 $Y=1.89 $X2=0
+ $Y2=0
cc_217 N_A_27_363#_c_187_n N_A_203_47#_c_460_n 0.00405726f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_218 N_A_27_363#_c_176_n N_A_203_47#_c_460_n 0.00138393f $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_219 N_A_27_363#_c_193_n N_A_203_47#_c_460_n 0.104184f $X=2.665 $Y=1.53 $X2=0
+ $Y2=0
cc_220 N_A_27_363#_c_241_p N_A_203_47#_c_460_n 0.0261499f $X=2.81 $Y=1.53 $X2=0
+ $Y2=0
cc_221 N_A_27_363#_c_184_n N_A_203_47#_c_460_n 0.0156538f $X=2.87 $Y=1.44 $X2=0
+ $Y2=0
cc_222 N_A_27_363#_c_185_n N_A_203_47#_c_461_n 0.00182829f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_223 N_A_27_363#_c_190_n N_A_203_47#_c_461_n 0.00529043f $X=0.605 $Y=1.88
+ $X2=0 $Y2=0
cc_224 N_A_27_363#_c_193_n N_A_203_47#_c_461_n 0.025576f $X=2.665 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_27_363#_c_195_n N_A_203_47#_c_461_n 9.19894e-19 $X=0.69 $Y=1.53 $X2=0
+ $Y2=0
cc_226 N_A_27_363#_c_176_n N_A_203_47#_c_463_n 0.00558349f $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_227 N_A_27_363#_c_241_p N_A_203_47#_c_463_n 0.00182791f $X=2.81 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_363#_c_183_n N_A_203_47#_c_463_n 0.00863156f $X=2.892 $Y=1.32
+ $X2=0 $Y2=0
cc_229 N_A_27_363#_c_184_n N_A_203_47#_c_463_n 0.00800041f $X=2.87 $Y=1.44 $X2=0
+ $Y2=0
cc_230 N_A_27_363#_M1005_g N_A_750_21#_M1000_g 0.0394664f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_231 N_A_27_363#_c_176_n N_A_750_21#_c_570_n 0.0394664f $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_232 N_A_27_363#_c_183_n N_A_750_21#_c_570_n 2.81272e-19 $X=2.892 $Y=1.32
+ $X2=0 $Y2=0
cc_233 N_A_27_363#_c_187_n N_A_604_47#_c_682_n 0.00515668f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_234 N_A_27_363#_c_176_n N_A_604_47#_c_683_n 0.00138963f $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_235 N_A_27_363#_M1005_g N_A_604_47#_c_683_n 0.0113891f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_236 N_A_27_363#_M1005_g N_A_604_47#_c_672_n 0.00872448f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_237 N_A_27_363#_c_176_n N_A_604_47#_c_679_n 6.06088e-19 $X=3.39 $Y=1.32 $X2=0
+ $Y2=0
cc_238 N_A_27_363#_c_183_n N_A_604_47#_c_679_n 4.18131e-19 $X=2.892 $Y=1.32
+ $X2=0 $Y2=0
cc_239 N_A_27_363#_M1005_g N_A_604_47#_c_673_n 0.0061787f $X=3.465 $Y=0.445
+ $X2=0 $Y2=0
cc_240 N_A_27_363#_c_190_n N_VPWR_M1001_d 0.00298278f $X=0.605 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_241 N_A_27_363#_c_185_n N_VPWR_c_795_n 0.009458f $X=0.965 $Y=1.74 $X2=0 $Y2=0
cc_242 N_A_27_363#_c_190_n N_VPWR_c_795_n 0.0124663f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_243 N_A_27_363#_c_191_n N_VPWR_c_795_n 0.0127533f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_244 N_A_27_363#_c_193_n N_VPWR_c_795_n 0.00196536f $X=2.665 $Y=1.53 $X2=0
+ $Y2=0
cc_245 N_A_27_363#_c_194_n N_VPWR_c_795_n 0.00327384f $X=0.835 $Y=1.53 $X2=0
+ $Y2=0
cc_246 N_A_27_363#_c_193_n N_VPWR_c_796_n 0.00140184f $X=2.665 $Y=1.53 $X2=0
+ $Y2=0
cc_247 N_A_27_363#_c_190_n N_VPWR_c_800_n 0.00206959f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_248 N_A_27_363#_c_191_n N_VPWR_c_800_n 0.0220573f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_249 N_A_27_363#_c_185_n N_VPWR_c_801_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_250 N_A_27_363#_c_187_n N_VPWR_c_802_n 0.00694986f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_251 N_A_27_363#_c_185_n N_VPWR_c_794_n 0.0113647f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_252 N_A_27_363#_c_187_n N_VPWR_c_794_n 0.00771671f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_253 N_A_27_363#_c_190_n N_VPWR_c_794_n 0.00444188f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_254 N_A_27_363#_c_191_n N_VPWR_c_794_n 0.011857f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_255 N_A_27_363#_c_178_n N_VGND_M1014_d 0.00151978f $X=0.605 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_256 N_A_27_363#_M1002_g N_VGND_c_914_n 0.00953934f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_257 N_A_27_363#_c_178_n N_VGND_c_914_n 0.0123958f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_258 N_A_27_363#_c_180_n N_VGND_c_914_n 0.0028901f $X=0.81 $Y=1.235 $X2=0
+ $Y2=0
cc_259 N_A_27_363#_c_182_n N_VGND_c_914_n 6.85506e-19 $X=0.94 $Y=1.235 $X2=0
+ $Y2=0
cc_260 N_A_27_363#_M1005_g N_VGND_c_916_n 0.0016369f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_261 N_A_27_363#_c_321_p N_VGND_c_920_n 0.00981821f $X=0.31 $Y=0.445 $X2=0
+ $Y2=0
cc_262 N_A_27_363#_c_178_n N_VGND_c_920_n 0.00243651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_263 N_A_27_363#_M1002_g N_VGND_c_921_n 0.0046653f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_264 N_A_27_363#_M1005_g N_VGND_c_922_n 0.00362991f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_265 N_A_27_363#_M1014_s N_VGND_c_924_n 0.00366338f $X=0.185 $Y=0.235 $X2=0
+ $Y2=0
cc_266 N_A_27_363#_M1002_g N_VGND_c_924_n 0.00934473f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_267 N_A_27_363#_M1005_g N_VGND_c_924_n 0.00539993f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_268 N_A_27_363#_c_321_p N_VGND_c_924_n 0.00634536f $X=0.31 $Y=0.445 $X2=0
+ $Y2=0
cc_269 N_A_27_363#_c_178_n N_VGND_c_924_n 0.00525284f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_270 N_D_c_332_n N_A_319_369#_c_373_n 0.0154881f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_271 N_D_c_334_n N_A_319_369#_c_379_n 0.0154881f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_272 N_D_c_335_n N_A_319_369#_c_379_n 0.009841f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_273 N_D_c_335_n N_A_319_369#_c_380_n 0.0134542f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_274 N_D_c_334_n N_A_319_369#_c_374_n 0.00821507f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_275 N_D_c_332_n N_A_319_369#_c_374_n 0.00663872f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_276 D N_A_319_369#_c_374_n 0.0156567f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_277 N_D_c_334_n N_A_319_369#_c_382_n 0.0121171f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_278 N_D_c_331_n N_A_319_369#_c_382_n 0.00443823f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_279 D N_A_319_369#_c_382_n 0.0138356f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_280 N_D_M1007_g N_A_319_369#_c_375_n 0.0222419f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_281 N_D_c_331_n N_A_319_369#_c_375_n 0.00632987f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_282 N_D_c_332_n N_A_319_369#_c_375_n 0.00343492f $X=1.955 $Y=1.16 $X2=0 $Y2=0
cc_283 D N_A_319_369#_c_375_n 0.0196854f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_284 N_D_M1007_g N_A_319_369#_c_376_n 0.0213174f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_285 N_D_M1007_g N_A_319_369#_c_377_n 0.0138443f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_286 N_D_c_334_n N_A_203_47#_c_452_n 0.00403725f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_287 N_D_M1007_g N_A_203_47#_c_452_n 0.00569292f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_288 N_D_c_331_n N_A_203_47#_c_452_n 0.00112186f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_289 D N_A_203_47#_c_452_n 0.0261672f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_290 N_D_c_335_n N_A_203_47#_c_459_n 0.00144922f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_291 N_D_c_335_n N_A_203_47#_c_460_n 0.00409389f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_292 N_D_c_335_n N_VPWR_c_796_n 0.00329547f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_293 N_D_c_335_n N_VPWR_c_801_n 0.00673617f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_294 N_D_c_335_n N_VPWR_c_794_n 0.00835409f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_295 N_D_M1007_g N_VGND_c_915_n 0.0111499f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_296 N_D_M1007_g N_VGND_c_921_n 0.00336882f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_297 N_D_M1007_g N_VGND_c_924_n 0.00532348f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_298 N_A_319_369#_c_377_n N_A_203_47#_M1010_g 0.0220789f $X=2.4 $Y=0.765 $X2=0
+ $Y2=0
cc_299 N_A_319_369#_c_380_n N_A_203_47#_c_452_n 9.98908e-19 $X=1.72 $Y=1.99
+ $X2=0 $Y2=0
cc_300 N_A_319_369#_c_382_n N_A_203_47#_c_452_n 0.00743802f $X=2.03 $Y=1.58
+ $X2=0 $Y2=0
cc_301 N_A_319_369#_c_375_n N_A_203_47#_c_452_n 0.0173676f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_302 N_A_319_369#_c_373_n N_A_203_47#_c_453_n 0.00350056f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_303 N_A_319_369#_c_380_n N_A_203_47#_c_459_n 0.0502658f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_304 N_A_319_369#_c_375_n N_A_203_47#_c_454_n 3.43721e-19 $X=2.03 $Y=0.72
+ $X2=0 $Y2=0
cc_305 N_A_319_369#_c_376_n N_A_203_47#_c_454_n 0.0144623f $X=2.4 $Y=0.93 $X2=0
+ $Y2=0
cc_306 N_A_319_369#_c_377_n N_A_203_47#_c_454_n 0.00124411f $X=2.4 $Y=0.765
+ $X2=0 $Y2=0
cc_307 N_A_319_369#_c_375_n N_A_203_47#_c_455_n 0.0212212f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_308 N_A_319_369#_c_376_n N_A_203_47#_c_455_n 7.77092e-19 $X=2.4 $Y=0.93 $X2=0
+ $Y2=0
cc_309 N_A_319_369#_c_379_n N_A_203_47#_c_460_n 0.00677393f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_310 N_A_319_369#_c_380_n N_A_203_47#_c_460_n 0.0211788f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_311 N_A_319_369#_c_382_n N_A_203_47#_c_460_n 0.00465602f $X=2.03 $Y=1.58
+ $X2=0 $Y2=0
cc_312 N_A_319_369#_c_380_n N_A_203_47#_c_461_n 0.00257398f $X=1.72 $Y=1.99
+ $X2=0 $Y2=0
cc_313 N_A_319_369#_c_379_n N_A_203_47#_c_463_n 3.59161e-19 $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_314 N_A_319_369#_c_379_n N_A_604_47#_c_682_n 9.84369e-19 $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_315 N_A_319_369#_c_379_n N_VPWR_c_796_n 0.00422565f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_316 N_A_319_369#_c_380_n N_VPWR_c_796_n 0.025165f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_317 N_A_319_369#_c_382_n N_VPWR_c_796_n 0.00394172f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_318 N_A_319_369#_c_380_n N_VPWR_c_801_n 0.0210596f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_319 N_A_319_369#_c_379_n N_VPWR_c_802_n 0.00702461f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_320 N_A_319_369#_M1008_s N_VPWR_c_794_n 0.00179197f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_321 N_A_319_369#_c_379_n N_VPWR_c_794_n 0.0074238f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_322 N_A_319_369#_c_380_n N_VPWR_c_794_n 0.00594162f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_323 N_A_319_369#_c_375_n N_VGND_M1007_d 5.4803e-19 $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_324 N_A_319_369#_c_375_n N_VGND_c_915_n 0.0120795f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_325 N_A_319_369#_c_376_n N_VGND_c_915_n 3.80743e-19 $X=2.4 $Y=0.93 $X2=0
+ $Y2=0
cc_326 N_A_319_369#_c_377_n N_VGND_c_915_n 0.00798806f $X=2.4 $Y=0.765 $X2=0
+ $Y2=0
cc_327 N_A_319_369#_c_375_n N_VGND_c_921_n 0.0109521f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_328 N_A_319_369#_c_376_n N_VGND_c_922_n 2.5317e-19 $X=2.4 $Y=0.93 $X2=0 $Y2=0
cc_329 N_A_319_369#_c_377_n N_VGND_c_922_n 0.00564095f $X=2.4 $Y=0.765 $X2=0
+ $Y2=0
cc_330 N_A_319_369#_M1007_s N_VGND_c_924_n 0.00285324f $X=1.645 $Y=0.235 $X2=0
+ $Y2=0
cc_331 N_A_319_369#_c_375_n N_VGND_c_924_n 0.0189897f $X=2.03 $Y=0.72 $X2=0
+ $Y2=0
cc_332 N_A_319_369#_c_377_n N_VGND_c_924_n 0.00527362f $X=2.4 $Y=0.765 $X2=0
+ $Y2=0
cc_333 N_A_203_47#_c_456_n N_A_750_21#_c_570_n 0.0476997f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_334 N_A_203_47#_c_453_n N_A_750_21#_c_570_n 8.26114e-19 $X=3.21 $Y=1.575
+ $X2=0 $Y2=0
cc_335 N_A_203_47#_c_463_n N_A_750_21#_c_570_n 6.27988e-19 $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_336 N_A_203_47#_c_456_n N_A_604_47#_c_682_n 0.0127286f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_337 N_A_203_47#_c_460_n N_A_604_47#_c_682_n 0.00338792f $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_338 N_A_203_47#_c_533_p N_A_604_47#_c_682_n 0.00120815f $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_339 N_A_203_47#_c_463_n N_A_604_47#_c_682_n 0.02443f $X=3.365 $Y=1.87 $X2=0
+ $Y2=0
cc_340 N_A_203_47#_c_454_n N_A_604_47#_c_683_n 0.00146696f $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_341 N_A_203_47#_c_455_n N_A_604_47#_c_683_n 0.0182656f $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_342 N_A_203_47#_M1010_g N_A_604_47#_c_672_n 7.58363e-19 $X=2.945 $Y=0.415
+ $X2=0 $Y2=0
cc_343 N_A_203_47#_c_454_n N_A_604_47#_c_672_n 2.13323e-19 $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_344 N_A_203_47#_c_455_n N_A_604_47#_c_672_n 0.0183748f $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_345 N_A_203_47#_c_456_n N_A_604_47#_c_679_n 0.0059256f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_346 N_A_203_47#_c_453_n N_A_604_47#_c_679_n 0.0104035f $X=3.21 $Y=1.575 $X2=0
+ $Y2=0
cc_347 N_A_203_47#_c_533_p N_A_604_47#_c_679_n 0.0017055f $X=3.365 $Y=1.87 $X2=0
+ $Y2=0
cc_348 N_A_203_47#_c_463_n N_A_604_47#_c_679_n 0.0290753f $X=3.365 $Y=1.87 $X2=0
+ $Y2=0
cc_349 N_A_203_47#_c_456_n N_A_604_47#_c_673_n 0.00178452f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_350 N_A_203_47#_c_453_n N_A_604_47#_c_673_n 0.012389f $X=3.21 $Y=1.575 $X2=0
+ $Y2=0
cc_351 N_A_203_47#_c_455_n N_A_604_47#_c_673_n 0.00778088f $X=3.21 $Y=0.915
+ $X2=0 $Y2=0
cc_352 N_A_203_47#_c_463_n N_A_604_47#_c_673_n 7.63243e-19 $X=3.365 $Y=1.87
+ $X2=0 $Y2=0
cc_353 N_A_203_47#_c_460_n N_VPWR_M1008_d 2.27104e-19 $X=3.22 $Y=1.87 $X2=0
+ $Y2=0
cc_354 N_A_203_47#_c_462_n N_VPWR_c_795_n 0.0127456f $X=1.2 $Y=1.87 $X2=0 $Y2=0
cc_355 N_A_203_47#_c_460_n N_VPWR_c_796_n 0.0196711f $X=3.22 $Y=1.87 $X2=0 $Y2=0
cc_356 N_A_203_47#_c_462_n N_VPWR_c_801_n 0.0192143f $X=1.2 $Y=1.87 $X2=0 $Y2=0
cc_357 N_A_203_47#_c_456_n N_VPWR_c_802_n 0.00448856f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_358 N_A_203_47#_c_456_n N_VPWR_c_794_n 0.00609959f $X=3.42 $Y=1.99 $X2=0
+ $Y2=0
cc_359 N_A_203_47#_c_460_n N_VPWR_c_794_n 0.0902341f $X=3.22 $Y=1.87 $X2=0 $Y2=0
cc_360 N_A_203_47#_c_461_n N_VPWR_c_794_n 0.0147801f $X=1.345 $Y=1.87 $X2=0
+ $Y2=0
cc_361 N_A_203_47#_c_462_n N_VPWR_c_794_n 0.00468601f $X=1.2 $Y=1.87 $X2=0 $Y2=0
cc_362 N_A_203_47#_c_533_p N_VPWR_c_794_n 0.0144105f $X=3.365 $Y=1.87 $X2=0
+ $Y2=0
cc_363 N_A_203_47#_c_460_n A_503_369# 0.00369043f $X=3.22 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_364 N_A_203_47#_M1010_g N_VGND_c_915_n 0.00181512f $X=2.945 $Y=0.415 $X2=0
+ $Y2=0
cc_365 N_A_203_47#_c_452_n N_VGND_c_921_n 0.00999887f $X=1.15 $Y=0.445 $X2=0
+ $Y2=0
cc_366 N_A_203_47#_M1010_g N_VGND_c_922_n 0.00439206f $X=2.945 $Y=0.415 $X2=0
+ $Y2=0
cc_367 N_A_203_47#_c_454_n N_VGND_c_922_n 0.00155706f $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_368 N_A_203_47#_c_455_n N_VGND_c_922_n 0.00358349f $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_369 N_A_203_47#_M1002_d N_VGND_c_924_n 0.00530224f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_370 N_A_203_47#_M1010_g N_VGND_c_924_n 0.00664952f $X=2.945 $Y=0.415 $X2=0
+ $Y2=0
cc_371 N_A_203_47#_c_452_n N_VGND_c_924_n 0.00639171f $X=1.15 $Y=0.445 $X2=0
+ $Y2=0
cc_372 N_A_203_47#_c_454_n N_VGND_c_924_n 0.00259944f $X=2.945 $Y=0.9 $X2=0
+ $Y2=0
cc_373 N_A_203_47#_c_455_n N_VGND_c_924_n 0.00661169f $X=3.21 $Y=0.915 $X2=0
+ $Y2=0
cc_374 N_A_750_21#_c_574_n N_A_604_47#_c_669_n 0.010664f $X=4.635 $Y=1.535 $X2=0
+ $Y2=0
cc_375 N_A_750_21#_c_575_n N_A_604_47#_c_669_n 0.00309332f $X=4.62 $Y=0.825
+ $X2=0 $Y2=0
cc_376 N_A_750_21#_c_591_p N_A_604_47#_c_669_n 6.70661e-19 $X=5.17 $Y=1.7 $X2=0
+ $Y2=0
cc_377 N_A_750_21#_c_570_n N_A_604_47#_c_677_n 0.01028f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_378 N_A_750_21#_c_574_n N_A_604_47#_c_677_n 0.00421619f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_379 N_A_750_21#_c_594_p N_A_604_47#_c_677_n 0.0154481f $X=5.04 $Y=1.96 $X2=0
+ $Y2=0
cc_380 N_A_750_21#_c_591_p N_A_604_47#_c_677_n 0.0234551f $X=5.17 $Y=1.7 $X2=0
+ $Y2=0
cc_381 N_A_750_21#_c_573_n N_A_604_47#_M1013_g 0.00740647f $X=4.62 $Y=0.38 $X2=0
+ $Y2=0
cc_382 N_A_750_21#_c_574_n N_A_604_47#_M1013_g 0.00577472f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_383 N_A_750_21#_c_575_n N_A_604_47#_M1013_g 0.00435148f $X=4.62 $Y=0.825
+ $X2=0 $Y2=0
cc_384 N_A_750_21#_c_574_n N_A_604_47#_c_671_n 0.00545235f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_385 N_A_750_21#_c_570_n N_A_604_47#_c_682_n 0.00613606f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_386 N_A_750_21#_M1000_g N_A_604_47#_c_683_n 0.00206262f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_387 N_A_750_21#_M1000_g N_A_604_47#_c_672_n 0.00870159f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_388 N_A_750_21#_c_570_n N_A_604_47#_c_679_n 0.03553f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_389 N_A_750_21#_c_579_n N_A_604_47#_c_679_n 0.0246758f $X=4.55 $Y=1.7 $X2=0
+ $Y2=0
cc_390 N_A_750_21#_M1000_g N_A_604_47#_c_673_n 0.00970956f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_391 N_A_750_21#_c_570_n N_A_604_47#_c_673_n 6.43776e-19 $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_392 N_A_750_21#_M1000_g N_A_604_47#_c_674_n 0.00591896f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_393 N_A_750_21#_c_570_n N_A_604_47#_c_674_n 0.0129533f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_394 N_A_750_21#_c_579_n N_A_604_47#_c_674_n 0.0239061f $X=4.55 $Y=1.7 $X2=0
+ $Y2=0
cc_395 N_A_750_21#_c_574_n N_A_604_47#_c_674_n 0.0256838f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_396 N_A_750_21#_M1000_g N_A_604_47#_c_675_n 0.0138805f $X=3.825 $Y=0.445
+ $X2=0 $Y2=0
cc_397 N_A_750_21#_c_570_n N_A_604_47#_c_675_n 0.00935438f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_398 N_A_750_21#_c_579_n N_A_604_47#_c_675_n 0.00919786f $X=4.55 $Y=1.7 $X2=0
+ $Y2=0
cc_399 N_A_750_21#_c_574_n N_A_604_47#_c_675_n 0.00131564f $X=4.635 $Y=1.535
+ $X2=0 $Y2=0
cc_400 N_A_750_21#_c_571_n N_RESET_B_c_762_n 0.0100656f $X=5.72 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_401 N_A_750_21#_c_573_n N_RESET_B_c_762_n 0.00167884f $X=4.62 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_402 N_A_750_21#_c_572_n N_RESET_B_c_763_n 0.0460168f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_403 N_A_750_21#_c_574_n N_RESET_B_c_763_n 9.44656e-19 $X=4.635 $Y=1.535 $X2=0
+ $Y2=0
cc_404 N_A_750_21#_c_619_p N_RESET_B_c_763_n 0.0149373f $X=5.555 $Y=1.62 $X2=0
+ $Y2=0
cc_405 N_A_750_21#_c_581_n N_RESET_B_c_763_n 0.00427849f $X=5.64 $Y=1.535 $X2=0
+ $Y2=0
cc_406 N_A_750_21#_c_591_p N_RESET_B_c_763_n 0.00125633f $X=5.17 $Y=1.7 $X2=0
+ $Y2=0
cc_407 N_A_750_21#_c_576_n N_RESET_B_c_763_n 8.84866e-19 $X=5.73 $Y=1.16 $X2=0
+ $Y2=0
cc_408 N_A_750_21#_c_572_n RESET_B 7.27155e-19 $X=5.745 $Y=1.41 $X2=0 $Y2=0
cc_409 N_A_750_21#_c_574_n RESET_B 0.0249612f $X=4.635 $Y=1.535 $X2=0 $Y2=0
cc_410 N_A_750_21#_c_591_p RESET_B 0.0278573f $X=5.17 $Y=1.7 $X2=0 $Y2=0
cc_411 N_A_750_21#_c_576_n RESET_B 0.0221162f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_412 N_A_750_21#_c_579_n N_VPWR_M1003_d 0.00479992f $X=4.55 $Y=1.7 $X2=0 $Y2=0
cc_413 N_A_750_21#_c_574_n N_VPWR_M1003_d 0.00115467f $X=4.635 $Y=1.535 $X2=0
+ $Y2=0
cc_414 N_A_750_21#_c_591_p N_VPWR_M1003_d 0.00188621f $X=5.17 $Y=1.7 $X2=0 $Y2=0
cc_415 N_A_750_21#_c_619_p N_VPWR_M1012_d 0.00694156f $X=5.555 $Y=1.62 $X2=0
+ $Y2=0
cc_416 N_A_750_21#_c_581_n N_VPWR_M1012_d 5.76203e-19 $X=5.64 $Y=1.535 $X2=0
+ $Y2=0
cc_417 N_A_750_21#_c_572_n N_VPWR_c_797_n 0.00312368f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_418 N_A_750_21#_c_572_n N_VPWR_c_853_n 0.0040108f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_419 N_A_750_21#_c_619_p N_VPWR_c_853_n 0.0165281f $X=5.555 $Y=1.62 $X2=0
+ $Y2=0
cc_420 N_A_750_21#_c_594_p N_VPWR_c_798_n 0.0163168f $X=5.04 $Y=1.96 $X2=0 $Y2=0
cc_421 N_A_750_21#_c_570_n N_VPWR_c_802_n 0.00667791f $X=3.9 $Y=1.99 $X2=0 $Y2=0
cc_422 N_A_750_21#_c_572_n N_VPWR_c_803_n 0.00652041f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_423 N_A_750_21#_M1019_d N_VPWR_c_794_n 0.0027906f $X=4.895 $Y=1.485 $X2=0
+ $Y2=0
cc_424 N_A_750_21#_c_570_n N_VPWR_c_794_n 0.0138324f $X=3.9 $Y=1.99 $X2=0 $Y2=0
cc_425 N_A_750_21#_c_572_n N_VPWR_c_794_n 0.0121842f $X=5.745 $Y=1.41 $X2=0
+ $Y2=0
cc_426 N_A_750_21#_c_579_n N_VPWR_c_794_n 0.00331262f $X=4.55 $Y=1.7 $X2=0 $Y2=0
cc_427 N_A_750_21#_c_594_p N_VPWR_c_794_n 0.0107499f $X=5.04 $Y=1.96 $X2=0 $Y2=0
cc_428 N_A_750_21#_c_591_p N_VPWR_c_794_n 0.00781507f $X=5.17 $Y=1.7 $X2=0 $Y2=0
cc_429 N_A_750_21#_c_570_n N_VPWR_c_807_n 0.0128891f $X=3.9 $Y=1.99 $X2=0 $Y2=0
cc_430 N_A_750_21#_c_579_n N_VPWR_c_807_n 0.0325801f $X=4.55 $Y=1.7 $X2=0 $Y2=0
cc_431 N_A_750_21#_c_594_p N_VPWR_c_807_n 0.0197406f $X=5.04 $Y=1.96 $X2=0 $Y2=0
cc_432 N_A_750_21#_c_571_n N_Q_c_891_n 0.00356318f $X=5.72 $Y=0.995 $X2=0 $Y2=0
cc_433 N_A_750_21#_c_572_n N_Q_c_891_n 0.00109067f $X=5.745 $Y=1.41 $X2=0 $Y2=0
cc_434 N_A_750_21#_c_576_n N_Q_c_891_n 0.00591221f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_435 N_A_750_21#_c_572_n N_Q_c_893_n 0.00317976f $X=5.745 $Y=1.41 $X2=0 $Y2=0
cc_436 N_A_750_21#_c_619_p N_Q_c_895_n 0.0141663f $X=5.555 $Y=1.62 $X2=0 $Y2=0
cc_437 N_A_750_21#_c_581_n N_Q_c_895_n 0.00297249f $X=5.64 $Y=1.535 $X2=0 $Y2=0
cc_438 N_A_750_21#_c_571_n Q 0.00189777f $X=5.72 $Y=0.995 $X2=0 $Y2=0
cc_439 N_A_750_21#_c_572_n Q 0.00651033f $X=5.745 $Y=1.41 $X2=0 $Y2=0
cc_440 N_A_750_21#_c_581_n Q 0.00523671f $X=5.64 $Y=1.535 $X2=0 $Y2=0
cc_441 N_A_750_21#_c_576_n Q 0.0218704f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_442 N_A_750_21#_M1000_g N_VGND_c_916_n 0.0114443f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_443 N_A_750_21#_c_573_n N_VGND_c_916_n 0.0222896f $X=4.62 $Y=0.38 $X2=0 $Y2=0
cc_444 N_A_750_21#_c_571_n N_VGND_c_917_n 0.00291966f $X=5.72 $Y=0.995 $X2=0
+ $Y2=0
cc_445 N_A_750_21#_c_573_n N_VGND_c_918_n 0.0209274f $X=4.62 $Y=0.38 $X2=0 $Y2=0
cc_446 N_A_750_21#_c_571_n N_VGND_c_974_n 0.00184845f $X=5.72 $Y=0.995 $X2=0
+ $Y2=0
cc_447 N_A_750_21#_c_576_n N_VGND_c_974_n 0.00412626f $X=5.73 $Y=1.16 $X2=0
+ $Y2=0
cc_448 N_A_750_21#_M1000_g N_VGND_c_922_n 0.0046653f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_A_750_21#_c_571_n N_VGND_c_923_n 0.00535523f $X=5.72 $Y=0.995 $X2=0
+ $Y2=0
cc_450 N_A_750_21#_M1013_s N_VGND_c_924_n 0.00209319f $X=4.495 $Y=0.235 $X2=0
+ $Y2=0
cc_451 N_A_750_21#_M1000_g N_VGND_c_924_n 0.00783311f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_452 N_A_750_21#_c_571_n N_VGND_c_924_n 0.010628f $X=5.72 $Y=0.995 $X2=0 $Y2=0
cc_453 N_A_750_21#_c_573_n N_VGND_c_924_n 0.0123993f $X=4.62 $Y=0.38 $X2=0 $Y2=0
cc_454 N_A_604_47#_M1013_g N_RESET_B_c_762_n 0.0427931f $X=4.83 $Y=0.56
+ $X2=-0.19 $Y2=-0.24
cc_455 N_A_604_47#_c_677_n N_RESET_B_c_763_n 0.00946913f $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_456 N_A_604_47#_M1013_g N_RESET_B_c_763_n 0.0213675f $X=4.83 $Y=0.56 $X2=0
+ $Y2=0
cc_457 N_A_604_47#_c_671_n N_RESET_B_c_763_n 0.00398928f $X=4.805 $Y=1.25 $X2=0
+ $Y2=0
cc_458 N_A_604_47#_M1013_g RESET_B 0.00402529f $X=4.83 $Y=0.56 $X2=0 $Y2=0
cc_459 N_A_604_47#_c_671_n RESET_B 0.00387184f $X=4.805 $Y=1.25 $X2=0 $Y2=0
cc_460 N_A_604_47#_c_677_n N_VPWR_c_797_n 9.88682e-19 $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_461 N_A_604_47#_c_677_n N_VPWR_c_798_n 0.00688798f $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_462 N_A_604_47#_c_682_n N_VPWR_c_802_n 0.0311316f $X=3.68 $Y=2.275 $X2=0
+ $Y2=0
cc_463 N_A_604_47#_M1017_d N_VPWR_c_794_n 0.00194144f $X=3.04 $Y=2.065 $X2=0
+ $Y2=0
cc_464 N_A_604_47#_c_677_n N_VPWR_c_794_n 0.00859707f $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_465 N_A_604_47#_c_682_n N_VPWR_c_794_n 0.0194526f $X=3.68 $Y=2.275 $X2=0
+ $Y2=0
cc_466 N_A_604_47#_c_677_n N_VPWR_c_807_n 0.00662978f $X=4.805 $Y=1.41 $X2=0
+ $Y2=0
cc_467 N_A_604_47#_c_682_n N_VPWR_c_807_n 0.0166799f $X=3.68 $Y=2.275 $X2=0
+ $Y2=0
cc_468 N_A_604_47#_c_679_n N_VPWR_c_807_n 0.00202439f $X=3.765 $Y=2.165 $X2=0
+ $Y2=0
cc_469 N_A_604_47#_c_682_n A_702_413# 0.00588737f $X=3.68 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_470 N_A_604_47#_c_679_n A_702_413# 0.00114824f $X=3.765 $Y=2.165 $X2=-0.19
+ $Y2=-0.24
cc_471 N_A_604_47#_M1013_g N_VGND_c_916_n 0.00210532f $X=4.83 $Y=0.56 $X2=0
+ $Y2=0
cc_472 N_A_604_47#_c_683_n N_VGND_c_916_n 0.0198459f $X=3.49 $Y=0.422 $X2=0
+ $Y2=0
cc_473 N_A_604_47#_c_672_n N_VGND_c_916_n 0.00279232f $X=3.575 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_604_47#_c_674_n N_VGND_c_916_n 0.0141331f $X=4.295 $Y=1.16 $X2=0
+ $Y2=0
cc_475 N_A_604_47#_c_675_n N_VGND_c_916_n 7.94156e-19 $X=4.295 $Y=1.16 $X2=0
+ $Y2=0
cc_476 N_A_604_47#_M1013_g N_VGND_c_918_n 0.00541359f $X=4.83 $Y=0.56 $X2=0
+ $Y2=0
cc_477 N_A_604_47#_c_683_n N_VGND_c_922_n 0.0313331f $X=3.49 $Y=0.422 $X2=0
+ $Y2=0
cc_478 N_A_604_47#_M1010_d N_VGND_c_924_n 0.0030893f $X=3.02 $Y=0.235 $X2=0
+ $Y2=0
cc_479 N_A_604_47#_M1013_g N_VGND_c_924_n 0.0110154f $X=4.83 $Y=0.56 $X2=0 $Y2=0
cc_480 N_A_604_47#_c_683_n N_VGND_c_924_n 0.0224738f $X=3.49 $Y=0.422 $X2=0
+ $Y2=0
cc_481 N_A_604_47#_c_683_n A_708_47# 0.0032618f $X=3.49 $Y=0.422 $X2=-0.19
+ $Y2=-0.24
cc_482 N_A_604_47#_c_672_n A_708_47# 8.90683e-19 $X=3.575 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_483 N_RESET_B_c_763_n N_VPWR_c_797_n 0.00821098f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_484 N_RESET_B_c_763_n N_VPWR_c_853_n 0.00308687f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_485 N_RESET_B_c_763_n N_VPWR_c_798_n 0.00622633f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_486 N_RESET_B_c_763_n N_VPWR_c_794_n 0.0104264f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_487 N_RESET_B_c_762_n N_VGND_c_917_n 0.00315649f $X=5.235 $Y=0.995 $X2=0
+ $Y2=0
cc_488 N_RESET_B_c_762_n N_VGND_c_918_n 0.00585385f $X=5.235 $Y=0.995 $X2=0
+ $Y2=0
cc_489 N_RESET_B_c_763_n N_VGND_c_974_n 0.00153517f $X=5.275 $Y=1.41 $X2=0 $Y2=0
cc_490 RESET_B N_VGND_c_974_n 0.00322068f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_491 N_RESET_B_c_762_n N_VGND_c_924_n 0.0106807f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_492 N_VPWR_c_794_n A_503_369# 0.00493898f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_493 N_VPWR_c_794_n A_702_413# 0.00249044f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_494 N_VPWR_c_794_n N_Q_M1006_d 0.00217517f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_495 N_VPWR_c_803_n N_Q_c_893_n 0.0317008f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_496 N_VPWR_c_794_n N_Q_c_893_n 0.0181675f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_497 N_VPWR_c_853_n N_Q_c_894_n 0.0171288f $X=5.51 $Y=1.97 $X2=0 $Y2=0
cc_498 N_Q_c_891_n N_VGND_c_923_n 0.0352943f $X=6.18 $Y=0.885 $X2=0 $Y2=0
cc_499 N_Q_M1011_d N_VGND_c_924_n 0.00209319f $X=5.795 $Y=0.235 $X2=0 $Y2=0
cc_500 N_Q_c_891_n N_VGND_c_924_n 0.0201325f $X=6.18 $Y=0.885 $X2=0 $Y2=0
cc_501 N_VGND_c_924_n A_500_47# 0.0121316f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_502 N_VGND_c_924_n A_708_47# 0.00481582f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_503 N_VGND_c_924_n A_981_47# 0.0109001f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
