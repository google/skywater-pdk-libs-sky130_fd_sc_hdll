# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__conb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.605000 1.740000 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775000 0.915000 1.295000 2.465000 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.275000  1.910000 0.605000 2.635000 ;
      RECT 0.775000  0.085000 1.115000 0.745000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__conb_1
END LIBRARY
