* File: sky130_fd_sc_hdll__bufbuf_8.pex.spice
* Created: Thu Aug 27 19:00:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_8%A 1 3 6 8
c27 8 0 1.49267e-19 $X=0.235 $Y=1.19
r28 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r29 4 11 40.1292 $w=4.26e-07 $l=2.36525e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.352 $Y2=1.16
r30 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r31 1 11 44.7281 $w=4.26e-07 $l=3.13449e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.352 $Y2=1.16
r32 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_8%A_27_47# 1 2 7 9 10 12 15 19 21 22 23 24
+ 27
c63 23 0 1.38193e-19 $X=0.66 $Y=1.53
c64 7 0 1.49267e-19 $X=1.03 $Y=1.41
r65 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.005
+ $Y=1.16 $X2=1.005 $Y2=1.16
r66 23 27 15.7832 $w=2.86e-07 $l=4.75079e-07 $layer=LI1_cond $X=0.66 $Y=1.53
+ $X2=0.9 $Y2=1.16
r67 23 24 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.66 $Y=1.53
+ $X2=0.425 $Y2=1.53
r68 21 27 14.5035 $w=2.86e-07 $l=4.44072e-07 $layer=LI1_cond $X=0.66 $Y=0.82
+ $X2=0.9 $Y2=1.16
r69 21 22 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.66 $Y=0.82
+ $X2=0.425 $Y2=0.82
r70 17 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.425 $Y2=1.53
r71 17 19 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.63
r72 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.425 $Y2=0.82
r73 13 15 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.47
r74 10 28 38.5336 $w=3.07e-07 $l=1.80748e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.022 $Y2=1.16
r75 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=0.56
r76 7 28 47.4309 $w=3.07e-07 $l=2.53969e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.022 $Y2=1.16
r77 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41 $X2=1.03
+ $Y2=1.985
r78 2 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r79 1 15 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_8%A_224_297# 1 2 9 11 13 16 18 20 21 23 26
+ 30 33 38 42 46 47 48 54
c105 38 0 1.39726e-19 $X=2.625 $Y=1.16
c106 26 0 1.25206e-19 $X=3.015 $Y=0.56
c107 21 0 1.26528e-19 $X=2.99 $Y=1.41
r108 54 55 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.99 $Y=1.217
+ $X2=3.015 $Y2=1.217
r109 51 52 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.495 $Y=1.217
+ $X2=2.52 $Y2=1.217
r110 50 51 64.997 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=2.05 $Y=1.217
+ $X2=2.495 $Y2=1.217
r111 49 50 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.025 $Y=1.217
+ $X2=2.05 $Y2=1.217
r112 46 47 6.64081 $w=4.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=1.63
+ $X2=1.265 $Y2=1.545
r113 42 44 15.7532 $w=4.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.265 $Y=0.4
+ $X2=1.265 $Y2=0.825
r114 39 54 53.3121 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.625 $Y=1.217
+ $X2=2.99 $Y2=1.217
r115 39 52 15.3364 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=2.625 $Y=1.217
+ $X2=2.52 $Y2=1.217
r116 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.625
+ $Y=1.16 $X2=2.625 $Y2=1.16
r117 36 48 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=1.175
+ $X2=1.395 $Y2=1.175
r118 36 38 63.4955 $w=1.98e-07 $l=1.145e-06 $layer=LI1_cond $X=1.48 $Y=1.175
+ $X2=2.625 $Y2=1.175
r119 34 48 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.395 $Y=1.275
+ $X2=1.395 $Y2=1.175
r120 34 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.395 $Y=1.275
+ $X2=1.395 $Y2=1.545
r121 33 48 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.395 $Y=1.075
+ $X2=1.395 $Y2=1.175
r122 33 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.395 $Y=1.075
+ $X2=1.395 $Y2=0.825
r123 28 46 3.48413 $w=4.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.265 $Y=1.76
+ $X2=1.265 $Y2=1.63
r124 28 30 14.7406 $w=4.28e-07 $l=5.5e-07 $layer=LI1_cond $X=1.265 $Y=1.76
+ $X2=1.265 $Y2=2.31
r125 24 55 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.015 $Y=1.025
+ $X2=3.015 $Y2=1.217
r126 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.015 $Y=1.025
+ $X2=3.015 $Y2=0.56
r127 21 54 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.99 $Y=1.41
+ $X2=2.99 $Y2=1.217
r128 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.99 $Y=1.41
+ $X2=2.99 $Y2=1.985
r129 18 52 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.52 $Y=1.41
+ $X2=2.52 $Y2=1.217
r130 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.52 $Y=1.41
+ $X2=2.52 $Y2=1.985
r131 14 51 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.495 $Y=1.025
+ $X2=2.495 $Y2=1.217
r132 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.495 $Y=1.025
+ $X2=2.495 $Y2=0.56
r133 11 50 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.05 $Y=1.41
+ $X2=2.05 $Y2=1.217
r134 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.05 $Y=1.41
+ $X2=2.05 $Y2=1.985
r135 7 49 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.025 $Y=1.025
+ $X2=2.025 $Y2=1.217
r136 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.025 $Y=1.025
+ $X2=2.025 $Y2=0.56
r137 2 46 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.63
r138 2 30 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=2.31
r139 1 42 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.13
+ $Y=0.235 $X2=1.265 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_8%A_338_47# 1 2 3 4 15 17 19 22 24 26 29 31
+ 33 36 38 40 43 45 47 50 52 54 57 59 61 62 64 67 71 75 79 80 81 82 85 89 93 95
+ 98 100 106 109 110 111 128
c242 128 0 1.39726e-19 $X=6.75 $Y=1.217
r243 128 129 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=6.75 $Y=1.217
+ $X2=6.775 $Y2=1.217
r244 127 128 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=6.28 $Y=1.217
+ $X2=6.75 $Y2=1.217
r245 126 127 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=6.255 $Y=1.217
+ $X2=6.28 $Y2=1.217
r246 125 126 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=5.81 $Y=1.217
+ $X2=6.255 $Y2=1.217
r247 124 125 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=5.785 $Y=1.217
+ $X2=5.81 $Y2=1.217
r248 121 122 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=5.315 $Y=1.217
+ $X2=5.34 $Y2=1.217
r249 120 121 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=4.87 $Y=1.217
+ $X2=5.315 $Y2=1.217
r250 119 120 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.845 $Y=1.217
+ $X2=4.87 $Y2=1.217
r251 118 119 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=4.4 $Y=1.217
+ $X2=4.845 $Y2=1.217
r252 117 118 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.375 $Y=1.217
+ $X2=4.4 $Y2=1.217
r253 116 117 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=3.93 $Y=1.217
+ $X2=4.375 $Y2=1.217
r254 115 116 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.905 $Y=1.217
+ $X2=3.93 $Y2=1.217
r255 112 113 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.435 $Y=1.217
+ $X2=3.46 $Y2=1.217
r256 107 124 47.9006 $w=3.22e-07 $l=3.2e-07 $layer=POLY_cond $X=5.465 $Y=1.217
+ $X2=5.785 $Y2=1.217
r257 107 122 18.7112 $w=3.22e-07 $l=1.25e-07 $layer=POLY_cond $X=5.465 $Y=1.217
+ $X2=5.34 $Y2=1.217
r258 106 107 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=5.465
+ $Y=1.16 $X2=5.465 $Y2=1.16
r259 104 115 50.8944 $w=3.22e-07 $l=3.4e-07 $layer=POLY_cond $X=3.565 $Y=1.217
+ $X2=3.905 $Y2=1.217
r260 104 113 15.7174 $w=3.22e-07 $l=1.05e-07 $layer=POLY_cond $X=3.565 $Y=1.217
+ $X2=3.46 $Y2=1.217
r261 103 106 105.364 $w=1.98e-07 $l=1.9e-06 $layer=LI1_cond $X=3.565 $Y=1.175
+ $X2=5.465 $Y2=1.175
r262 103 104 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.565
+ $Y=1.16 $X2=3.565 $Y2=1.16
r263 101 111 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=1.175
+ $X2=3.225 $Y2=1.175
r264 101 103 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=3.31 $Y=1.175
+ $X2=3.565 $Y2=1.175
r265 99 111 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.225 $Y=1.275
+ $X2=3.225 $Y2=1.175
r266 99 100 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.225 $Y=1.275
+ $X2=3.225 $Y2=1.445
r267 98 111 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.225 $Y=1.075
+ $X2=3.225 $Y2=1.175
r268 97 98 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.225 $Y=0.905
+ $X2=3.225 $Y2=1.075
r269 96 110 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.92 $Y=1.53
+ $X2=2.73 $Y2=1.53
r270 95 100 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.14 $Y=1.53
+ $X2=3.225 $Y2=1.445
r271 95 96 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.14 $Y=1.53
+ $X2=2.92 $Y2=1.53
r272 94 109 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.92 $Y=0.82
+ $X2=2.73 $Y2=0.82
r273 93 97 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.14 $Y=0.82
+ $X2=3.225 $Y2=0.905
r274 93 94 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.14 $Y=0.82
+ $X2=2.92 $Y2=0.82
r275 89 91 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.73 $Y=1.63
+ $X2=2.73 $Y2=2.31
r276 87 110 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=1.615
+ $X2=2.73 $Y2=1.53
r277 87 89 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.73 $Y=1.615
+ $X2=2.73 $Y2=1.63
r278 83 109 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=0.735
+ $X2=2.73 $Y2=0.82
r279 83 85 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.73 $Y=0.735
+ $X2=2.73 $Y2=0.4
r280 81 110 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.54 $Y=1.53
+ $X2=2.73 $Y2=1.53
r281 81 82 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.54 $Y=1.53
+ $X2=1.98 $Y2=1.53
r282 79 109 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.54 $Y=0.82
+ $X2=2.73 $Y2=0.82
r283 79 80 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.54 $Y=0.82
+ $X2=1.98 $Y2=0.82
r284 75 77 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.815 $Y=1.63
+ $X2=1.815 $Y2=2.31
r285 73 82 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.815 $Y=1.615
+ $X2=1.98 $Y2=1.53
r286 73 75 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.815 $Y=1.615
+ $X2=1.815 $Y2=1.63
r287 69 80 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.815 $Y=0.735
+ $X2=1.98 $Y2=0.82
r288 69 71 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.815 $Y=0.735
+ $X2=1.815 $Y2=0.4
r289 65 129 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.775 $Y=1.025
+ $X2=6.775 $Y2=1.217
r290 65 67 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.775 $Y=1.025
+ $X2=6.775 $Y2=0.56
r291 62 128 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.75 $Y=1.41
+ $X2=6.75 $Y2=1.217
r292 62 64 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.75 $Y=1.41
+ $X2=6.75 $Y2=1.985
r293 59 127 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.28 $Y=1.41
+ $X2=6.28 $Y2=1.217
r294 59 61 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.28 $Y=1.41
+ $X2=6.28 $Y2=1.985
r295 55 126 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.255 $Y=1.025
+ $X2=6.255 $Y2=1.217
r296 55 57 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.255 $Y=1.025
+ $X2=6.255 $Y2=0.56
r297 52 125 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.81 $Y=1.41
+ $X2=5.81 $Y2=1.217
r298 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.81 $Y=1.41
+ $X2=5.81 $Y2=1.985
r299 48 124 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.785 $Y=1.025
+ $X2=5.785 $Y2=1.217
r300 48 50 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.785 $Y=1.025
+ $X2=5.785 $Y2=0.56
r301 45 122 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.34 $Y=1.41
+ $X2=5.34 $Y2=1.217
r302 45 47 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.34 $Y=1.41
+ $X2=5.34 $Y2=1.985
r303 41 121 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.315 $Y=1.025
+ $X2=5.315 $Y2=1.217
r304 41 43 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.315 $Y=1.025
+ $X2=5.315 $Y2=0.56
r305 38 120 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.87 $Y=1.41
+ $X2=4.87 $Y2=1.217
r306 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.87 $Y=1.41
+ $X2=4.87 $Y2=1.985
r307 34 119 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.845 $Y=1.025
+ $X2=4.845 $Y2=1.217
r308 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.845 $Y=1.025
+ $X2=4.845 $Y2=0.56
r309 31 118 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.4 $Y=1.41
+ $X2=4.4 $Y2=1.217
r310 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.4 $Y=1.41
+ $X2=4.4 $Y2=1.985
r311 27 117 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.375 $Y=1.025
+ $X2=4.375 $Y2=1.217
r312 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.375 $Y=1.025
+ $X2=4.375 $Y2=0.56
r313 24 116 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.93 $Y=1.41
+ $X2=3.93 $Y2=1.217
r314 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.93 $Y=1.41
+ $X2=3.93 $Y2=1.985
r315 20 115 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.905 $Y=1.025
+ $X2=3.905 $Y2=1.217
r316 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.905 $Y=1.025
+ $X2=3.905 $Y2=0.56
r317 17 113 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.46 $Y=1.41
+ $X2=3.46 $Y2=1.217
r318 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.46 $Y=1.41
+ $X2=3.46 $Y2=1.985
r319 13 112 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.435 $Y=1.025
+ $X2=3.435 $Y2=1.217
r320 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.435 $Y=1.025
+ $X2=3.435 $Y2=0.56
r321 4 91 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=1.485 $X2=2.755 $Y2=2.31
r322 4 89 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=1.485 $X2=2.755 $Y2=1.63
r323 3 77 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.69
+ $Y=1.485 $X2=1.815 $Y2=2.31
r324 3 75 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.69
+ $Y=1.485 $X2=1.815 $Y2=1.63
r325 2 85 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.235 $X2=2.755 $Y2=0.4
r326 1 71 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.69
+ $Y=0.235 $X2=1.815 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_8%VPWR 1 2 3 4 5 6 7 26 30 34 38 42 46 50
+ 53 54 56 57 59 60 62 63 65 66 68 69 70 95 96 99
c113 1 0 1.38193e-19 $X=0.585 $Y=1.485
r114 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r116 93 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r117 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r118 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r119 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r120 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r121 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r122 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r123 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r124 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r125 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r126 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r127 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r128 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r129 75 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r130 74 77 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r131 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r132 72 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.73 $Y2=2.72
r133 72 74 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=1.15 $Y2=2.72
r134 70 100 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r135 68 92 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.9 $Y=2.72
+ $X2=6.67 $Y2=2.72
r136 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.9 $Y=2.72
+ $X2=6.985 $Y2=2.72
r137 67 95 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=7.07 $Y=2.72 $X2=7.13
+ $Y2=2.72
r138 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.07 $Y=2.72
+ $X2=6.985 $Y2=2.72
r139 65 89 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.96 $Y=2.72
+ $X2=5.75 $Y2=2.72
r140 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=2.72
+ $X2=6.045 $Y2=2.72
r141 64 92 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=6.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r142 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=2.72
+ $X2=6.045 $Y2=2.72
r143 62 86 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.02 $Y=2.72
+ $X2=4.83 $Y2=2.72
r144 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.02 $Y=2.72
+ $X2=5.105 $Y2=2.72
r145 61 89 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.19 $Y=2.72
+ $X2=5.75 $Y2=2.72
r146 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=2.72
+ $X2=5.105 $Y2=2.72
r147 59 83 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.08 $Y=2.72
+ $X2=3.91 $Y2=2.72
r148 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=2.72
+ $X2=4.165 $Y2=2.72
r149 58 86 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.25 $Y=2.72
+ $X2=4.83 $Y2=2.72
r150 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.25 $Y=2.72
+ $X2=4.165 $Y2=2.72
r151 56 80 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.14 $Y=2.72
+ $X2=2.99 $Y2=2.72
r152 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=2.72
+ $X2=3.225 $Y2=2.72
r153 55 83 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.31 $Y=2.72 $X2=3.91
+ $Y2=2.72
r154 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=2.72
+ $X2=3.225 $Y2=2.72
r155 53 77 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.2 $Y=2.72
+ $X2=2.07 $Y2=2.72
r156 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.72
+ $X2=2.285 $Y2=2.72
r157 52 80 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.37 $Y=2.72
+ $X2=2.99 $Y2=2.72
r158 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=2.72
+ $X2=2.285 $Y2=2.72
r159 48 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=2.635
+ $X2=6.985 $Y2=2.72
r160 48 50 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.985 $Y=2.635
+ $X2=6.985 $Y2=2
r161 44 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=2.635
+ $X2=6.045 $Y2=2.72
r162 44 46 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.045 $Y=2.635
+ $X2=6.045 $Y2=2
r163 40 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=2.635
+ $X2=5.105 $Y2=2.72
r164 40 42 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.105 $Y=2.635
+ $X2=5.105 $Y2=2
r165 36 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=2.635
+ $X2=4.165 $Y2=2.72
r166 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.165 $Y=2.635
+ $X2=4.165 $Y2=2
r167 32 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=2.635
+ $X2=3.225 $Y2=2.72
r168 32 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.225 $Y=2.635
+ $X2=3.225 $Y2=2
r169 28 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.285 $Y=2.635
+ $X2=2.285 $Y2=2.72
r170 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.285 $Y=2.635
+ $X2=2.285 $Y2=2
r171 24 99 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r172 24 26 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=1.95
r173 7 50 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.84
+ $Y=1.485 $X2=6.985 $Y2=2
r174 6 46 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.9
+ $Y=1.485 $X2=6.045 $Y2=2
r175 5 42 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.96
+ $Y=1.485 $X2=5.105 $Y2=2
r176 4 38 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.02
+ $Y=1.485 $X2=4.165 $Y2=2
r177 3 34 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.08
+ $Y=1.485 $X2=3.225 $Y2=2
r178 2 30 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.14
+ $Y=1.485 $X2=2.285 $Y2=2
r179 1 26 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_8%X 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45
+ 49 51 55 59 63 65 69 73 77 79 81 82 83 84 85 86 88 89
c171 79 0 1.95897e-19 $X=6.86 $Y=1.53
c172 38 0 1.26528e-19 $X=3.86 $Y=1.53
c173 36 0 1.25206e-19 $X=3.86 $Y=0.82
r174 88 89 6.69888 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=7.05 $Y=1.19
+ $X2=7.05 $Y2=1.445
r175 87 88 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=7.05 $Y=0.905
+ $X2=7.05 $Y2=1.19
r176 80 86 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.68 $Y=1.53
+ $X2=6.49 $Y2=1.53
r177 79 89 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.86 $Y=1.53
+ $X2=7.05 $Y2=1.53
r178 79 80 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.86 $Y=1.53
+ $X2=6.68 $Y2=1.53
r179 78 85 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.68 $Y=0.82
+ $X2=6.49 $Y2=0.82
r180 77 87 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=6.86 $Y=0.82
+ $X2=7.05 $Y2=0.905
r181 77 78 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.86 $Y=0.82
+ $X2=6.68 $Y2=0.82
r182 73 75 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.49 $Y=1.63
+ $X2=6.49 $Y2=2.31
r183 71 86 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=1.615
+ $X2=6.49 $Y2=1.53
r184 71 73 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=6.49 $Y=1.615
+ $X2=6.49 $Y2=1.63
r185 67 85 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=0.735
+ $X2=6.49 $Y2=0.82
r186 67 69 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.49 $Y=0.735
+ $X2=6.49 $Y2=0.4
r187 66 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.74 $Y=1.53
+ $X2=5.55 $Y2=1.53
r188 65 86 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.3 $Y=1.53 $X2=6.49
+ $Y2=1.53
r189 65 66 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.3 $Y=1.53
+ $X2=5.74 $Y2=1.53
r190 64 83 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.74 $Y=0.82
+ $X2=5.55 $Y2=0.82
r191 63 85 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.3 $Y=0.82 $X2=6.49
+ $Y2=0.82
r192 63 64 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.3 $Y=0.82
+ $X2=5.74 $Y2=0.82
r193 59 61 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=5.55 $Y=1.63
+ $X2=5.55 $Y2=2.31
r194 57 84 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=1.615
+ $X2=5.55 $Y2=1.53
r195 57 59 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=5.55 $Y=1.615
+ $X2=5.55 $Y2=1.63
r196 53 83 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=0.735
+ $X2=5.55 $Y2=0.82
r197 53 55 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.55 $Y=0.735
+ $X2=5.55 $Y2=0.4
r198 52 82 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.8 $Y=1.53 $X2=4.61
+ $Y2=1.53
r199 51 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.36 $Y=1.53
+ $X2=5.55 $Y2=1.53
r200 51 52 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.36 $Y=1.53
+ $X2=4.8 $Y2=1.53
r201 50 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.8 $Y=0.82 $X2=4.61
+ $Y2=0.82
r202 49 83 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.36 $Y=0.82
+ $X2=5.55 $Y2=0.82
r203 49 50 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.36 $Y=0.82
+ $X2=4.8 $Y2=0.82
r204 45 47 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=4.61 $Y=1.63
+ $X2=4.61 $Y2=2.31
r205 43 82 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=1.615
+ $X2=4.61 $Y2=1.53
r206 43 45 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=4.61 $Y=1.615
+ $X2=4.61 $Y2=1.63
r207 39 81 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=0.735
+ $X2=4.61 $Y2=0.82
r208 39 41 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.61 $Y=0.735
+ $X2=4.61 $Y2=0.4
r209 37 82 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.42 $Y=1.53
+ $X2=4.61 $Y2=1.53
r210 37 38 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.42 $Y=1.53
+ $X2=3.86 $Y2=1.53
r211 35 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.42 $Y=0.82
+ $X2=4.61 $Y2=0.82
r212 35 36 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.42 $Y=0.82
+ $X2=3.86 $Y2=0.82
r213 31 33 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.67 $Y=1.63
+ $X2=3.67 $Y2=2.31
r214 29 38 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.67 $Y=1.615
+ $X2=3.86 $Y2=1.53
r215 29 31 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.67 $Y=1.615
+ $X2=3.67 $Y2=1.63
r216 25 36 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.67 $Y=0.735
+ $X2=3.86 $Y2=0.82
r217 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.67 $Y=0.735
+ $X2=3.67 $Y2=0.4
r218 8 75 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.37
+ $Y=1.485 $X2=6.515 $Y2=2.31
r219 8 73 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.37
+ $Y=1.485 $X2=6.515 $Y2=1.63
r220 7 61 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=1.485 $X2=5.575 $Y2=2.31
r221 7 59 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=1.485 $X2=5.575 $Y2=1.63
r222 6 47 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=4.49
+ $Y=1.485 $X2=4.635 $Y2=2.31
r223 6 45 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.49
+ $Y=1.485 $X2=4.635 $Y2=1.63
r224 5 33 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.55
+ $Y=1.485 $X2=3.695 $Y2=2.31
r225 5 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.55
+ $Y=1.485 $X2=3.695 $Y2=1.63
r226 4 69 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=6.33
+ $Y=0.235 $X2=6.515 $Y2=0.4
r227 3 55 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=5.39
+ $Y=0.235 $X2=5.575 $Y2=0.4
r228 2 41 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=4.45
+ $Y=0.235 $X2=4.635 $Y2=0.4
r229 1 27 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=3.51
+ $Y=0.235 $X2=3.695 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUFBUF_8%VGND 1 2 3 4 5 6 7 26 30 34 38 42 46 50
+ 53 54 56 57 59 60 62 63 65 66 68 69 70 95 96 99 102
r126 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r127 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r128 93 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r129 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r130 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r131 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r132 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r133 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r134 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r135 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r136 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r137 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r138 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r139 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r140 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r141 75 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r142 74 77 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r143 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r144 72 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r145 72 74 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0
+ $X2=1.15 $Y2=0
r146 70 100 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r147 70 102 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r148 68 92 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.9 $Y=0 $X2=6.67
+ $Y2=0
r149 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.9 $Y=0 $X2=6.985
+ $Y2=0
r150 67 95 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=7.07 $Y=0 $X2=7.13
+ $Y2=0
r151 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.07 $Y=0 $X2=6.985
+ $Y2=0
r152 65 89 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.96 $Y=0 $X2=5.75
+ $Y2=0
r153 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=0 $X2=6.045
+ $Y2=0
r154 64 92 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6.67
+ $Y2=0
r155 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=0 $X2=6.045
+ $Y2=0
r156 62 86 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.02 $Y=0 $X2=4.83
+ $Y2=0
r157 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.02 $Y=0 $X2=5.105
+ $Y2=0
r158 61 89 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.19 $Y=0 $X2=5.75
+ $Y2=0
r159 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=0 $X2=5.105
+ $Y2=0
r160 59 83 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=3.91
+ $Y2=0
r161 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=0 $X2=4.165
+ $Y2=0
r162 58 86 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.25 $Y=0 $X2=4.83
+ $Y2=0
r163 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.25 $Y=0 $X2=4.165
+ $Y2=0
r164 56 80 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=2.99
+ $Y2=0
r165 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.225
+ $Y2=0
r166 55 83 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.31 $Y=0 $X2=3.91
+ $Y2=0
r167 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=0 $X2=3.225
+ $Y2=0
r168 53 77 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.2 $Y=0 $X2=2.07
+ $Y2=0
r169 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0 $X2=2.285
+ $Y2=0
r170 52 80 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.99
+ $Y2=0
r171 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.285
+ $Y2=0
r172 48 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=0.085
+ $X2=6.985 $Y2=0
r173 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.985 $Y=0.085
+ $X2=6.985 $Y2=0.4
r174 44 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=0.085
+ $X2=6.045 $Y2=0
r175 44 46 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.045 $Y=0.085
+ $X2=6.045 $Y2=0.4
r176 40 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=0.085
+ $X2=5.105 $Y2=0
r177 40 42 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.105 $Y=0.085
+ $X2=5.105 $Y2=0.4
r178 36 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=0.085
+ $X2=4.165 $Y2=0
r179 36 38 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.165 $Y=0.085
+ $X2=4.165 $Y2=0.4
r180 32 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=0.085
+ $X2=3.225 $Y2=0
r181 32 34 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.225 $Y=0.085
+ $X2=3.225 $Y2=0.4
r182 28 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.285 $Y=0.085
+ $X2=2.285 $Y2=0
r183 28 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.285 $Y=0.085
+ $X2=2.285 $Y2=0.4
r184 24 99 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r185 24 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.4
r186 7 50 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.85
+ $Y=0.235 $X2=6.985 $Y2=0.4
r187 6 46 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=5.86
+ $Y=0.235 $X2=6.045 $Y2=0.4
r188 5 42 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.92
+ $Y=0.235 $X2=5.105 $Y2=0.4
r189 4 38 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.98
+ $Y=0.235 $X2=4.165 $Y2=0.4
r190 3 34 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.09
+ $Y=0.235 $X2=3.225 $Y2=0.4
r191 2 30 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.1
+ $Y=0.235 $X2=2.285 $Y2=0.4
r192 1 26 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

