# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__ebufn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__ebufn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 0.765000 0.830000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.954300 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.765000 1.380000 1.425000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.445000 6.335000 1.725000 ;
        RECT 4.495000 0.615000 6.335000 0.855000 ;
        RECT 6.105000 0.855000 6.335000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.440000 0.085000 ;
        RECT 0.515000  0.085000 0.980000 0.595000 ;
        RECT 2.495000  0.085000 2.875000 0.485000 ;
        RECT 3.435000  0.085000 3.815000 0.485000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.440000 2.805000 ;
        RECT 0.515000 1.845000 0.980000 2.635000 ;
        RECT 2.080000 2.275000 2.460000 2.635000 ;
        RECT 3.070000 2.275000 3.400000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.280000 0.345000 0.665000 ;
      RECT 0.085000 0.665000 0.320000 1.765000 ;
      RECT 0.085000 1.765000 0.345000 2.465000 ;
      RECT 1.200000 0.255000 1.825000 0.595000 ;
      RECT 1.200000 1.595000 1.825000 1.765000 ;
      RECT 1.200000 1.765000 1.455000 2.465000 ;
      RECT 1.550000 0.595000 1.825000 1.025000 ;
      RECT 1.550000 1.025000 4.160000 1.275000 ;
      RECT 1.550000 1.275000 1.825000 1.595000 ;
      RECT 1.665000 1.935000 6.285000 2.105000 ;
      RECT 1.665000 2.105000 1.910000 2.465000 ;
      RECT 1.995000 0.255000 2.325000 0.655000 ;
      RECT 1.995000 0.655000 4.325000 0.855000 ;
      RECT 1.995000 1.895000 6.285000 1.935000 ;
      RECT 2.680000 2.105000 2.850000 2.465000 ;
      RECT 3.095000 0.275000 3.265000 0.655000 ;
      RECT 3.620000 2.105000 6.285000 2.465000 ;
      RECT 4.035000 0.255000 6.285000 0.445000 ;
      RECT 4.035000 0.445000 4.325000 0.655000 ;
      RECT 4.330000 1.025000 5.935000 1.275000 ;
    LAYER mcon ;
      RECT 0.150000 1.105000 0.320000 1.275000 ;
      RECT 4.710000 1.105000 4.880000 1.275000 ;
    LAYER met1 ;
      RECT 0.085000 1.075000 0.380000 1.165000 ;
      RECT 0.085000 1.165000 4.940000 1.305000 ;
      RECT 4.650000 1.075000 4.940000 1.165000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_4
