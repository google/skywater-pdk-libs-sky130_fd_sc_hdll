* File: sky130_fd_sc_hdll__a2bb2oi_1.pex.spice
* Created: Wed Sep  2 08:19:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A1_N 1 3 4 6 7 8 13
r24 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r25 7 8 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.335 $Y=1.19 $X2=0.335
+ $Y2=1.53
r26 7 13 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=0.335 $Y=1.19
+ $X2=0.335 $Y2=1.16
r27 4 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.435 $Y2=1.16
r28 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r29 1 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.435 $Y2=1.16
r30 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A2_N 1 3 4 6 7 15
r30 11 15 9.13257 $w=2.63e-07 $l=2.1e-07 $layer=LI1_cond $X=0.94 $Y=1.142
+ $X2=1.15 $Y2=1.142
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r32 7 15 4.56628 $w=2.63e-07 $l=1.05e-07 $layer=LI1_cond $X=1.255 $Y=1.142
+ $X2=1.15 $Y2=1.142
r33 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1 $Y=0.995
+ $X2=0.94 $Y2=1.16
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1 $Y=0.995 $X2=1
+ $Y2=0.56
r35 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.94 $Y2=1.16
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A_119_47# 1 2 7 9 10 12 13 16 17 20 24
+ 25 29
r66 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.16 $X2=1.73 $Y2=1.16
r67 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.73 $Y=1.445
+ $X2=1.73 $Y2=1.16
r68 26 29 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.73 $Y=0.83
+ $X2=1.73 $Y2=1.16
r69 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.645 $Y=1.53
+ $X2=1.73 $Y2=1.445
r70 24 25 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.645 $Y=1.53
+ $X2=1.305 $Y2=1.53
r71 20 22 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.115 $Y=1.64
+ $X2=1.115 $Y2=2.32
r72 18 25 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=1.115 $Y=1.615
+ $X2=1.305 $Y2=1.53
r73 18 20 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=1.115 $Y=1.615
+ $X2=1.115 $Y2=1.64
r74 16 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.645 $Y=0.745
+ $X2=1.73 $Y2=0.83
r75 16 17 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.645 $Y=0.745
+ $X2=0.815 $Y2=0.745
r76 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.73 $Y=0.66
+ $X2=0.815 $Y2=0.745
r77 13 15 7.17647 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.73 $Y=0.66 $X2=0.73
+ $Y2=0.56
r78 10 30 39.7049 $w=4.06e-07 $l=2.29783e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.825 $Y2=1.16
r79 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.98 $Y2=0.56
r80 7 30 44.8379 $w=4.06e-07 $l=3.08221e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.825 $Y2=1.16
r81 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r82 2 22 400 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.485 $X2=1.14 $Y2=2.32
r83 2 20 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.485 $X2=1.14 $Y2=1.64
r84 1 15 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_1%B2 1 3 4 6 7 8 9 10 27
r40 25 27 2.50531 $w=2.28e-07 $l=5e-08 $layer=LI1_cond $X=2.5 $Y=1.11 $X2=2.5
+ $Y2=1.16
r41 17 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.16 $X2=2.47 $Y2=1.16
r42 9 25 0.150319 $w=2.28e-07 $l=3e-09 $layer=LI1_cond $X=2.5 $Y=1.107 $X2=2.5
+ $Y2=1.11
r43 9 33 6.41961 $w=2.28e-07 $l=1.12e-07 $layer=LI1_cond $X=2.5 $Y=1.107 $X2=2.5
+ $Y2=0.995
r44 9 10 16.9359 $w=2.28e-07 $l=3.38e-07 $layer=LI1_cond $X=2.5 $Y=1.192 $X2=2.5
+ $Y2=1.53
r45 9 27 1.6034 $w=2.28e-07 $l=3.2e-08 $layer=LI1_cond $X=2.5 $Y=1.192 $X2=2.5
+ $Y2=1.16
r46 8 33 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.53 $Y=0.85
+ $X2=2.53 $Y2=0.995
r47 7 8 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.53 $Y=0.51 $X2=2.53
+ $Y2=0.85
r48 4 17 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.53 $Y=0.995
+ $X2=2.47 $Y2=1.16
r49 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.53 $Y=0.995 $X2=2.53
+ $Y2=0.56
r50 1 17 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.47 $Y2=1.16
r51 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.505 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_1%B1 1 3 4 6 7 14
c26 4 0 8.41034e-20 $X=2.985 $Y=1.41
r27 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.02
+ $Y=1.16 $X2=3.02 $Y2=1.16
r28 7 14 1.06104 $w=6.18e-07 $l=5.5e-08 $layer=LI1_cond $X=3.075 $Y=1.305
+ $X2=3.02 $Y2=1.305
r29 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=3.02 $Y2=1.16
r30 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=2.985 $Y2=1.985
r31 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.96 $Y=0.995
+ $X2=3.02 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.96 $Y=0.995 $X2=2.96
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_1%VPWR 1 2 9 12 13 14 17 27 28 36
r45 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 25 28 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 22 25 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 21 24 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 19 21 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 17 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 14 36 16.8131 $w=4.98e-07 $l=6.45e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=1.99
r54 14 19 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.212 $Y=2.72
+ $X2=0.425 $Y2=2.72
r55 14 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 12 24 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.665 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 12 13 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.665 $Y=2.72
+ $X2=2.79 $Y2=2.72
r58 11 27 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 11 13 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=2.79 $Y2=2.72
r60 7 13 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=2.635
+ $X2=2.79 $Y2=2.72
r61 7 9 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.79 $Y=2.635
+ $X2=2.79 $Y2=2.36
r62 2 9 600 $w=1.7e-07 $l=9.49342e-07 $layer=licon1_PDIFF $count=1 $X=2.595
+ $Y=1.485 $X2=2.75 $Y2=2.36
r63 1 36 300 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_1%Y 1 2 8 10 11 12 13 20 32 37
r37 12 20 7.26197 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=1.702 $Y=2.21
+ $X2=1.702 $Y2=1.98
r38 11 37 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=1.87
+ $X2=2.07 $Y2=1.87
r39 11 32 6.32834 $w=1.68e-07 $l=9.7e-08 $layer=LI1_cond $X=1.702 $Y=1.87
+ $X2=1.605 $Y2=1.87
r40 11 20 1.77461 $w=5.33e-07 $l=2.5e-08 $layer=LI1_cond $X=1.702 $Y=1.955
+ $X2=1.702 $Y2=1.98
r41 9 13 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.13 $Y=0.68 $X2=2.13
+ $Y2=0.51
r42 9 10 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.13 $Y=0.68
+ $X2=2.13 $Y2=0.825
r43 8 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=1.785
+ $X2=2.07 $Y2=1.87
r44 8 10 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.07 $Y=1.785 $X2=2.07
+ $Y2=0.825
r45 2 20 300 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.485 $X2=1.72 $Y2=1.98
r46 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A_409_297# 1 2 8 9 10 11 13 18
c33 11 0 8.41034e-20 $X=3.262 $Y=1.955
r34 16 18 7.01487 $w=2.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.27 $Y=2.35
+ $X2=2.41 $Y2=2.35
r35 11 21 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.262 $Y=1.955
+ $X2=3.262 $Y2=1.87
r36 11 13 15.5919 $w=2.53e-07 $l=3.45e-07 $layer=LI1_cond $X=3.262 $Y=1.955
+ $X2=3.262 $Y2=2.3
r37 9 21 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.135 $Y=1.87
+ $X2=3.262 $Y2=1.87
r38 9 10 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.135 $Y=1.87
+ $X2=2.495 $Y2=1.87
r39 8 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.41 $Y=2.235
+ $X2=2.41 $Y2=2.35
r40 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.41 $Y=1.955
+ $X2=2.495 $Y2=1.87
r41 7 8 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.41 $Y=1.955 $X2=2.41
+ $Y2=2.235
r42 2 21 600 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=1.485 $X2=3.22 $Y2=1.87
r43 2 13 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=1.485 $X2=3.22 $Y2=2.3
r44 1 16 600 $w=1.7e-07 $l=9.40798e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.27 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_1%VGND 1 2 3 12 15 16 17 20 35 36 46 52 54
r47 50 52 8.74535 $w=5.73e-07 $l=1.05e-07 $layer=LI1_cond $X=1.61 $Y=0.202
+ $X2=1.715 $Y2=0.202
r48 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r49 48 50 1.24808 $w=5.73e-07 $l=6e-08 $layer=LI1_cond $X=1.55 $Y=0.202 $X2=1.61
+ $Y2=0.202
r50 45 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r51 44 48 8.32055 $w=5.73e-07 $l=4e-07 $layer=LI1_cond $X=1.15 $Y=0.202 $X2=1.55
+ $Y2=0.202
r52 44 46 8.74535 $w=5.73e-07 $l=1.05e-07 $layer=LI1_cond $X=1.15 $Y=0.202
+ $X2=1.045 $Y2=0.202
r53 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r55 33 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r56 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r57 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r58 30 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r59 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r60 29 52 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.715
+ $Y2=0
r61 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r62 26 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r63 25 46 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.045
+ $Y2=0
r64 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r65 23 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r66 20 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r67 17 54 8.44056 $w=4.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r68 17 23 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.212 $Y=0 $X2=0.425
+ $Y2=0
r69 17 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r70 15 32 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.005 $Y=0 $X2=2.99
+ $Y2=0
r71 15 16 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.005 $Y=0 $X2=3.195
+ $Y2=0
r72 14 35 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.45
+ $Y2=0
r73 14 16 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.195
+ $Y2=0
r74 10 16 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=0.085
+ $X2=3.195 $Y2=0
r75 10 12 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.195 $Y=0.085
+ $X2=3.195 $Y2=0.38
r76 3 12 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.035
+ $Y=0.235 $X2=3.22 $Y2=0.38
r77 2 48 91 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.235 $X2=1.55 $Y2=0.38
r78 1 54 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

