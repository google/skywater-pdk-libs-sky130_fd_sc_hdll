* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__clkinvlp_4 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.4e+11p pd=5.08e+06u as=7.9e+11p ps=7.58e+06u
M1001 Y A a_110_47# VNB nshort w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=1.155e+11p ps=1.52e+06u
M1002 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_110_47# A VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=2.8875e+11p ps=3.25e+06u
M1004 VGND A a_268_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.52e+06u
M1005 a_268_47# A Y VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends
