* File: sky130_fd_sc_hdll__o21bai_1.pxi.spice
* Created: Thu Aug 27 19:19:56 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21BAI_1%B1_N N_B1_N_c_56_n N_B1_N_M1002_g N_B1_N_c_57_n
+ N_B1_N_c_58_n N_B1_N_M1006_g N_B1_N_c_53_n N_B1_N_c_54_n B1_N N_B1_N_c_55_n
+ PM_SKY130_FD_SC_HDLL__O21BAI_1%B1_N
x_PM_SKY130_FD_SC_HDLL__O21BAI_1%A_105_352# N_A_105_352#_M1002_d
+ N_A_105_352#_M1006_s N_A_105_352#_c_101_n N_A_105_352#_M1007_g
+ N_A_105_352#_c_94_n N_A_105_352#_M1004_g N_A_105_352#_c_95_n
+ N_A_105_352#_c_96_n N_A_105_352#_c_104_n N_A_105_352#_c_97_n
+ N_A_105_352#_c_105_n N_A_105_352#_c_98_n N_A_105_352#_c_99_n
+ N_A_105_352#_c_100_n PM_SKY130_FD_SC_HDLL__O21BAI_1%A_105_352#
x_PM_SKY130_FD_SC_HDLL__O21BAI_1%A2 N_A2_c_153_n N_A2_M1001_g N_A2_c_154_n
+ N_A2_M1003_g A2 A2 PM_SKY130_FD_SC_HDLL__O21BAI_1%A2
x_PM_SKY130_FD_SC_HDLL__O21BAI_1%A1 N_A1_c_183_n N_A1_M1000_g N_A1_c_184_n
+ N_A1_M1005_g A1 A1 PM_SKY130_FD_SC_HDLL__O21BAI_1%A1
x_PM_SKY130_FD_SC_HDLL__O21BAI_1%VPWR N_VPWR_M1006_d N_VPWR_M1000_d
+ N_VPWR_c_205_n N_VPWR_c_206_n N_VPWR_c_207_n VPWR N_VPWR_c_208_n
+ N_VPWR_c_209_n N_VPWR_c_210_n N_VPWR_c_204_n
+ PM_SKY130_FD_SC_HDLL__O21BAI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O21BAI_1%Y N_Y_M1004_s N_Y_M1007_d N_Y_c_237_n
+ N_Y_c_239_n Y PM_SKY130_FD_SC_HDLL__O21BAI_1%Y
x_PM_SKY130_FD_SC_HDLL__O21BAI_1%VGND N_VGND_M1002_s N_VGND_M1003_d
+ N_VGND_c_270_n N_VGND_c_271_n N_VGND_c_272_n N_VGND_c_273_n N_VGND_c_274_n
+ VGND N_VGND_c_275_n N_VGND_c_276_n PM_SKY130_FD_SC_HDLL__O21BAI_1%VGND
x_PM_SKY130_FD_SC_HDLL__O21BAI_1%A_327_47# N_A_327_47#_M1004_d
+ N_A_327_47#_M1005_d N_A_327_47#_c_325_n N_A_327_47#_c_307_n
+ N_A_327_47#_c_308_n N_A_327_47#_c_309_n
+ PM_SKY130_FD_SC_HDLL__O21BAI_1%A_327_47#
cc_1 VNB N_B1_N_c_53_n 0.0146653f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_2 VNB N_B1_N_c_54_n 0.032184f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_3 VNB N_B1_N_c_55_n 0.0411574f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_4 VNB N_A_105_352#_c_94_n 0.0201038f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.97
cc_5 VNB N_A_105_352#_c_95_n 0.0431759f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.17
cc_6 VNB N_A_105_352#_c_96_n 0.0142923f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.345
cc_7 VNB N_A_105_352#_c_97_n 0.00587684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_105_352#_c_98_n 0.00107229f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.325
cc_9 VNB N_A_105_352#_c_99_n 0.00383545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_105_352#_c_100_n 0.00251215f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_153_n 0.0206979f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.325
cc_12 VNB N_A2_c_154_n 0.0174787f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.675
cc_13 VNB A2 0.00805763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_183_n 0.0273545f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.325
cc_15 VNB N_A1_c_184_n 0.0222311f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.675
cc_16 VNB A1 0.0169962f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.61
cc_17 VNB N_VPWR_c_204_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_237_n 0.00195089f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_270_n 0.0102019f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.61
cc_20 VNB N_VGND_c_271_n 0.032448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_272_n 0.00469858f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.17
cc_22 VNB N_VGND_c_273_n 0.0508202f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.17
cc_23 VNB N_VGND_c_274_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_24 VNB N_VGND_c_275_n 0.0252698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_276_n 0.207843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_327_47#_c_307_n 0.017008f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.97
cc_27 VNB N_A_327_47#_c_308_n 0.0031057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_327_47#_c_309_n 0.0185545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_B1_N_c_56_n 0.0137644f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.535
cc_30 VPB N_B1_N_c_57_n 0.0254806f $X=-0.19 $Y=1.305 $X2=0.845 $Y2=1.61
cc_31 VPB N_B1_N_c_58_n 0.0149581f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.61
cc_32 VPB N_B1_N_M1006_g 0.0446907f $X=-0.19 $Y=1.305 $X2=0.935 $Y2=1.97
cc_33 VPB N_B1_N_c_53_n 0.00538841f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_34 VPB N_B1_N_c_54_n 0.00501256f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_35 VPB B1_N 0.0614815f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_36 VPB N_A_105_352#_c_101_n 0.0177465f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.61
cc_37 VPB N_A_105_352#_c_95_n 0.0154557f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.17
cc_38 VPB N_A_105_352#_c_96_n 0.00725888f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.345
cc_39 VPB N_A_105_352#_c_104_n 0.00503075f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_40 VPB N_A_105_352#_c_105_n 0.00376695f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.16
cc_41 VPB N_A_105_352#_c_98_n 0.00331143f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_42 VPB N_A2_c_153_n 0.0248855f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.325
cc_43 VPB N_A1_c_183_n 0.0318092f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.325
cc_44 VPB N_VPWR_c_205_n 0.00896885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_206_n 0.0168816f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.17
cc_46 VPB N_VPWR_c_207_n 0.0541346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_208_n 0.0319134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_209_n 0.0278912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_210_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_204_n 0.0592181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_Y_c_237_n 0.00150073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_Y_c_239_n 0.00438941f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.17
cc_53 N_B1_N_c_57_n N_A_105_352#_c_101_n 0.0039572f $X=0.845 $Y=1.61 $X2=0 $Y2=0
cc_54 N_B1_N_M1006_g N_A_105_352#_c_101_n 0.0213546f $X=0.935 $Y=1.97 $X2=0
+ $Y2=0
cc_55 N_B1_N_c_57_n N_A_105_352#_c_95_n 0.0123728f $X=0.845 $Y=1.61 $X2=0 $Y2=0
cc_56 N_B1_N_c_53_n N_A_105_352#_c_95_n 3.11035e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_57 N_B1_N_c_54_n N_A_105_352#_c_95_n 0.0205724f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_58 N_B1_N_c_58_n N_A_105_352#_c_104_n 0.00445625f $X=0.635 $Y=1.61 $X2=0
+ $Y2=0
cc_59 N_B1_N_M1006_g N_A_105_352#_c_104_n 0.0093092f $X=0.935 $Y=1.97 $X2=0
+ $Y2=0
cc_60 B1_N N_A_105_352#_c_104_n 0.0407329f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_61 N_B1_N_c_53_n N_A_105_352#_c_97_n 0.0219349f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_62 N_B1_N_c_54_n N_A_105_352#_c_97_n 0.00428175f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_63 N_B1_N_c_57_n N_A_105_352#_c_105_n 0.0159307f $X=0.845 $Y=1.61 $X2=0 $Y2=0
cc_64 N_B1_N_c_58_n N_A_105_352#_c_105_n 0.0087797f $X=0.635 $Y=1.61 $X2=0 $Y2=0
cc_65 N_B1_N_M1006_g N_A_105_352#_c_105_n 0.00858486f $X=0.935 $Y=1.97 $X2=0
+ $Y2=0
cc_66 N_B1_N_c_53_n N_A_105_352#_c_105_n 6.56352e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_67 B1_N N_A_105_352#_c_105_n 0.0137262f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_68 N_B1_N_c_56_n N_A_105_352#_c_98_n 0.00428175f $X=0.535 $Y=1.535 $X2=0
+ $Y2=0
cc_69 N_B1_N_c_57_n N_A_105_352#_c_98_n 0.00247496f $X=0.845 $Y=1.61 $X2=0 $Y2=0
cc_70 B1_N N_A_105_352#_c_98_n 0.00829424f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_71 N_B1_N_c_55_n N_A_105_352#_c_100_n 0.00428175f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_72 N_B1_N_M1006_g N_VPWR_c_205_n 0.013544f $X=0.935 $Y=1.97 $X2=0 $Y2=0
cc_73 N_B1_N_M1006_g N_VPWR_c_208_n 0.00759451f $X=0.935 $Y=1.97 $X2=0 $Y2=0
cc_74 B1_N N_VPWR_c_208_n 0.0170586f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_75 N_B1_N_M1006_g N_VPWR_c_204_n 0.0148511f $X=0.935 $Y=1.97 $X2=0 $Y2=0
cc_76 B1_N N_VPWR_c_204_n 0.010222f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_77 N_B1_N_c_55_n N_Y_c_237_n 0.00599004f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B1_N_c_57_n N_Y_c_239_n 3.54712e-19 $X=0.845 $Y=1.61 $X2=0 $Y2=0
cc_79 N_B1_N_c_53_n N_VGND_c_271_n 0.0236731f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B1_N_c_54_n N_VGND_c_271_n 0.00102501f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B1_N_c_55_n N_VGND_c_271_n 0.0211895f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_82 N_B1_N_c_55_n N_VGND_c_273_n 0.00585385f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_83 N_B1_N_c_55_n N_VGND_c_276_n 0.0132583f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A_105_352#_c_101_n N_A2_c_153_n 0.0086027f $X=1.535 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_105_352#_c_96_n N_A2_c_153_n 0.0246834f $X=1.535 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_105_352#_c_94_n N_A2_c_154_n 0.00895029f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_105_352#_c_96_n A2 0.00194037f $X=1.535 $Y=1.202 $X2=0 $Y2=0
cc_88 N_A_105_352#_c_101_n N_VPWR_c_205_n 0.00695832f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_89 N_A_105_352#_c_95_n N_VPWR_c_205_n 0.00473925f $X=1.435 $Y=1.16 $X2=0
+ $Y2=0
cc_90 N_A_105_352#_c_104_n N_VPWR_c_205_n 0.0112115f $X=0.7 $Y=1.96 $X2=0 $Y2=0
cc_91 N_A_105_352#_c_104_n N_VPWR_c_208_n 0.00852856f $X=0.7 $Y=1.96 $X2=0 $Y2=0
cc_92 N_A_105_352#_c_101_n N_VPWR_c_209_n 0.00702461f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_93 N_A_105_352#_c_101_n N_VPWR_c_204_n 0.0129385f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_94 N_A_105_352#_c_104_n N_VPWR_c_204_n 0.0104443f $X=0.7 $Y=1.96 $X2=0 $Y2=0
cc_95 N_A_105_352#_c_101_n N_Y_c_237_n 0.00125894f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_105_352#_c_94_n N_Y_c_237_n 0.00886537f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_105_352#_c_95_n N_Y_c_237_n 0.0187522f $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_105_352#_c_96_n N_Y_c_237_n 0.00844148f $X=1.535 $Y=1.202 $X2=0 $Y2=0
cc_99 N_A_105_352#_c_97_n N_Y_c_237_n 0.0333811f $X=0.917 $Y=1.142 $X2=0 $Y2=0
cc_100 N_A_105_352#_c_99_n N_Y_c_237_n 0.0261377f $X=0.775 $Y=0.66 $X2=0 $Y2=0
cc_101 N_A_105_352#_c_101_n N_Y_c_239_n 0.0216819f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_105_352#_c_95_n N_Y_c_239_n 0.0011741f $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_105_352#_c_96_n N_Y_c_239_n 5.91391e-19 $X=1.535 $Y=1.202 $X2=0 $Y2=0
cc_104 N_A_105_352#_c_105_n N_Y_c_239_n 0.00794898f $X=0.917 $Y=1.535 $X2=0
+ $Y2=0
cc_105 N_A_105_352#_c_98_n N_Y_c_239_n 0.0077217f $X=0.98 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_105_352#_c_94_n N_VGND_c_273_n 0.00585385f $X=1.56 $Y=0.995 $X2=0
+ $Y2=0
cc_107 N_A_105_352#_c_99_n N_VGND_c_273_n 0.00685041f $X=0.775 $Y=0.66 $X2=0
+ $Y2=0
cc_108 N_A_105_352#_c_94_n N_VGND_c_276_n 0.0123242f $X=1.56 $Y=0.995 $X2=0
+ $Y2=0
cc_109 N_A_105_352#_c_99_n N_VGND_c_276_n 0.00866271f $X=0.775 $Y=0.66 $X2=0
+ $Y2=0
cc_110 N_A_105_352#_c_94_n N_A_327_47#_c_308_n 2.01734e-19 $X=1.56 $Y=0.995
+ $X2=0 $Y2=0
cc_111 N_A2_c_153_n N_A1_c_183_n 0.0743574f $X=2.035 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_112 A2 N_A1_c_183_n 6.84e-19 $X=2.01 $Y=1.19 $X2=-0.19 $Y2=-0.24
cc_113 N_A2_c_154_n N_A1_c_184_n 0.0205136f $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A2_c_153_n A1 8.91766e-19 $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_115 A2 A1 0.017913f $X=2.01 $Y=1.19 $X2=0 $Y2=0
cc_116 N_A2_c_153_n N_VPWR_c_207_n 0.00234541f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A2_c_153_n N_VPWR_c_209_n 0.00429201f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A2_c_153_n N_VPWR_c_204_n 0.00616095f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A2_c_153_n N_Y_c_237_n 0.0013144f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_120 A2 N_Y_c_237_n 0.0130926f $X=2.01 $Y=1.19 $X2=0 $Y2=0
cc_121 N_A2_c_153_n N_Y_c_239_n 0.00959919f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_122 A2 N_Y_c_239_n 0.0350129f $X=2.01 $Y=1.19 $X2=0 $Y2=0
cc_123 N_A2_c_153_n Y 0.0196172f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A2_c_154_n N_VGND_c_272_n 0.00412826f $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A2_c_154_n N_VGND_c_273_n 0.00439206f $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A2_c_154_n N_VGND_c_276_n 0.00631555f $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A2_c_153_n N_A_327_47#_c_307_n 4.31598e-19 $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A2_c_154_n N_A_327_47#_c_307_n 0.0106913f $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_129 A2 N_A_327_47#_c_307_n 0.0159183f $X=2.01 $Y=1.19 $X2=0 $Y2=0
cc_130 N_A2_c_153_n N_A_327_47#_c_308_n 0.00293476f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_131 A2 N_A_327_47#_c_308_n 0.0246764f $X=2.01 $Y=1.19 $X2=0 $Y2=0
cc_132 N_A2_c_154_n N_A_327_47#_c_309_n 6.1012e-19 $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A1_c_183_n N_VPWR_c_207_n 0.0315511f $X=2.495 $Y=1.41 $X2=0 $Y2=0
cc_134 A1 N_VPWR_c_207_n 0.0258868f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_135 N_A1_c_183_n N_VPWR_c_209_n 0.00251889f $X=2.495 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A1_c_183_n N_VPWR_c_204_n 0.0047299f $X=2.495 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A1_c_183_n N_Y_c_239_n 0.00137626f $X=2.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A1_c_184_n N_VGND_c_272_n 0.00384701f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A1_c_184_n N_VGND_c_275_n 0.00398883f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A1_c_184_n N_VGND_c_276_n 0.0068457f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A1_c_183_n N_A_327_47#_c_307_n 0.00327376f $X=2.495 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A1_c_184_n N_A_327_47#_c_307_n 0.00883093f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_143 A1 N_A_327_47#_c_307_n 0.0436897f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A1_c_184_n N_A_327_47#_c_309_n 0.00859991f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_145 N_VPWR_c_204_n N_Y_M1007_d 0.00290066f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_146 N_VPWR_M1006_d N_Y_c_239_n 0.00336693f $X=1.025 $Y=1.76 $X2=0 $Y2=0
cc_147 N_VPWR_c_205_n N_Y_c_239_n 0.00939049f $X=1.235 $Y=1.96 $X2=0 $Y2=0
cc_148 N_VPWR_c_209_n Y 0.0314093f $X=2.47 $Y=2.72 $X2=0 $Y2=0
cc_149 N_VPWR_c_204_n Y 0.0190535f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_150 N_VPWR_c_204_n A_425_297# 0.0109731f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_151 N_Y_c_237_n N_VGND_c_273_n 0.0144241f $X=1.35 $Y=0.545 $X2=0 $Y2=0
cc_152 N_Y_M1004_s N_VGND_c_276_n 0.00570496f $X=1.175 $Y=0.235 $X2=0 $Y2=0
cc_153 N_Y_c_237_n N_VGND_c_276_n 0.00839556f $X=1.35 $Y=0.545 $X2=0 $Y2=0
cc_154 N_Y_c_237_n N_A_327_47#_c_308_n 0.00153713f $X=1.35 $Y=0.545 $X2=0 $Y2=0
cc_155 N_Y_c_239_n N_A_327_47#_c_308_n 0.00132365f $X=1.895 $Y=1.625 $X2=0 $Y2=0
cc_156 N_VGND_c_276_n N_A_327_47#_M1004_d 0.00303164f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_157 N_VGND_c_276_n N_A_327_47#_M1005_d 0.00209863f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_158 N_VGND_c_273_n N_A_327_47#_c_325_n 0.0198051f $X=2.195 $Y=0 $X2=0 $Y2=0
cc_159 N_VGND_c_276_n N_A_327_47#_c_325_n 0.0126169f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_160 N_VGND_M1003_d N_A_327_47#_c_307_n 0.00261935f $X=2.135 $Y=0.235 $X2=0
+ $Y2=0
cc_161 N_VGND_c_272_n N_A_327_47#_c_307_n 0.0125492f $X=2.28 $Y=0.39 $X2=0 $Y2=0
cc_162 N_VGND_c_273_n N_A_327_47#_c_307_n 0.00253972f $X=2.195 $Y=0 $X2=0 $Y2=0
cc_163 N_VGND_c_275_n N_A_327_47#_c_307_n 0.00194552f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_164 N_VGND_c_276_n N_A_327_47#_c_307_n 0.00984903f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_165 N_VGND_c_272_n N_A_327_47#_c_309_n 0.0212768f $X=2.28 $Y=0.39 $X2=0 $Y2=0
cc_166 N_VGND_c_275_n N_A_327_47#_c_309_n 0.022204f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_167 N_VGND_c_276_n N_A_327_47#_c_309_n 0.0139896f $X=2.99 $Y=0 $X2=0 $Y2=0
