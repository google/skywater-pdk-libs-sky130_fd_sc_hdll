* File: sky130_fd_sc_hdll__o221a_4.spice
* Created: Thu Aug 27 19:20:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o221a_4.pex.spice"
.subckt sky130_fd_sc_hdll__o221a_4  VNB VPB C1 B1 B2 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1002 N_A_27_47#_M1002_d N_C1_M1002_g N_A_117_297#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1019 N_A_27_47#_M1019_d N_C1_M1019_g N_A_117_297#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1014 N_A_27_47#_M1019_d N_B1_M1014_g N_A_307_47#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1015 N_A_307_47#_M1014_s N_B2_M1015_g N_A_27_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1024 N_A_307_47#_M1024_d N_B2_M1024_g N_A_27_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1027 N_A_27_47#_M1027_d N_B1_M1027_g N_A_307_47#_M1024_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_307_47#_M1000_d N_A1_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1018 N_A_307_47#_M1000_d N_A2_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1025 N_A_307_47#_M1025_d N_A2_M1025_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1010 N_A_307_47#_M1025_d N_A1_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_117_297#_M1003_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1003_d N_A_117_297#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1008_d N_A_117_297#_M1008_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1021 N_X_M1008_d N_A_117_297#_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_C1_M1001_g N_A_117_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90006.8 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_C1_M1009_g N_A_117_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90006.3 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1009_d N_B1_M1006_g N_A_305_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90005.9 A=0.18 P=2.36 MULT=1
MM1011 N_A_305_297#_M1006_s N_B2_M1011_g N_A_117_297#_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90005.4 A=0.18 P=2.36 MULT=1
MM1016 N_A_305_297#_M1016_d N_B2_M1016_g N_A_117_297#_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1022_d N_B1_M1022_g N_A_305_297#_M1016_d VPB PHIGHVT L=0.18 W=1
+ AD=0.405 AS=0.145 PD=1.81 PS=1.29 NRD=2.9353 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90004.5 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1022_d N_A1_M1005_g N_A_785_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.405 AS=0.145 PD=1.81 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1013 N_A_785_297#_M1005_s N_A2_M1013_g N_A_117_297#_M1013_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004 SB=90003 A=0.18 P=2.36 MULT=1
MM1020 N_A_785_297#_M1020_d N_A2_M1020_g N_A_117_297#_M1013_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.5 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1026 N_VPWR_M1026_d N_A1_M1026_g N_A_785_297#_M1020_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.9 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1004 N_X_M1004_d N_A_117_297#_M1004_g N_VPWR_M1026_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.4 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1012 N_X_M1004_d N_A_117_297#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.9 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1017 N_X_M1017_d N_A_117_297#_M1017_g N_VPWR_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.3 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1023 N_X_M1017_d N_A_117_297#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.8 SB=90000.2 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=13.161 P=19.61
pX29_noxref noxref_16 B1 B1 PROBETYPE=1
pX30_noxref noxref_17 B2 B2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o221a_4.pxi.spice"
*
.ends
*
*
