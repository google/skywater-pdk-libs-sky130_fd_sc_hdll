* NGSPICE file created from sky130_fd_sc_hdll__nor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nor3_2 A B C VGND VNB VPB VPWR Y
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u
M1001 VGND C Y VNB nshort w=650000u l=150000u
+  ad=8.6125e+11p pd=9.15e+06u as=7.215e+11p ps=6.12e+06u
M1002 a_27_297# B a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.3e+11p ps=7.66e+06u
M1003 a_309_297# C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 a_309_297# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y C a_309_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

