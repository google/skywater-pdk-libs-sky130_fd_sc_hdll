* File: sky130_fd_sc_hdll__inputiso1n_1.spice
* Created: Thu Aug 27 19:08:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__inputiso1n_1.pex.spice"
.subckt sky130_fd_sc_hdll__inputiso1n_1  VNB VPB SLEEP_B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* SLEEP_B	SLEEP_B
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_SLEEP_B_M1000_g N_A_27_53#_M1000_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1806 AS=0.1302 PD=1.28 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_229_297#_M1006_d N_A_27_53#_M1006_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1806 PD=0.74 PS=1.28 NRD=0 NRS=30 M=1 R=2.8 SA=75001.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_229_297#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0927336 AS=0.0672 PD=0.816449 PS=0.74 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75001.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_229_297#_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.143516 PD=1.86 PS=1.26355 NRD=0.912 NRS=11.988 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_53#_M1002_d N_SLEEP_B_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1218 AS=0.1134 PD=1.42 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1003 A_319_297# N_A_27_53#_M1003_g N_A_229_297#_M1003_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=42.1974 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g A_319_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0918972 AS=0.0609 PD=0.804507 PS=0.71 NRD=76.83 NRS=42.1974 M=1 R=2.33333
+ SA=90000.6 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1007 N_X_M1007_d N_A_229_297#_M1007_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.218803 PD=2.58 PS=1.91549 NRD=2.9353 NRS=1.9503 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_55 VPB 0 8.49032e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__inputiso1n_1.pxi.spice"
*
.ends
*
*
