* File: sky130_fd_sc_hdll__a21oi_1.pxi.spice
* Created: Wed Sep  2 08:17:41 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21OI_1%B1 N_B1_c_38_n N_B1_M1000_g N_B1_c_35_n
+ N_B1_M1001_g B1 B1 N_B1_c_37_n PM_SKY130_FD_SC_HDLL__A21OI_1%B1
x_PM_SKY130_FD_SC_HDLL__A21OI_1%A1 N_A1_c_63_n N_A1_M1003_g N_A1_c_64_n
+ N_A1_M1002_g A1 A1 A1 A1 N_A1_c_66_n PM_SKY130_FD_SC_HDLL__A21OI_1%A1
x_PM_SKY130_FD_SC_HDLL__A21OI_1%A2 N_A2_c_101_n N_A2_M1005_g N_A2_c_103_n
+ N_A2_M1004_g A2 N_A2_c_102_n A2 PM_SKY130_FD_SC_HDLL__A21OI_1%A2
x_PM_SKY130_FD_SC_HDLL__A21OI_1%Y N_Y_M1001_d N_Y_M1000_s N_Y_c_126_n
+ N_Y_c_133_n Y Y PM_SKY130_FD_SC_HDLL__A21OI_1%Y
x_PM_SKY130_FD_SC_HDLL__A21OI_1%A_121_297# N_A_121_297#_M1000_d
+ N_A_121_297#_M1004_d N_A_121_297#_c_153_n N_A_121_297#_c_152_n
+ N_A_121_297#_c_150_n N_A_121_297#_c_151_n
+ PM_SKY130_FD_SC_HDLL__A21OI_1%A_121_297#
x_PM_SKY130_FD_SC_HDLL__A21OI_1%VPWR N_VPWR_M1003_d N_VPWR_c_179_n VPWR
+ N_VPWR_c_180_n N_VPWR_c_181_n N_VPWR_c_178_n N_VPWR_c_183_n
+ PM_SKY130_FD_SC_HDLL__A21OI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A21OI_1%VGND N_VGND_M1001_s N_VGND_M1005_d
+ N_VGND_c_207_n N_VGND_c_208_n N_VGND_c_209_n VGND N_VGND_c_210_n
+ N_VGND_c_211_n N_VGND_c_212_n N_VGND_c_213_n
+ PM_SKY130_FD_SC_HDLL__A21OI_1%VGND
cc_1 VNB N_B1_c_35_n 0.0193645f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB B1 0.0240596f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_B1_c_37_n 0.0405658f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_4 VNB N_A1_c_63_n 0.0254906f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_5 VNB N_A1_c_64_n 0.0165891f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_6 VNB A1 0.0013765f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_7 VNB N_A1_c_66_n 0.00233559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A2_c_101_n 0.0224192f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_9 VNB N_A2_c_102_n 0.0464807f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_Y_c_126_n 0.00268807f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_11 VNB N_VPWR_c_178_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_207_n 0.0119672f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_13 VNB N_VGND_c_208_n 0.0151005f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_209_n 0.028986f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_15 VNB N_VGND_c_210_n 0.0322453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_211_n 0.0150312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_212_n 0.154839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_213_n 0.00577043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VPB N_B1_c_38_n 0.0208881f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_20 VPB B1 0.00295004f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_21 VPB N_B1_c_37_n 0.0179665f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_22 VPB N_A1_c_63_n 0.0269329f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_23 VPB N_A1_c_66_n 0.00125452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_A2_c_103_n 0.0214614f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_25 VPB N_A2_c_102_n 0.0171244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_Y_c_126_n 0.0101665f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_27 VPB Y 0.0301226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_121_297#_c_150_n 0.022587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_A_121_297#_c_151_n 0.0171747f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.202
cc_30 VPB N_VPWR_c_179_n 0.0048706f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_31 VPB N_VPWR_c_180_n 0.0315326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_181_n 0.0286457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_178_n 0.0570554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_183_n 0.00372273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 N_B1_c_38_n N_A1_c_63_n 0.0196871f $X=0.515 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_36 N_B1_c_37_n N_A1_c_63_n 0.0203458f $X=0.515 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_37 N_B1_c_35_n N_A1_c_64_n 0.0172043f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_38 N_B1_c_35_n A1 2.4351e-19 $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_39 N_B1_c_37_n N_A1_c_66_n 3.13134e-19 $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_40 N_B1_c_38_n N_Y_c_126_n 0.0217443f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_41 N_B1_c_35_n N_Y_c_126_n 0.00438956f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_42 B1 N_Y_c_126_n 0.0550022f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_43 N_B1_c_37_n N_Y_c_126_n 0.0185725f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_44 N_B1_c_35_n N_Y_c_133_n 0.00765221f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_45 B1 N_Y_c_133_n 0.0114674f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_46 N_B1_c_38_n N_A_121_297#_c_152_n 0.0100219f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_47 N_B1_c_38_n N_VPWR_c_180_n 0.00604689f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_48 N_B1_c_38_n N_VPWR_c_178_n 0.0113332f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_49 B1 N_VGND_M1001_s 0.00520684f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_50 B1 N_VGND_c_207_n 2.61981e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_51 N_B1_c_35_n N_VGND_c_208_n 0.00478313f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_52 B1 N_VGND_c_208_n 0.0165104f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_53 N_B1_c_37_n N_VGND_c_208_n 0.00357437f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_54 N_B1_c_35_n N_VGND_c_210_n 0.00468917f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_55 N_B1_c_35_n N_VGND_c_212_n 0.00812511f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_56 B1 N_VGND_c_212_n 0.00158303f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_A1_c_64_n N_A2_c_101_n 0.0350147f $X=1.02 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_58 A1 N_A2_c_101_n 0.00815043f $X=1.09 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_59 N_A1_c_63_n N_A2_c_103_n 0.0352145f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A1_c_63_n A2 2.77823e-19 $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A1_c_66_n A2 0.0210026f $X=1.18 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A1_c_63_n N_A2_c_102_n 0.0250003f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_63 N_A1_c_66_n N_A2_c_102_n 0.00260893f $X=1.18 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A1_c_63_n N_Y_c_126_n 0.00729299f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A1_c_64_n N_Y_c_126_n 0.00127053f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_66 A1 N_Y_c_126_n 0.00756136f $X=1.09 $Y=0.425 $X2=0 $Y2=0
cc_67 N_A1_c_66_n N_Y_c_126_n 0.0256541f $X=1.18 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A1_c_63_n N_Y_c_133_n 9.44913e-19 $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A1_c_64_n N_Y_c_133_n 0.00456065f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_70 A1 N_Y_c_133_n 0.0320402f $X=1.09 $Y=0.425 $X2=0 $Y2=0
cc_71 N_A1_c_63_n N_A_121_297#_c_153_n 0.0224781f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A1_c_66_n N_A_121_297#_c_153_n 0.0243825f $X=1.18 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A1_c_63_n N_A_121_297#_c_152_n 0.00800211f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A1_c_66_n N_A_121_297#_c_152_n 0.00121593f $X=1.18 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A1_c_63_n N_A_121_297#_c_151_n 5.44221e-19 $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A1_c_63_n N_VPWR_c_179_n 0.0027771f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A1_c_63_n N_VPWR_c_180_n 0.00513064f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A1_c_63_n N_VPWR_c_178_n 0.00687734f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A1_c_64_n N_VGND_c_210_n 0.00545968f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_80 A1 N_VGND_c_210_n 0.00784567f $X=1.09 $Y=0.425 $X2=0 $Y2=0
cc_81 N_A1_c_64_n N_VGND_c_212_n 0.0100218f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_82 A1 N_VGND_c_212_n 0.00804886f $X=1.09 $Y=0.425 $X2=0 $Y2=0
cc_83 A1 A_219_47# 0.00761283f $X=1.09 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_84 N_A2_c_103_n N_A_121_297#_c_153_n 0.0202731f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A2_c_103_n N_A_121_297#_c_152_n 5.06552e-19 $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A2_c_103_n N_A_121_297#_c_150_n 0.004385f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_87 A2 N_A_121_297#_c_150_n 0.0190296f $X=1.585 $Y=1.105 $X2=0 $Y2=0
cc_88 N_A2_c_102_n N_A_121_297#_c_150_n 0.00684083f $X=1.49 $Y=1.202 $X2=0 $Y2=0
cc_89 N_A2_c_103_n N_A_121_297#_c_151_n 0.00792688f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A2_c_103_n N_VPWR_c_179_n 0.00404464f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A2_c_103_n N_VPWR_c_181_n 0.00489915f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A2_c_103_n N_VPWR_c_178_n 0.00787416f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A2_c_101_n N_VGND_c_209_n 0.00813487f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_94 A2 N_VGND_c_209_n 0.0176537f $X=1.585 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A2_c_102_n N_VGND_c_209_n 0.00694792f $X=1.49 $Y=1.202 $X2=0 $Y2=0
cc_96 N_A2_c_101_n N_VGND_c_210_n 0.00585385f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A2_c_101_n N_VGND_c_212_n 0.0121693f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_98 N_Y_c_126_n N_A_121_297#_M1000_d 0.0029996f $X=0.617 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_99 N_Y_c_126_n N_A_121_297#_c_152_n 0.0103775f $X=0.617 $Y=1.495 $X2=0 $Y2=0
cc_100 Y N_VPWR_c_180_n 0.0180804f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_101 N_Y_M1000_s N_VPWR_c_178_n 0.004171f $X=0.15 $Y=1.485 $X2=0 $Y2=0
cc_102 Y N_VPWR_c_178_n 0.0104586f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_103 N_Y_c_133_n N_VGND_c_210_n 0.0160204f $X=0.772 $Y=0.645 $X2=0 $Y2=0
cc_104 N_Y_M1001_d N_VGND_c_212_n 0.00490202f $X=0.615 $Y=0.235 $X2=0 $Y2=0
cc_105 N_Y_c_133_n N_VGND_c_212_n 0.012285f $X=0.772 $Y=0.645 $X2=0 $Y2=0
cc_106 N_A_121_297#_c_153_n N_VPWR_M1003_d 0.00599137f $X=1.515 $Y=1.775
+ $X2=-0.19 $Y2=1.305
cc_107 N_A_121_297#_c_153_n N_VPWR_c_179_n 0.016034f $X=1.515 $Y=1.775 $X2=0
+ $Y2=0
cc_108 N_A_121_297#_c_151_n N_VPWR_c_179_n 0.0187589f $X=1.73 $Y=2.33 $X2=0
+ $Y2=0
cc_109 N_A_121_297#_c_153_n N_VPWR_c_180_n 0.00297848f $X=1.515 $Y=1.775 $X2=0
+ $Y2=0
cc_110 N_A_121_297#_c_152_n N_VPWR_c_180_n 0.0210187f $X=0.92 $Y=1.775 $X2=0
+ $Y2=0
cc_111 N_A_121_297#_c_153_n N_VPWR_c_181_n 0.00236055f $X=1.515 $Y=1.775 $X2=0
+ $Y2=0
cc_112 N_A_121_297#_c_151_n N_VPWR_c_181_n 0.0230089f $X=1.73 $Y=2.33 $X2=0
+ $Y2=0
cc_113 N_A_121_297#_M1000_d N_VPWR_c_178_n 0.00239662f $X=0.605 $Y=1.485 $X2=0
+ $Y2=0
cc_114 N_A_121_297#_M1004_d N_VPWR_c_178_n 0.00221957f $X=1.58 $Y=1.485 $X2=0
+ $Y2=0
cc_115 N_A_121_297#_c_153_n N_VPWR_c_178_n 0.0107109f $X=1.515 $Y=1.775 $X2=0
+ $Y2=0
cc_116 N_A_121_297#_c_152_n N_VPWR_c_178_n 0.0140066f $X=0.92 $Y=1.775 $X2=0
+ $Y2=0
cc_117 N_A_121_297#_c_151_n N_VPWR_c_178_n 0.014122f $X=1.73 $Y=2.33 $X2=0 $Y2=0
cc_118 N_VGND_c_212_n A_219_47# 0.00580835f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24
