* File: sky130_fd_sc_hdll__nand3b_4.spice
* Created: Wed Sep  2 08:38:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand3b_4.pex.spice"
.subckt sky130_fd_sc_hdll__nand3b_4  VNB VPB A_N B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_A_N_M1023_g N_A_27_47#_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.169 PD=1.92 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_225_47#_M1005_d N_A_27_47#_M1005_g N_Y_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1006 N_A_225_47#_M1006_d N_A_27_47#_M1006_g N_Y_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75003 A=0.0975 P=1.6 MULT=1
MM1008 N_A_225_47#_M1006_d N_A_27_47#_M1008_g N_Y_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1018 N_A_225_47#_M1018_d N_A_27_47#_M1018_g N_Y_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1003 N_A_225_47#_M1018_d N_B_M1003_g N_A_683_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1004 N_A_225_47#_M1004_d N_B_M1004_g N_A_683_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.5 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1016 N_A_225_47#_M1004_d N_B_M1016_g N_A_683_47#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1024 N_A_225_47#_M1024_d N_B_M1024_g N_A_683_47#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_C_M1011_g N_A_683_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_C_M1012_g N_A_683_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1012_d N_C_M1019_g N_A_683_47#_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1022_d N_C_M1022_g N_A_683_47#_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.234 AS=0.104 PD=2.02 PS=0.97 NRD=13.836 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_A_N_M1007_g N_A_27_47#_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.27 PD=2.54 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_27_47#_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_27_47#_M1009_g N_Y_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1009_d N_A_27_47#_M1014_g N_Y_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_A_27_47#_M1020_g N_Y_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VPWR_M1020_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1013 N_Y_M1001_d N_B_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.5
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1017 N_Y_M1017_d N_B_M1017_g N_VPWR_M1013_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1025 N_Y_M1017_d N_B_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1010 N_Y_M1000_d N_C_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1015_d N_C_M1015_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1021 N_Y_M1015_d N_C_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.37 PD=1.29 PS=2.74 NRD=0.9653 NRS=16.7253 M=1 R=5.55556 SA=90001.6
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX26_noxref VNB VPB NWDIODE A=13.161 P=19.61
*
.include "sky130_fd_sc_hdll__nand3b_4.pxi.spice"
*
.ends
*
*
