* File: sky130_fd_sc_hdll__bufbuf_8.spice
* Created: Thu Aug 27 19:00:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__bufbuf_8.pex.spice"
.subckt sky130_fd_sc_hdll__bufbuf_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_M1018_g N_A_27_47#_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0914579 AS=0.1302 PD=0.812523 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1024 N_A_224_297#_M1024_d N_A_27_47#_M1024_g N_VGND_M1018_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.141542 PD=1.82 PS=1.25748 NRD=0 NRS=20.304 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_224_297#_M1005_g N_A_338_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1005_d N_A_224_297#_M1011_g N_A_338_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_224_297#_M1012_g N_A_338_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75003.9 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1012_d N_A_338_47#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_338_47#_M1003_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1003_d N_A_338_47#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_338_47#_M1007_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1007_d N_A_338_47#_M1013_g N_X_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_338_47#_M1015_g N_X_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.9
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1015_d N_A_338_47#_M1020_g N_X_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.4
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1023_d N_A_338_47#_M1023_g N_X_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.126595 AS=0.1728 PD=1.05756 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1021 N_A_224_297#_M1021_d N_A_27_47#_M1021_g N_VPWR_M1010_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.197805 PD=2.54 PS=1.65244 NRD=0.9653 NRS=13.7703 M=1
+ R=5.55556 SA=90000.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_224_297#_M1009_g N_A_338_47#_M1009_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1009_d N_A_224_297#_M1014_g N_A_338_47#_M1014_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1017_d N_A_224_297#_M1017_g N_A_338_47#_M1014_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001.1 SB=90003.9 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1017_d N_A_338_47#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_338_47#_M1002_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90003 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1002_d N_A_338_47#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_338_47#_M1008_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1008_d N_A_338_47#_M1016_g N_X_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1019_d N_A_338_47#_M1019_g N_X_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.9 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1019_d N_A_338_47#_M1022_g N_X_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1025 N_VPWR_M1025_d N_A_338_47#_M1025_g N_X_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.9 SB=90000.2 A=0.18 P=2.36 MULT=1
DX26_noxref VNB VPB NWDIODE A=12.4227 P=18.69
pX27_noxref noxref_10 X X PROBETYPE=1
pX28_noxref noxref_11 X X PROBETYPE=1
c_128 VPB 0 1.95897e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__bufbuf_8.pxi.spice"
*
.ends
*
*
