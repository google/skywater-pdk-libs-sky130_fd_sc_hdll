* File: sky130_fd_sc_hdll__o211a_2.pxi.spice
* Created: Thu Aug 27 19:18:17 2020
* 
x_PM_SKY130_FD_SC_HDLL__O211A_2%C1 N_C1_c_59_n N_C1_M1002_g N_C1_c_60_n
+ N_C1_M1001_g C1 C1 PM_SKY130_FD_SC_HDLL__O211A_2%C1
x_PM_SKY130_FD_SC_HDLL__O211A_2%B1 N_B1_c_80_n N_B1_M1004_g N_B1_c_81_n
+ N_B1_M1008_g B1 B1 PM_SKY130_FD_SC_HDLL__O211A_2%B1
x_PM_SKY130_FD_SC_HDLL__O211A_2%A2 N_A2_c_109_n N_A2_M1010_g N_A2_c_110_n
+ N_A2_M1005_g A2 N_A2_c_111_n A2 PM_SKY130_FD_SC_HDLL__O211A_2%A2
x_PM_SKY130_FD_SC_HDLL__O211A_2%A1 N_A1_c_136_n N_A1_M1011_g N_A1_c_137_n
+ N_A1_M1009_g A1 A1 PM_SKY130_FD_SC_HDLL__O211A_2%A1
x_PM_SKY130_FD_SC_HDLL__O211A_2%A_27_47# N_A_27_47#_M1001_s N_A_27_47#_M1002_s
+ N_A_27_47#_M1008_d N_A_27_47#_c_167_n N_A_27_47#_M1006_g N_A_27_47#_c_172_n
+ N_A_27_47#_M1000_g N_A_27_47#_c_173_n N_A_27_47#_M1003_g N_A_27_47#_c_168_n
+ N_A_27_47#_M1007_g N_A_27_47#_c_174_n N_A_27_47#_c_169_n N_A_27_47#_c_190_n
+ N_A_27_47#_c_176_n N_A_27_47#_c_219_p N_A_27_47#_c_195_n N_A_27_47#_c_203_n
+ N_A_27_47#_c_204_n N_A_27_47#_c_177_n N_A_27_47#_c_170_n N_A_27_47#_c_193_n
+ N_A_27_47#_c_171_n PM_SKY130_FD_SC_HDLL__O211A_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O211A_2%VPWR N_VPWR_M1002_d N_VPWR_M1011_d
+ N_VPWR_M1003_d N_VPWR_c_259_n N_VPWR_c_260_n N_VPWR_c_261_n VPWR
+ N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_264_n N_VPWR_c_258_n N_VPWR_c_266_n
+ N_VPWR_c_267_n N_VPWR_c_268_n PM_SKY130_FD_SC_HDLL__O211A_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O211A_2%X N_X_M1006_d N_X_M1000_s N_X_c_335_n
+ N_X_c_315_n N_X_c_321_n N_X_c_323_n N_X_c_317_n X N_X_c_313_n X
+ PM_SKY130_FD_SC_HDLL__O211A_2%X
x_PM_SKY130_FD_SC_HDLL__O211A_2%A_206_47# N_A_206_47#_M1004_d
+ N_A_206_47#_M1005_d N_A_206_47#_c_360_n
+ PM_SKY130_FD_SC_HDLL__O211A_2%A_206_47#
x_PM_SKY130_FD_SC_HDLL__O211A_2%VGND N_VGND_M1005_s N_VGND_M1009_d
+ N_VGND_M1007_s N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n
+ N_VGND_c_384_n N_VGND_c_385_n VGND N_VGND_c_386_n N_VGND_c_387_n
+ N_VGND_c_388_n N_VGND_c_389_n PM_SKY130_FD_SC_HDLL__O211A_2%VGND
cc_1 VNB N_C1_c_59_n 0.0377383f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_2 VNB N_C1_c_60_n 0.0216657f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_3 VNB C1 0.011737f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_B1_c_80_n 0.0222863f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_5 VNB N_B1_c_81_n 0.0296502f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_6 VNB B1 0.00240786f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.16
cc_7 VNB N_A2_c_109_n 0.0314802f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_8 VNB N_A2_c_110_n 0.0225937f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_9 VNB N_A2_c_111_n 0.00290298f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_10 VNB N_A1_c_136_n 0.0251885f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_11 VNB N_A1_c_137_n 0.0174905f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_12 VNB A1 0.00563763f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_13 VNB N_A_27_47#_c_167_n 0.0177201f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_14 VNB N_A_27_47#_c_168_n 0.0202771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_169_n 0.00289902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_170_n 0.0239964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_171_n 0.044742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_258_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_313_n 0.0077428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB X 0.026374f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_206_47#_c_360_n 0.0128595f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_22 VNB N_VGND_c_380_n 0.00904014f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_23 VNB N_VGND_c_381_n 0.00452783f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_382_n 0.0162245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_383_n 0.00563028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_384_n 0.0190178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_385_n 0.00448835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_386_n 0.0429299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_387_n 0.0197271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_388_n 0.00641049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_389_n 0.222435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_C1_c_59_n 0.0386527f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_33 VPB C1 0.00101332f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_34 VPB N_B1_c_81_n 0.0341443f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_35 VPB B1 4.62185e-19 $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.16
cc_36 VPB N_A2_c_109_n 0.036226f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_37 VPB N_A2_c_111_n 0.00103114f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_38 VPB N_A1_c_136_n 0.0272796f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_39 VPB A1 0.00167584f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_40 VPB N_A_27_47#_c_172_n 0.0171083f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_41 VPB N_A_27_47#_c_173_n 0.0182903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_174_n 0.0269609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_169_n 0.00167261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_47#_c_176_n 0.0111775f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_177_n 0.00611171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_171_n 0.0240767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_259_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_48 VPB N_VPWR_c_260_n 6.85619e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_261_n 0.0141218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_262_n 0.0153288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_263_n 0.0381016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_264_n 0.0112609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_258_n 0.0459914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_266_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_267_n 0.00666211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_268_n 0.00868132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_X_c_315_n 0.00917881f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_58 VPB X 0.0271672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 N_C1_c_60_n N_B1_c_80_n 0.0280466f $X=0.525 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_60 N_C1_c_59_n N_B1_c_81_n 0.050064f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_61 N_C1_c_59_n B1 2.93152e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_62 N_C1_c_59_n N_A_27_47#_c_169_n 0.0195612f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_63 N_C1_c_60_n N_A_27_47#_c_169_n 0.00890804f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_64 C1 N_A_27_47#_c_169_n 0.0237386f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_65 N_C1_c_59_n N_A_27_47#_c_176_n 0.0286838f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_66 C1 N_A_27_47#_c_176_n 0.0191266f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_67 N_C1_c_59_n N_A_27_47#_c_170_n 0.00882475f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_68 N_C1_c_60_n N_A_27_47#_c_170_n 0.0148717f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_69 C1 N_A_27_47#_c_170_n 0.0216856f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_70 N_C1_c_59_n N_VPWR_c_259_n 0.0152888f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_71 N_C1_c_59_n N_VPWR_c_262_n 0.00447018f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_72 N_C1_c_59_n N_VPWR_c_258_n 0.00855297f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_73 N_C1_c_60_n N_VGND_c_386_n 0.00390689f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_74 N_C1_c_60_n N_VGND_c_389_n 0.0064453f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_75 N_B1_c_81_n N_A2_c_109_n 0.0143247f $X=0.98 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_76 B1 N_A2_c_109_n 0.00100644f $X=1.155 $Y=1.19 $X2=-0.19 $Y2=-0.24
cc_77 N_B1_c_81_n N_A2_c_111_n 0.00118216f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_78 B1 N_A2_c_111_n 0.0258174f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_79 N_B1_c_80_n N_A_27_47#_c_169_n 0.00834851f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B1_c_81_n N_A_27_47#_c_169_n 0.00233795f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_81 B1 N_A_27_47#_c_169_n 0.0256222f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_82 N_B1_c_81_n N_A_27_47#_c_190_n 0.025329f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_83 B1 N_A_27_47#_c_190_n 0.0115562f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_84 N_B1_c_80_n N_A_27_47#_c_170_n 0.00741427f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B1_c_81_n N_A_27_47#_c_193_n 0.00346193f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_86 B1 N_A_27_47#_c_193_n 0.0143708f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_87 N_B1_c_81_n N_VPWR_c_259_n 0.0119178f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B1_c_81_n N_VPWR_c_263_n 0.00642146f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B1_c_81_n N_VPWR_c_258_n 0.0121178f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B1_c_80_n N_A_206_47#_c_360_n 0.0064694f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B1_c_81_n N_A_206_47#_c_360_n 0.00554716f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_92 B1 N_A_206_47#_c_360_n 0.0260705f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_93 N_B1_c_80_n N_VGND_c_380_n 0.00800344f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B1_c_80_n N_VGND_c_386_n 0.00478524f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B1_c_80_n N_VGND_c_389_n 0.00895262f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A2_c_109_n N_A1_c_136_n 0.0953836f $X=1.94 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_97 N_A2_c_111_n N_A1_c_136_n 3.04787e-19 $X=1.81 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_98 N_A2_c_110_n N_A1_c_137_n 0.0223705f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A2_c_109_n A1 0.00245884f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A2_c_111_n A1 0.0227993f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A2_c_109_n N_A_27_47#_c_195_n 0.0238554f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A2_c_111_n N_A_27_47#_c_195_n 0.00752405f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A2_c_109_n N_A_27_47#_c_193_n 0.00555548f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A2_c_111_n N_A_27_47#_c_193_n 0.0236223f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A2_c_109_n N_VPWR_c_260_n 0.00285921f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A2_c_109_n N_VPWR_c_263_n 0.00702461f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A2_c_109_n N_VPWR_c_258_n 0.0139635f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A2_c_109_n N_A_206_47#_c_360_n 0.00674721f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A2_c_110_n N_A_206_47#_c_360_n 0.015527f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A2_c_111_n N_A_206_47#_c_360_n 0.0310041f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A2_c_110_n N_VGND_c_380_n 0.00345652f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A2_c_110_n N_VGND_c_384_n 0.00425094f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A2_c_110_n N_VGND_c_389_n 0.00708936f $X=1.965 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A1_c_137_n N_A_27_47#_c_167_n 0.0217484f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A1_c_136_n N_A_27_47#_c_172_n 0.0344846f $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A1_c_136_n N_A_27_47#_c_195_n 0.0219704f $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_117 A1 N_A_27_47#_c_195_n 0.0321415f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_118 N_A1_c_136_n N_A_27_47#_c_203_n 0.00106976f $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A1_c_136_n N_A_27_47#_c_204_n 3.53241e-19 $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_120 A1 N_A_27_47#_c_204_n 0.0274615f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A1_c_136_n N_A_27_47#_c_171_n 0.0222646f $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_122 A1 N_A_27_47#_c_171_n 0.00230199f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_123 N_A1_c_136_n N_VPWR_c_260_n 0.0277303f $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A1_c_136_n N_VPWR_c_263_n 0.00447018f $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A1_c_136_n N_VPWR_c_258_n 0.00758362f $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A1_c_137_n N_X_c_317_n 0.00101088f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A1_c_136_n N_A_206_47#_c_360_n 0.00248491f $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A1_c_137_n N_A_206_47#_c_360_n 0.00443781f $X=2.425 $Y=0.995 $X2=0
+ $Y2=0
cc_129 A1 N_A_206_47#_c_360_n 0.0137833f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_130 N_A1_c_136_n N_VGND_c_381_n 0.00124351f $X=2.35 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A1_c_137_n N_VGND_c_381_n 0.00165107f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_132 A1 N_VGND_c_381_n 0.00492859f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_133 N_A1_c_137_n N_VGND_c_384_n 0.0055867f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A1_c_137_n N_VGND_c_389_n 0.0100826f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_169_n N_VPWR_M1002_d 6.24752e-19 $X=0.645 $Y=1.51 $X2=-0.19
+ $Y2=-0.24
cc_136 N_A_27_47#_c_190_n N_VPWR_M1002_d 0.00366026f $X=1.125 $Y=1.637 $X2=-0.19
+ $Y2=-0.24
cc_137 N_A_27_47#_c_176_n N_VPWR_M1002_d 0.00153672f $X=0.76 $Y=1.637 $X2=-0.19
+ $Y2=-0.24
cc_138 N_A_27_47#_c_195_n N_VPWR_M1011_d 0.0103923f $X=2.855 $Y=1.622 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_c_176_n N_VPWR_c_259_n 0.0215081f $X=0.76 $Y=1.637 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_172_n N_VPWR_c_260_n 0.0184614f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_173_n N_VPWR_c_260_n 6.38696e-19 $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_195_n N_VPWR_c_260_n 0.0263794f $X=2.855 $Y=1.622 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_c_172_n N_VPWR_c_261_n 0.00681171f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_173_n N_VPWR_c_261_n 0.00327033f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_174_n N_VPWR_c_262_n 0.0185597f $X=0.26 $Y=1.82 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_219_p N_VPWR_c_263_n 0.0477916f $X=1.655 $Y=1.89 $X2=0 $Y2=0
cc_147 N_A_27_47#_M1002_s N_VPWR_c_258_n 0.00412552f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_M1008_d N_VPWR_c_258_n 0.00935418f $X=1.07 $Y=1.485 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_172_n N_VPWR_c_258_n 0.0113479f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_173_n N_VPWR_c_258_n 0.00389766f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_174_n N_VPWR_c_258_n 0.0101311f $X=0.26 $Y=1.82 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_219_p N_VPWR_c_258_n 0.0266834f $X=1.655 $Y=1.89 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_172_n N_VPWR_c_268_n 5.3452e-19 $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_173_n N_VPWR_c_268_n 0.0102824f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_195_n A_406_297# 0.00808081f $X=2.855 $Y=1.622 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A_27_47#_c_173_n N_X_c_315_n 0.0167137f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_177_n N_X_c_315_n 0.00654338f $X=3.38 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_171_n N_X_c_315_n 4.64597e-19 $X=3.42 $Y=1.202 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_177_n N_X_c_321_n 0.0066142f $X=3.38 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_171_n N_X_c_321_n 0.00114188f $X=3.42 $Y=1.202 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_168_n N_X_c_323_n 0.0117891f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_177_n N_X_c_323_n 0.0121177f $X=3.38 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_171_n N_X_c_323_n 0.00204241f $X=3.42 $Y=1.202 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_167_n N_X_c_317_n 0.00943863f $X=2.915 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_204_n N_X_c_317_n 0.00429544f $X=3.025 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_177_n N_X_c_317_n 0.0185703f $X=3.38 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_171_n N_X_c_317_n 0.00405352f $X=3.42 $Y=1.202 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_173_n X 0.0166417f $X=3.42 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_168_n X 0.00683075f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_177_n X 0.0240749f $X=3.38 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_171_n X 0.011647f $X=3.42 $Y=1.202 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_169_n A_120_47# 6.89224e-19 $X=0.645 $Y=1.51 $X2=-0.19
+ $Y2=-0.24
cc_173 N_A_27_47#_c_170_n A_120_47# 0.00580726f $X=0.265 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_27_47#_c_167_n N_A_206_47#_c_360_n 6.34793e-19 $X=2.915 $Y=0.995
+ $X2=0 $Y2=0
cc_175 N_A_27_47#_c_170_n N_A_206_47#_c_360_n 0.0164039f $X=0.265 $Y=0.38 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_167_n N_VGND_c_381_n 0.0039553f $X=2.915 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_168_n N_VGND_c_383_n 0.00867164f $X=3.425 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_170_n N_VGND_c_386_n 0.0314814f $X=0.265 $Y=0.38 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_167_n N_VGND_c_387_n 0.00518588f $X=2.915 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_168_n N_VGND_c_387_n 0.00422112f $X=3.425 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1001_s N_VGND_c_389_n 0.00256266f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_167_n N_VGND_c_389_n 0.0093943f $X=2.915 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_168_n N_VGND_c_389_n 0.00703456f $X=3.425 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_170_n N_VGND_c_389_n 0.0234808f $X=0.265 $Y=0.38 $X2=0 $Y2=0
cc_185 N_VPWR_c_258_n A_406_297# 0.00983149f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_186 N_VPWR_c_258_n N_X_M1000_s 0.00449905f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_187 N_VPWR_c_261_n N_X_c_335_n 0.0129667f $X=3.445 $Y=2.72 $X2=0 $Y2=0
cc_188 N_VPWR_c_258_n N_X_c_335_n 0.00719373f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_189 N_VPWR_M1003_d N_X_c_315_n 0.01373f $X=3.51 $Y=1.485 $X2=0 $Y2=0
cc_190 N_VPWR_c_261_n N_X_c_315_n 0.00236302f $X=3.445 $Y=2.72 $X2=0 $Y2=0
cc_191 N_VPWR_c_264_n N_X_c_315_n 0.00407384f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_258_n N_X_c_315_n 0.0121989f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_268_n N_X_c_315_n 0.023377f $X=3.66 $Y=2.34 $X2=0 $Y2=0
cc_194 N_VPWR_M1003_d X 0.00905309f $X=3.51 $Y=1.485 $X2=0 $Y2=0
cc_195 N_X_c_317_n N_A_206_47#_c_360_n 0.00442188f $X=3.16 $Y=0.36 $X2=0 $Y2=0
cc_196 N_X_c_323_n N_VGND_M1007_s 0.0100321f $X=3.765 $Y=0.7 $X2=0 $Y2=0
cc_197 N_X_c_313_n N_VGND_M1007_s 0.00532384f $X=3.9 $Y=0.785 $X2=0 $Y2=0
cc_198 X N_VGND_M1007_s 0.00253356f $X=3.915 $Y=0.85 $X2=0 $Y2=0
cc_199 N_X_c_317_n N_VGND_c_381_n 0.0206442f $X=3.16 $Y=0.36 $X2=0 $Y2=0
cc_200 N_X_c_313_n N_VGND_c_382_n 0.00328407f $X=3.9 $Y=0.785 $X2=0 $Y2=0
cc_201 N_X_c_323_n N_VGND_c_383_n 0.0157355f $X=3.765 $Y=0.7 $X2=0 $Y2=0
cc_202 N_X_c_313_n N_VGND_c_383_n 0.00912618f $X=3.9 $Y=0.785 $X2=0 $Y2=0
cc_203 N_X_c_323_n N_VGND_c_387_n 0.00327755f $X=3.765 $Y=0.7 $X2=0 $Y2=0
cc_204 N_X_c_317_n N_VGND_c_387_n 0.0230251f $X=3.16 $Y=0.36 $X2=0 $Y2=0
cc_205 N_X_M1006_d N_VGND_c_389_n 0.00294735f $X=2.99 $Y=0.235 $X2=0 $Y2=0
cc_206 N_X_c_323_n N_VGND_c_389_n 0.00653146f $X=3.765 $Y=0.7 $X2=0 $Y2=0
cc_207 N_X_c_317_n N_VGND_c_389_n 0.0141909f $X=3.16 $Y=0.36 $X2=0 $Y2=0
cc_208 N_X_c_313_n N_VGND_c_389_n 0.00550142f $X=3.9 $Y=0.785 $X2=0 $Y2=0
cc_209 A_120_47# N_VGND_c_389_n 0.00657074f $X=0.6 $Y=0.235 $X2=0.645 $Y2=1.637
cc_210 N_A_206_47#_c_360_n N_VGND_M1005_s 0.00621664f $X=2.21 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_211 N_A_206_47#_c_360_n N_VGND_c_380_n 0.022938f $X=2.21 $Y=0.73 $X2=0 $Y2=0
cc_212 N_A_206_47#_c_360_n N_VGND_c_384_n 0.00762762f $X=2.21 $Y=0.73 $X2=0
+ $Y2=0
cc_213 N_A_206_47#_c_360_n N_VGND_c_386_n 0.0102777f $X=2.21 $Y=0.73 $X2=0 $Y2=0
cc_214 N_A_206_47#_M1004_d N_VGND_c_389_n 0.00310899f $X=1.03 $Y=0.235 $X2=0
+ $Y2=0
cc_215 N_A_206_47#_M1005_d N_VGND_c_389_n 0.00362021f $X=2.04 $Y=0.235 $X2=0
+ $Y2=0
cc_216 N_A_206_47#_c_360_n N_VGND_c_389_n 0.0316647f $X=2.21 $Y=0.73 $X2=0 $Y2=0
