* File: sky130_fd_sc_hdll__a2bb2o_1.pxi.spice
* Created: Thu Aug 27 18:54:43 2020
* 
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%A_79_21# N_A_79_21#_M1002_d N_A_79_21#_M1000_s
+ N_A_79_21#_c_74_n N_A_79_21#_M1011_g N_A_79_21#_c_75_n N_A_79_21#_M1003_g
+ N_A_79_21#_c_76_n N_A_79_21#_c_82_n N_A_79_21#_c_129_p N_A_79_21#_c_83_n
+ N_A_79_21#_c_84_n N_A_79_21#_c_85_n N_A_79_21#_c_77_n N_A_79_21#_c_78_n
+ N_A_79_21#_c_87_n N_A_79_21#_c_79_n PM_SKY130_FD_SC_HDLL__A2BB2O_1%A_79_21#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%A1_N N_A1_N_c_165_n N_A1_N_M1004_g
+ N_A1_N_M1008_g A1_N A1_N PM_SKY130_FD_SC_HDLL__A2BB2O_1%A1_N
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%A2_N N_A2_N_c_195_n N_A2_N_M1009_g
+ N_A2_N_M1006_g A2_N A2_N PM_SKY130_FD_SC_HDLL__A2BB2O_1%A2_N
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%A_243_47# N_A_243_47#_M1008_d
+ N_A_243_47#_M1009_d N_A_243_47#_c_223_n N_A_243_47#_c_231_n
+ N_A_243_47#_M1000_g N_A_243_47#_M1002_g N_A_243_47#_c_225_n
+ N_A_243_47#_c_226_n N_A_243_47#_c_281_p N_A_243_47#_c_227_n
+ N_A_243_47#_c_228_n N_A_243_47#_c_232_n N_A_243_47#_c_229_n
+ N_A_243_47#_c_234_n PM_SKY130_FD_SC_HDLL__A2BB2O_1%A_243_47#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%B2 N_B2_M1001_g N_B2_c_293_n N_B2_c_294_n
+ N_B2_M1010_g B2 N_B2_c_292_n PM_SKY130_FD_SC_HDLL__A2BB2O_1%B2
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%B1 N_B1_M1007_g N_B1_c_333_n N_B1_c_334_n
+ N_B1_M1005_g B1 B1 B1 N_B1_c_332_n PM_SKY130_FD_SC_HDLL__A2BB2O_1%B1
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%X N_X_M1011_s N_X_M1003_s X X X
+ PM_SKY130_FD_SC_HDLL__A2BB2O_1%X
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%VPWR N_VPWR_M1003_d N_VPWR_M1010_d
+ N_VPWR_c_375_n N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n VPWR VPWR
+ N_VPWR_c_379_n VPWR N_VPWR_c_380_n N_VPWR_c_374_n N_VPWR_c_382_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%A_525_413# N_A_525_413#_M1000_d
+ N_A_525_413#_M1005_d N_A_525_413#_c_432_n N_A_525_413#_c_433_n
+ N_A_525_413#_c_434_n N_A_525_413#_c_435_n N_A_525_413#_c_439_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_1%A_525_413#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_1%VGND N_VGND_M1011_d N_VGND_M1006_d
+ N_VGND_M1007_d N_VGND_c_471_n N_VGND_c_472_n VGND VGND N_VGND_c_473_n VGND
+ N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_1%VGND
cc_1 VNB N_A_79_21#_c_74_n 0.0210357f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_75_n 0.0289922f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB N_A_79_21#_c_76_n 0.00199762f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_4 VNB N_A_79_21#_c_77_n 3.09199e-19 $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=1.895
cc_5 VNB N_A_79_21#_c_78_n 0.00130934f $X=-0.19 $Y=-0.24 $X2=2.77 $Y2=0.445
cc_6 VNB N_A_79_21#_c_79_n 0.0134631f $X=-0.19 $Y=-0.24 $X2=2.77 $Y2=0.785
cc_7 VNB N_A1_N_c_165_n 0.0207793f $X=-0.19 $Y=-0.24 $X2=2.635 $Y2=0.235
cc_8 VNB N_A1_N_M1008_g 0.0325896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB A1_N 0.00795212f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_A2_N_c_195_n 0.0219332f $X=-0.19 $Y=-0.24 $X2=2.635 $Y2=0.235
cc_11 VNB N_A2_N_M1006_g 0.0327467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB A2_N 0.00268823f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_13 VNB N_A_243_47#_c_223_n 0.00249771f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_14 VNB N_A_243_47#_M1002_g 0.0253447f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_15 VNB N_A_243_47#_c_225_n 0.0529479f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_16 VNB N_A_243_47#_c_226_n 0.0176332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_243_47#_c_227_n 0.0164821f $X=-0.19 $Y=-0.24 $X2=2.13 $Y2=2.285
cc_18 VNB N_A_243_47#_c_228_n 0.00698017f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=2.285
cc_19 VNB N_A_243_47#_c_229_n 0.00127188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B2_M1001_g 0.0438234f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB B2 0.00818883f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_22 VNB N_B2_c_292_n 0.00387715f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.805
cc_23 VNB N_B1_M1007_g 0.0355524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB B1 0.0142666f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_25 VNB N_B1_c_332_n 0.0325379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.046235f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_27 VNB N_VPWR_c_374_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_471_n 0.0158789f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_29 VNB N_VGND_c_472_n 0.022289f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_30 VNB N_VGND_c_473_n 0.0150788f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.89
cc_31 VNB N_VGND_c_474_n 0.031149f $X=-0.19 $Y=-0.24 $X2=2.365 $Y2=2.275
cc_32 VNB N_VGND_c_475_n 0.0111145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_476_n 0.0188556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_477_n 0.021135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_478_n 0.222597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_A_79_21#_c_75_n 0.0322703f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_37 VPB N_A_79_21#_c_76_n 0.00120716f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_38 VPB N_A_79_21#_c_82_n 0.00304263f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.89
cc_39 VPB N_A_79_21#_c_83_n 0.00868184f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=2.2
cc_40 VPB N_A_79_21#_c_84_n 0.0230789f $X=-0.19 $Y=1.305 $X2=2.13 $Y2=2.285
cc_41 VPB N_A_79_21#_c_85_n 0.004893f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=2.285
cc_42 VPB N_A_79_21#_c_77_n 0.00641068f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=1.895
cc_43 VPB N_A_79_21#_c_87_n 0.0166826f $X=-0.19 $Y=1.305 $X2=2.3 $Y2=2.275
cc_44 VPB N_A1_N_c_165_n 0.0243727f $X=-0.19 $Y=1.305 $X2=2.635 $Y2=0.235
cc_45 VPB A1_N 0.00279235f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_46 VPB N_A2_N_c_195_n 0.0281516f $X=-0.19 $Y=1.305 $X2=2.635 $Y2=0.235
cc_47 VPB A2_N 0.00309963f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_48 VPB N_A_243_47#_c_223_n 0.040005f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_49 VPB N_A_243_47#_c_231_n 0.0270873f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_50 VPB N_A_243_47#_c_232_n 0.0103582f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=0.87
cc_51 VPB N_A_243_47#_c_229_n 0.00466275f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_243_47#_c_234_n 0.00180429f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=0.785
cc_53 VPB N_B2_c_293_n 0.0141703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_B2_c_294_n 0.0214609f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_55 VPB B2 0.00335832f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_56 VPB N_B2_c_292_n 0.0249379f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.805
cc_57 VPB N_B1_c_333_n 0.0392684f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_B1_c_334_n 0.0260478f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_59 VPB B1 0.0147782f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_60 VPB N_B1_c_332_n 0.00384665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB X 0.0468332f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_62 VPB N_VPWR_c_375_n 0.00937122f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_63 VPB N_VPWR_c_376_n 0.00248358f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.805
cc_64 VPB N_VPWR_c_377_n 0.0562396f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_65 VPB N_VPWR_c_378_n 0.00378955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_379_n 0.0150576f $X=-0.19 $Y=1.305 $X2=2.13 $Y2=2.285
cc_67 VPB N_VPWR_c_380_n 0.0216505f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.16
cc_68 VPB N_VPWR_c_374_n 0.064228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_382_n 0.005797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_525_413#_c_432_n 3.53856e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_71 VPB N_A_525_413#_c_433_n 0.0253089f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_72 VPB N_A_525_413#_c_434_n 0.00570438f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_73 VPB N_A_525_413#_c_435_n 0.00268843f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.805
cc_74 N_A_79_21#_c_75_n N_A1_N_c_165_n 0.0369473f $X=0.495 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_79_21#_c_76_n N_A1_N_c_165_n 0.00539986f $X=0.6 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_79_21#_c_82_n N_A1_N_c_165_n 0.0118782f $X=1.155 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_79_21#_c_83_n N_A1_N_c_165_n 0.00274485f $X=1.265 $Y=2.2 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_79_21#_c_74_n N_A1_N_M1008_g 0.0166714f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_75_n A1_N 0.00221246f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_76_n A1_N 0.0338634f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_82_n A1_N 0.0194121f $X=1.155 $Y=1.89 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_82_n N_A2_N_c_195_n 0.00315845f $X=1.155 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_79_21#_c_83_n N_A2_N_c_195_n 0.0014283f $X=1.265 $Y=2.2 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_79_21#_c_84_n N_A2_N_c_195_n 0.00751161f $X=2.13 $Y=2.285 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_79_21#_c_87_n N_A2_N_c_195_n 0.00366357f $X=2.3 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_79_21#_c_77_n N_A_243_47#_c_223_n 0.0247748f $X=2.49 $Y=1.895 $X2=0
+ $Y2=0
cc_87 N_A_79_21#_c_87_n N_A_243_47#_c_231_n 0.0139179f $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_88 N_A_79_21#_c_78_n N_A_243_47#_M1002_g 5.47682e-19 $X=2.77 $Y=0.445 $X2=0
+ $Y2=0
cc_89 N_A_79_21#_c_79_n N_A_243_47#_M1002_g 0.0100975f $X=2.77 $Y=0.785 $X2=0
+ $Y2=0
cc_90 N_A_79_21#_c_77_n N_A_243_47#_c_225_n 0.00882306f $X=2.49 $Y=1.895 $X2=0
+ $Y2=0
cc_91 N_A_79_21#_c_87_n N_A_243_47#_c_225_n 0.00492052f $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_92 N_A_79_21#_c_79_n N_A_243_47#_c_225_n 0.00112065f $X=2.77 $Y=0.785 $X2=0
+ $Y2=0
cc_93 N_A_79_21#_c_77_n N_A_243_47#_c_226_n 0.0107783f $X=2.49 $Y=1.895 $X2=0
+ $Y2=0
cc_94 N_A_79_21#_c_79_n N_A_243_47#_c_226_n 0.00306755f $X=2.77 $Y=0.785 $X2=0
+ $Y2=0
cc_95 N_A_79_21#_c_78_n N_A_243_47#_c_227_n 0.00183297f $X=2.77 $Y=0.445 $X2=0
+ $Y2=0
cc_96 N_A_79_21#_c_79_n N_A_243_47#_c_227_n 0.0113123f $X=2.77 $Y=0.785 $X2=0
+ $Y2=0
cc_97 N_A_79_21#_c_84_n N_A_243_47#_c_232_n 0.0101096f $X=2.13 $Y=2.285 $X2=0
+ $Y2=0
cc_98 N_A_79_21#_c_77_n N_A_243_47#_c_232_n 0.0138681f $X=2.49 $Y=1.895 $X2=0
+ $Y2=0
cc_99 N_A_79_21#_c_87_n N_A_243_47#_c_232_n 0.00705702f $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_100 N_A_79_21#_c_77_n N_A_243_47#_c_229_n 0.0487793f $X=2.49 $Y=1.895 $X2=0
+ $Y2=0
cc_101 N_A_79_21#_c_79_n N_A_243_47#_c_229_n 0.00353808f $X=2.77 $Y=0.785 $X2=0
+ $Y2=0
cc_102 N_A_79_21#_c_82_n N_A_243_47#_c_234_n 0.0051555f $X=1.155 $Y=1.89 $X2=0
+ $Y2=0
cc_103 N_A_79_21#_c_84_n N_A_243_47#_c_234_n 0.00805606f $X=2.13 $Y=2.285 $X2=0
+ $Y2=0
cc_104 N_A_79_21#_c_77_n N_A_243_47#_c_234_n 0.00611524f $X=2.49 $Y=1.895 $X2=0
+ $Y2=0
cc_105 N_A_79_21#_c_87_n N_A_243_47#_c_234_n 5.78476e-19 $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_106 N_A_79_21#_c_77_n N_B2_M1001_g 0.00174754f $X=2.49 $Y=1.895 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_78_n N_B2_M1001_g 0.00111676f $X=2.77 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_79_n N_B2_M1001_g 0.00325332f $X=2.77 $Y=0.785 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_77_n N_B2_c_293_n 0.00115391f $X=2.49 $Y=1.895 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_77_n B2 0.0307643f $X=2.49 $Y=1.895 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_79_n B1 0.00406739f $X=2.77 $Y=0.785 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_74_n X 0.0197919f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_75_n X 0.0134543f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_76_n X 0.0594311f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_129_p X 0.013769f $X=0.685 $Y=1.89 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_76_n N_VPWR_M1003_d 0.00390096f $X=0.6 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_117 N_A_79_21#_c_82_n N_VPWR_M1003_d 0.0118658f $X=1.155 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_118 N_A_79_21#_c_129_p N_VPWR_M1003_d 5.4783e-19 $X=0.685 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_79_21#_c_75_n N_VPWR_c_375_n 0.0125971f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_82_n N_VPWR_c_375_n 0.0113742f $X=1.155 $Y=1.89 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_129_p N_VPWR_c_375_n 0.00622534f $X=0.685 $Y=1.89 $X2=0
+ $Y2=0
cc_122 N_A_79_21#_c_85_n N_VPWR_c_375_n 0.00896244f $X=1.375 $Y=2.285 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_c_82_n N_VPWR_c_377_n 0.00356258f $X=1.155 $Y=1.89 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_84_n N_VPWR_c_377_n 0.0304585f $X=2.13 $Y=2.285 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_85_n N_VPWR_c_377_n 0.00969682f $X=1.375 $Y=2.285 $X2=0
+ $Y2=0
cc_126 N_A_79_21#_c_87_n N_VPWR_c_377_n 0.0215386f $X=2.3 $Y=2.275 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_75_n N_VPWR_c_379_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_79_21#_M1000_s N_VPWR_c_374_n 0.00241861f $X=2.175 $Y=2.065 $X2=0
+ $Y2=0
cc_129 N_A_79_21#_c_75_n N_VPWR_c_374_n 0.00835414f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_82_n N_VPWR_c_374_n 0.00758377f $X=1.155 $Y=1.89 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_129_p N_VPWR_c_374_n 8.39522e-19 $X=0.685 $Y=1.89 $X2=0
+ $Y2=0
cc_132 N_A_79_21#_c_84_n N_VPWR_c_374_n 0.0264428f $X=2.13 $Y=2.285 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_85_n N_VPWR_c_374_n 0.00800038f $X=1.375 $Y=2.285 $X2=0
+ $Y2=0
cc_134 N_A_79_21#_c_87_n N_VPWR_c_374_n 0.0153548f $X=2.3 $Y=2.275 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_82_n A_241_297# 0.00405998f $X=1.155 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_136 N_A_79_21#_c_87_n N_A_525_413#_c_432_n 0.0124315f $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_137 N_A_79_21#_c_77_n N_A_525_413#_c_434_n 0.00474796f $X=2.49 $Y=1.895 $X2=0
+ $Y2=0
cc_138 N_A_79_21#_c_87_n N_A_525_413#_c_434_n 0.00930488f $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_139 N_A_79_21#_c_87_n N_A_525_413#_c_439_n 0.0111686f $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_140 N_A_79_21#_c_74_n N_VGND_c_473_n 0.00468308f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_78_n N_VGND_c_474_n 0.0110645f $X=2.77 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_79_n N_VGND_c_474_n 0.00446391f $X=2.77 $Y=0.785 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_74_n N_VGND_c_475_n 0.0103325f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_75_n N_VGND_c_475_n 0.00231239f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_76_n N_VGND_c_475_n 0.0053584f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_79_n N_VGND_c_477_n 6.41288e-19 $X=2.77 $Y=0.785 $X2=0 $Y2=0
cc_147 N_A_79_21#_M1002_d N_VGND_c_478_n 0.00413042f $X=2.635 $Y=0.235 $X2=0
+ $Y2=0
cc_148 N_A_79_21#_c_74_n N_VGND_c_478_n 0.00895861f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_78_n N_VGND_c_478_n 0.00640047f $X=2.77 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_79_21#_c_79_n N_VGND_c_478_n 0.00729903f $X=2.77 $Y=0.785 $X2=0 $Y2=0
cc_151 N_A1_N_c_165_n N_A2_N_c_195_n 0.054623f $X=1.115 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_152 A1_N N_A2_N_c_195_n 0.00741123f $X=1.105 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_153 N_A1_N_M1008_g N_A2_N_M1006_g 0.0240691f $X=1.14 $Y=0.445 $X2=0 $Y2=0
cc_154 N_A1_N_c_165_n A2_N 3.56086e-19 $X=1.115 $Y=1.41 $X2=0 $Y2=0
cc_155 A1_N A2_N 0.0296811f $X=1.105 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A1_N_M1008_g N_A_243_47#_c_228_n 0.00536216f $X=1.14 $Y=0.445 $X2=0
+ $Y2=0
cc_157 A1_N N_A_243_47#_c_228_n 0.00541889f $X=1.105 $Y=1.105 $X2=0 $Y2=0
cc_158 A1_N N_A_243_47#_c_234_n 0.00308021f $X=1.105 $Y=1.105 $X2=0 $Y2=0
cc_159 A1_N N_VPWR_M1003_d 0.00168449f $X=1.105 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_160 N_A1_N_c_165_n N_VPWR_c_377_n 0.00241764f $X=1.115 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A1_N_c_165_n N_VPWR_c_374_n 0.00363302f $X=1.115 $Y=1.41 $X2=0 $Y2=0
cc_162 A1_N A_241_297# 0.00226506f $X=1.105 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_163 N_A1_N_c_165_n N_VGND_c_475_n 3.19739e-19 $X=1.115 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A1_N_M1008_g N_VGND_c_475_n 0.00548195f $X=1.14 $Y=0.445 $X2=0 $Y2=0
cc_165 A1_N N_VGND_c_475_n 0.00188799f $X=1.105 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A1_N_M1008_g N_VGND_c_476_n 0.00585385f $X=1.14 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A1_N_M1008_g N_VGND_c_478_n 0.0113114f $X=1.14 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A2_N_c_195_n N_A_243_47#_c_223_n 5.38281e-19 $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_169 N_A2_N_c_195_n N_A_243_47#_c_225_n 0.0127581f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A2_N_M1006_g N_A_243_47#_c_225_n 0.00521083f $X=1.56 $Y=0.445 $X2=0
+ $Y2=0
cc_171 A2_N N_A_243_47#_c_225_n 0.00196206f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_172 N_A2_N_c_195_n N_A_243_47#_c_227_n 0.00363831f $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_173 N_A2_N_M1006_g N_A_243_47#_c_227_n 0.0136001f $X=1.56 $Y=0.445 $X2=0
+ $Y2=0
cc_174 A2_N N_A_243_47#_c_227_n 0.0173932f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_175 N_A2_N_c_195_n N_A_243_47#_c_229_n 0.00503897f $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A2_N_M1006_g N_A_243_47#_c_229_n 0.00175871f $X=1.56 $Y=0.445 $X2=0
+ $Y2=0
cc_177 A2_N N_A_243_47#_c_229_n 0.0182487f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_178 A2_N N_A_243_47#_c_234_n 0.00325851f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_179 N_A2_N_M1006_g N_VGND_c_476_n 0.00428022f $X=1.56 $Y=0.445 $X2=0 $Y2=0
cc_180 N_A2_N_M1006_g N_VGND_c_477_n 0.00834626f $X=1.56 $Y=0.445 $X2=0 $Y2=0
cc_181 N_A2_N_M1006_g N_VGND_c_478_n 0.00716774f $X=1.56 $Y=0.445 $X2=0 $Y2=0
cc_182 N_A_243_47#_M1002_g N_B2_M1001_g 0.0173449f $X=2.56 $Y=0.445 $X2=0 $Y2=0
cc_183 N_A_243_47#_c_223_n N_B2_c_293_n 0.0173449f $X=2.535 $Y=1.89 $X2=0 $Y2=0
cc_184 N_A_243_47#_c_231_n N_B2_c_294_n 0.0296932f $X=2.535 $Y=1.99 $X2=0 $Y2=0
cc_185 N_A_243_47#_c_226_n B2 0.00403862f $X=2.535 $Y=1.065 $X2=0 $Y2=0
cc_186 N_A_243_47#_c_226_n N_B2_c_292_n 0.0173449f $X=2.535 $Y=1.065 $X2=0 $Y2=0
cc_187 N_A_243_47#_c_231_n N_VPWR_c_377_n 0.00513788f $X=2.535 $Y=1.99 $X2=0
+ $Y2=0
cc_188 N_A_243_47#_c_231_n N_VPWR_c_374_n 0.00828969f $X=2.535 $Y=1.99 $X2=0
+ $Y2=0
cc_189 N_A_243_47#_c_231_n N_A_525_413#_c_432_n 0.00156703f $X=2.535 $Y=1.99
+ $X2=0 $Y2=0
cc_190 N_A_243_47#_c_223_n N_A_525_413#_c_434_n 0.00107876f $X=2.535 $Y=1.89
+ $X2=0 $Y2=0
cc_191 N_A_243_47#_c_231_n N_A_525_413#_c_439_n 0.0031145f $X=2.535 $Y=1.99
+ $X2=0 $Y2=0
cc_192 N_A_243_47#_c_227_n N_VGND_M1006_d 0.00182057f $X=2.04 $Y=0.74 $X2=0
+ $Y2=0
cc_193 N_A_243_47#_M1002_g N_VGND_c_474_n 0.00434414f $X=2.56 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_A_243_47#_c_281_p N_VGND_c_476_n 0.0112554f $X=1.35 $Y=0.445 $X2=0
+ $Y2=0
cc_195 N_A_243_47#_c_227_n N_VGND_c_476_n 0.00381617f $X=2.04 $Y=0.74 $X2=0
+ $Y2=0
cc_196 N_A_243_47#_M1002_g N_VGND_c_477_n 0.0108036f $X=2.56 $Y=0.445 $X2=0
+ $Y2=0
cc_197 N_A_243_47#_c_225_n N_VGND_c_477_n 0.00697993f $X=2.435 $Y=1.065 $X2=0
+ $Y2=0
cc_198 N_A_243_47#_c_227_n N_VGND_c_477_n 0.0420473f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_243_47#_M1008_d N_VGND_c_478_n 0.00412745f $X=1.215 $Y=0.235 $X2=0
+ $Y2=0
cc_200 N_A_243_47#_M1002_g N_VGND_c_478_n 0.00742902f $X=2.56 $Y=0.445 $X2=0
+ $Y2=0
cc_201 N_A_243_47#_c_281_p N_VGND_c_478_n 0.00644035f $X=1.35 $Y=0.445 $X2=0
+ $Y2=0
cc_202 N_A_243_47#_c_227_n N_VGND_c_478_n 0.00819503f $X=2.04 $Y=0.74 $X2=0
+ $Y2=0
cc_203 N_B2_M1001_g N_B1_M1007_g 0.0432259f $X=2.98 $Y=0.445 $X2=0 $Y2=0
cc_204 N_B2_c_293_n N_B1_c_333_n 0.0086983f $X=3.005 $Y=1.89 $X2=0 $Y2=0
cc_205 N_B2_c_294_n N_B1_c_334_n 0.0205581f $X=3.005 $Y=1.99 $X2=0 $Y2=0
cc_206 N_B2_M1001_g B1 0.00493429f $X=2.98 $Y=0.445 $X2=0 $Y2=0
cc_207 B2 B1 0.0412625f $X=2.985 $Y=1.445 $X2=0 $Y2=0
cc_208 N_B2_c_292_n B1 0.00186087f $X=3.04 $Y=1.47 $X2=0 $Y2=0
cc_209 B2 N_B1_c_332_n 0.00131497f $X=2.985 $Y=1.445 $X2=0 $Y2=0
cc_210 N_B2_c_292_n N_B1_c_332_n 0.0203097f $X=3.04 $Y=1.47 $X2=0 $Y2=0
cc_211 N_B2_c_294_n N_VPWR_c_376_n 0.00499876f $X=3.005 $Y=1.99 $X2=0 $Y2=0
cc_212 N_B2_c_294_n N_VPWR_c_377_n 0.00513173f $X=3.005 $Y=1.99 $X2=0 $Y2=0
cc_213 N_B2_c_294_n N_VPWR_c_374_n 0.00679831f $X=3.005 $Y=1.99 $X2=0 $Y2=0
cc_214 N_B2_c_294_n N_A_525_413#_c_432_n 0.00526001f $X=3.005 $Y=1.99 $X2=0
+ $Y2=0
cc_215 N_B2_c_293_n N_A_525_413#_c_433_n 0.0036561f $X=3.005 $Y=1.89 $X2=0 $Y2=0
cc_216 N_B2_c_294_n N_A_525_413#_c_433_n 0.00689197f $X=3.005 $Y=1.99 $X2=0
+ $Y2=0
cc_217 B2 N_A_525_413#_c_433_n 0.0154584f $X=2.985 $Y=1.445 $X2=0 $Y2=0
cc_218 N_B2_c_292_n N_A_525_413#_c_433_n 0.0010573f $X=3.04 $Y=1.47 $X2=0 $Y2=0
cc_219 N_B2_c_293_n N_A_525_413#_c_434_n 0.00113449f $X=3.005 $Y=1.89 $X2=0
+ $Y2=0
cc_220 N_B2_c_294_n N_A_525_413#_c_434_n 0.00138352f $X=3.005 $Y=1.99 $X2=0
+ $Y2=0
cc_221 B2 N_A_525_413#_c_434_n 0.00393971f $X=2.985 $Y=1.445 $X2=0 $Y2=0
cc_222 N_B2_c_294_n N_A_525_413#_c_439_n 0.00244193f $X=3.005 $Y=1.99 $X2=0
+ $Y2=0
cc_223 N_B2_M1001_g N_VGND_c_472_n 0.00220228f $X=2.98 $Y=0.445 $X2=0 $Y2=0
cc_224 N_B2_M1001_g N_VGND_c_474_n 0.00585385f $X=2.98 $Y=0.445 $X2=0 $Y2=0
cc_225 N_B2_M1001_g N_VGND_c_478_n 0.0110141f $X=2.98 $Y=0.445 $X2=0 $Y2=0
cc_226 N_B1_c_334_n N_VPWR_c_376_n 0.00900356f $X=3.485 $Y=1.99 $X2=0 $Y2=0
cc_227 N_B1_c_334_n N_VPWR_c_380_n 0.00468263f $X=3.485 $Y=1.99 $X2=0 $Y2=0
cc_228 N_B1_c_334_n N_VPWR_c_374_n 0.00646284f $X=3.485 $Y=1.99 $X2=0 $Y2=0
cc_229 N_B1_c_334_n N_A_525_413#_c_432_n 7.38983e-19 $X=3.485 $Y=1.99 $X2=0
+ $Y2=0
cc_230 N_B1_c_333_n N_A_525_413#_c_433_n 0.00543479f $X=3.485 $Y=1.89 $X2=0
+ $Y2=0
cc_231 N_B1_c_334_n N_A_525_413#_c_433_n 0.0101339f $X=3.485 $Y=1.99 $X2=0 $Y2=0
cc_232 B1 N_A_525_413#_c_433_n 0.0192526f $X=3.455 $Y=0.765 $X2=0 $Y2=0
cc_233 N_B1_c_332_n N_A_525_413#_c_433_n 0.00102541f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_234 N_B1_c_334_n N_A_525_413#_c_435_n 0.00585773f $X=3.485 $Y=1.99 $X2=0
+ $Y2=0
cc_235 N_B1_M1007_g N_VGND_c_472_n 0.0146687f $X=3.46 $Y=0.445 $X2=0 $Y2=0
cc_236 B1 N_VGND_c_472_n 0.00891566f $X=3.455 $Y=0.765 $X2=0 $Y2=0
cc_237 N_B1_c_332_n N_VGND_c_472_n 0.00137613f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_238 N_B1_M1007_g N_VGND_c_474_n 0.00407992f $X=3.46 $Y=0.445 $X2=0 $Y2=0
cc_239 N_B1_M1007_g N_VGND_c_478_n 0.00395858f $X=3.46 $Y=0.445 $X2=0 $Y2=0
cc_240 B1 N_VGND_c_478_n 0.00492962f $X=3.455 $Y=0.765 $X2=0 $Y2=0
cc_241 X N_VPWR_c_375_n 0.0177194f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_242 X N_VPWR_c_379_n 0.0182101f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_243 N_X_M1003_s N_VPWR_c_374_n 0.00430086f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_244 X N_VPWR_c_374_n 0.00993603f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_245 X N_VGND_c_473_n 0.018001f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_246 N_X_M1011_s N_VGND_c_478_n 0.00387172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_247 X N_VGND_c_478_n 0.00993603f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_248 N_VPWR_c_374_n N_A_525_413#_M1000_d 0.00233855f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_249 N_VPWR_c_374_n N_A_525_413#_M1005_d 0.00354071f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_376_n N_A_525_413#_c_432_n 0.00493711f $X=3.24 $Y=2.34 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_376_n N_A_525_413#_c_433_n 0.0177704f $X=3.24 $Y=2.34 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_377_n N_A_525_413#_c_433_n 0.00297063f $X=3.155 $Y=2.72 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_380_n N_A_525_413#_c_433_n 0.00310557f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_374_n N_A_525_413#_c_433_n 0.0109181f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_376_n N_A_525_413#_c_435_n 0.0173145f $X=3.24 $Y=2.34 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_380_n N_A_525_413#_c_435_n 0.0124472f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_374_n N_A_525_413#_c_435_n 0.00684138f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_376_n N_A_525_413#_c_439_n 0.0109524f $X=3.24 $Y=2.34 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_377_n N_A_525_413#_c_439_n 0.0145661f $X=3.155 $Y=2.72 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_374_n N_A_525_413#_c_439_n 0.0119869f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_261 N_VGND_c_478_n A_611_47# 0.013552f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
