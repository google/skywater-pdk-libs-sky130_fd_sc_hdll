* File: sky130_fd_sc_hdll__dfrtp_4.pex.spice
* Created: Thu Aug 27 19:04:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%CLK 1 2 3 5 6 8 13 14
c37 3 0 9.59708e-20 $X=0.495 $Y=1.74
c38 1 0 2.71124e-20 $X=0.305 $Y=1.325
r39 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=1.16
+ $X2=0.265 $Y2=1.53
r40 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r41 6 18 86.21 $w=2.7e-07 $l=5.0709e-07 $layer=POLY_cond $X=0.52 $Y=0.73
+ $X2=0.352 $Y2=1.16
r42 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r43 3 9 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.305 $Y2=1.665
r44 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r45 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r46 1 18 38.9026 $w=2.7e-07 $l=1.87029e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.352 $Y2=1.16
r47 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.305 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%A_27_47# 1 2 8 9 11 14 17 20 22 23 25 26
+ 28 29 30 31 33 36 40 44 45 46 49 52 53 54 55 58 64 72 75 76 81
c245 81 0 4.78096e-20 $X=6.57 $Y=1.11
c246 64 0 1.76704e-20 $X=6.61 $Y=1.19
c247 54 0 1.58851e-19 $X=6.465 $Y=1.19
c248 30 0 7.17362e-20 $X=6.32 $Y=1.89
c249 23 0 1.85946e-19 $X=2.92 $Y=1.32
r250 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.57
+ $Y=1.11 $X2=6.57 $Y2=1.11
r251 75 78 37.1829 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=0.93
+ $X2=2.76 $Y2=1.095
r252 75 77 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=0.93
+ $X2=2.76 $Y2=0.765
r253 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.735
+ $Y=0.93 $X2=2.735 $Y2=0.93
r254 71 72 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r255 68 71 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=0.805 $Y=1.235
+ $X2=0.965 $Y2=1.235
r256 64 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.61 $Y=1.19
+ $X2=6.61 $Y2=1.19
r257 62 76 7.49088 $w=3.98e-07 $l=2.6e-07 $layer=LI1_cond $X=2.735 $Y=1.19
+ $X2=2.735 $Y2=0.93
r258 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.68 $Y=1.19
+ $X2=2.68 $Y2=1.19
r259 58 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.805
+ $Y=1.235 $X2=0.805 $Y2=1.235
r260 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.745 $Y=1.19
+ $X2=0.745 $Y2=1.19
r261 55 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.825 $Y=1.19
+ $X2=2.68 $Y2=1.19
r262 54 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.465 $Y=1.19
+ $X2=6.61 $Y2=1.19
r263 54 55 4.50494 $w=1.4e-07 $l=3.64e-06 $layer=MET1_cond $X=6.465 $Y=1.19
+ $X2=2.825 $Y2=1.19
r264 53 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.89 $Y=1.19
+ $X2=0.745 $Y2=1.19
r265 52 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.535 $Y=1.19
+ $X2=2.68 $Y2=1.19
r266 52 53 2.03589 $w=1.4e-07 $l=1.645e-06 $layer=MET1_cond $X=2.535 $Y=1.19
+ $X2=0.89 $Y2=1.19
r267 51 58 30.3143 $w=2.28e-07 $l=6.05e-07 $layer=LI1_cond $X=0.775 $Y=1.795
+ $X2=0.775 $Y2=1.19
r268 50 58 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.775 $Y=0.805
+ $X2=0.775 $Y2=1.19
r269 47 49 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.217 $Y2=1.88
r270 46 51 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.775 $Y2=1.795
r271 46 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.345 $Y2=1.88
r272 44 50 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.775 $Y2=0.805
r273 44 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.345 $Y2=0.72
r274 38 45 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.345 $Y2=0.72
r275 38 40 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.217 $Y2=0.51
r276 34 80 38.8967 $w=3.59e-07 $l=1.76125e-07 $layer=POLY_cond $X=6.51 $Y=0.945
+ $X2=6.487 $Y2=1.11
r277 34 36 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.51 $Y=0.945
+ $X2=6.51 $Y2=0.415
r278 31 33 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.32 $Y=1.99
+ $X2=6.32 $Y2=2.275
r279 30 31 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.32 $Y=1.89 $X2=6.32
+ $Y2=1.99
r280 29 80 47.6452 $w=3.59e-07 $l=3.58915e-07 $layer=POLY_cond $X=6.32 $Y=1.395
+ $X2=6.487 $Y2=1.11
r281 29 30 164.131 $w=2e-07 $l=4.95e-07 $layer=POLY_cond $X=6.32 $Y=1.395
+ $X2=6.32 $Y2=1.89
r282 26 28 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.405 $Y=1.99
+ $X2=3.405 $Y2=2.275
r283 25 26 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.405 $Y=1.89 $X2=3.405
+ $Y2=1.99
r284 24 25 164.131 $w=2e-07 $l=4.95e-07 $layer=POLY_cond $X=3.405 $Y=1.395
+ $X2=3.405 $Y2=1.89
r285 22 24 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=3.305 $Y=1.32
+ $X2=3.405 $Y2=1.395
r286 22 23 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.305 $Y=1.32
+ $X2=2.92 $Y2=1.32
r287 20 77 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.84 $Y=0.415
+ $X2=2.84 $Y2=0.765
r288 17 23 27.7801 $w=1.5e-07 $l=1.35403e-07 $layer=POLY_cond $X=2.817 $Y=1.245
+ $X2=2.92 $Y2=1.32
r289 17 78 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=2.817 $Y=1.245
+ $X2=2.817 $Y2=1.095
r290 12 72 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r291 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r292 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r293 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r294 7 71 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r295 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r296 2 49 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r297 1 40 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%D 3 6 7 9 10 11 16 20
c56 11 0 1.94832e-19 $X=2.19 $Y=1.3
c57 6 0 1.76402e-19 $X=2.35 $Y=1.89
r58 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.89
+ $Y=1.465 $X2=1.89 $Y2=1.465
r59 16 20 1.4951 $w=5.18e-07 $l=6.5e-08 $layer=LI1_cond $X=1.715 $Y=1.53
+ $X2=1.715 $Y2=1.465
r60 10 19 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.19 $Y=1.465 $X2=1.89
+ $Y2=1.465
r61 10 11 3.18546 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.465
+ $X2=2.19 $Y2=1.3
r62 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.35 $Y=1.99 $X2=2.35
+ $Y2=2.275
r63 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.35 $Y=1.89 $X2=2.35
+ $Y2=1.99
r64 5 11 33.332 $w=1.75e-07 $l=4.02119e-07 $layer=POLY_cond $X=2.35 $Y=1.63
+ $X2=2.19 $Y2=1.3
r65 5 6 86.2101 $w=2e-07 $l=2.6e-07 $layer=POLY_cond $X=2.35 $Y=1.63 $X2=2.35
+ $Y2=1.89
r66 1 11 33.332 $w=1.75e-07 $l=7.5e-08 $layer=POLY_cond $X=2.265 $Y=1.3 $X2=2.19
+ $Y2=1.3
r67 1 3 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.265 $Y=1.3
+ $X2=2.265 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%A_211_363# 1 2 7 9 12 14 16 17 19 21 24 25
+ 27 28 32 35 36 37 38 45 47 55 63 65
c210 63 0 3.94709e-20 $X=6.815 $Y=1.74
c211 55 0 1.61046e-19 $X=3.37 $Y=0.9
c212 45 0 1.76402e-19 $X=3.19 $Y=1.87
c213 36 0 9.59708e-20 $X=1.345 $Y=1.87
c214 35 0 1.17518e-19 $X=3.045 $Y=1.87
c215 27 0 1.76704e-20 $X=6.47 $Y=1.58
c216 24 0 1.25508e-19 $X=6.04 $Y=0.87
r217 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.815
+ $Y=1.74 $X2=6.815 $Y2=1.74
r218 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.74 $X2=2.845 $Y2=1.74
r219 48 63 3.59637 $w=4.41e-07 $l=1.3e-07 $layer=LI1_cond $X=6.75 $Y=1.87
+ $X2=6.75 $Y2=1.74
r220 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.61 $Y=1.87
+ $X2=6.61 $Y2=1.87
r221 45 52 10.1947 $w=3.88e-07 $l=3.45e-07 $layer=LI1_cond $X=3.19 $Y=1.77
+ $X2=2.845 $Y2=1.77
r222 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.19 $Y=1.87
+ $X2=3.19 $Y2=1.87
r223 41 65 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.2 $Y=1.87
+ $X2=1.2 $Y2=0.51
r224 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.87 $X2=1.2
+ $Y2=1.87
r225 38 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.335 $Y=1.87
+ $X2=3.19 $Y2=1.87
r226 37 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.465 $Y=1.87
+ $X2=6.61 $Y2=1.87
r227 37 38 3.87375 $w=1.4e-07 $l=3.13e-06 $layer=MET1_cond $X=6.465 $Y=1.87
+ $X2=3.335 $Y2=1.87
r228 36 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.87
+ $X2=1.2 $Y2=1.87
r229 35 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.045 $Y=1.87
+ $X2=3.19 $Y2=1.87
r230 35 36 2.10396 $w=1.4e-07 $l=1.7e-06 $layer=MET1_cond $X=3.045 $Y=1.87
+ $X2=1.345 $Y2=1.87
r231 33 55 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.295 $Y=0.9
+ $X2=3.37 $Y2=0.9
r232 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=0.9 $X2=3.295 $Y2=0.9
r233 29 32 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=3.19 $Y=0.875
+ $X2=3.295 $Y2=0.875
r234 27 63 4.4263 $w=4.41e-07 $l=3.50999e-07 $layer=LI1_cond $X=6.47 $Y=1.58
+ $X2=6.75 $Y2=1.74
r235 27 28 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.47 $Y=1.58
+ $X2=6.125 $Y2=1.58
r236 25 57 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=6.04 $Y=0.87
+ $X2=5.865 $Y2=0.87
r237 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.04
+ $Y=0.87 $X2=6.04 $Y2=0.87
r238 22 28 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.02 $Y=1.495
+ $X2=6.125 $Y2=1.58
r239 22 24 33.0087 $w=2.08e-07 $l=6.25e-07 $layer=LI1_cond $X=6.02 $Y=1.495
+ $X2=6.02 $Y2=0.87
r240 21 45 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.19 $Y=1.575
+ $X2=3.19 $Y2=1.77
r241 20 29 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.19 $Y=0.985
+ $X2=3.19 $Y2=0.875
r242 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.19 $Y=0.985
+ $X2=3.19 $Y2=1.575
r243 17 62 48.1208 $w=2.95e-07 $l=2.54951e-07 $layer=POLY_cond $X=6.85 $Y=1.99
+ $X2=6.84 $Y2=1.74
r244 17 19 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.85 $Y=1.99
+ $X2=6.85 $Y2=2.275
r245 14 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.865 $Y=0.705
+ $X2=5.865 $Y2=0.87
r246 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.865 $Y=0.705
+ $X2=5.865 $Y2=0.415
r247 10 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.37 $Y=0.765
+ $X2=3.37 $Y2=0.9
r248 10 12 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.37 $Y=0.765
+ $X2=3.37 $Y2=0.415
r249 7 51 46.5577 $w=3.26e-07 $l=2.54951e-07 $layer=POLY_cond $X=2.86 $Y=1.99
+ $X2=2.87 $Y2=1.74
r250 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.86 $Y=1.99
+ $X2=2.86 $Y2=2.275
r251 2 41 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r252 1 65 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%A_811_289# 1 2 7 9 12 14 20 22 24 25 26 29
+ 32 35 36
c106 36 0 2.93959e-20 $X=5.59 $Y=1.61
c107 35 0 1.0473e-19 $X=5.52 $Y=0.835
c108 22 0 4.23403e-20 $X=5.59 $Y=1.525
r109 32 34 3.06272 $w=3.98e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0.36
+ $X2=5.565 $Y2=0.445
r110 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.03 $Y=2.005
+ $X2=6.03 $Y2=2.3
r111 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.945 $Y=1.92
+ $X2=6.03 $Y2=2.005
r112 25 26 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.945 $Y=1.92
+ $X2=5.675 $Y2=1.92
r113 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.59 $Y=1.835
+ $X2=5.675 $Y2=1.92
r114 23 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.59 $Y=1.695
+ $X2=5.59 $Y2=1.61
r115 23 24 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.59 $Y=1.695
+ $X2=5.59 $Y2=1.835
r116 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.59 $Y=1.525
+ $X2=5.59 $Y2=1.61
r117 22 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.59 $Y=1.525
+ $X2=5.59 $Y2=0.835
r118 20 35 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=5.52 $Y=0.68
+ $X2=5.52 $Y2=0.835
r119 20 34 8.73626 $w=3.08e-07 $l=2.35e-07 $layer=LI1_cond $X=5.52 $Y=0.68
+ $X2=5.52 $Y2=0.445
r120 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.19
+ $Y=1.61 $X2=4.19 $Y2=1.61
r121 14 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=1.61
+ $X2=5.59 $Y2=1.61
r122 14 16 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=5.505 $Y=1.61
+ $X2=4.19 $Y2=1.61
r123 10 17 38.8084 $w=2.75e-07 $l=1.80748e-07 $layer=POLY_cond $X=4.25 $Y=1.445
+ $X2=4.217 $Y2=1.61
r124 10 12 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.25 $Y=1.445
+ $X2=4.25 $Y2=0.445
r125 7 17 72.3531 $w=2.75e-07 $l=4.09829e-07 $layer=POLY_cond $X=4.155 $Y=1.99
+ $X2=4.217 $Y2=1.61
r126 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.155 $Y=1.99
+ $X2=4.155 $Y2=2.275
r127 2 29 600 $w=1.7e-07 $l=7.32871e-07 $layer=licon1_PDIFF $count=1 $X=5.865
+ $Y=1.645 $X2=6.03 $Y2=2.3
r128 1 32 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.445
+ $Y=0.235 $X2=5.6 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%RESET_B 3 5 6 8 10 11 13 16 18 23 24 25 28
+ 29 30 33 42 49 54
c154 29 0 6.20412e-20 $X=4.67 $Y=0.93
c155 28 0 1.0473e-19 $X=4.67 $Y=0.93
r156 46 49 9.96707 $w=3.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.955 $Y=1.22
+ $X2=8.275 $Y2=1.22
r157 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.955 $Y=1.165
+ $X2=7.955 $Y2=1.165
r158 43 54 0.0466954 $w=5.22e-07 $l=1.95e-07 $layer=MET1_cond $X=8.25 $Y=1.007
+ $X2=8.055 $Y2=1.007
r159 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.25 $Y=0.85
+ $X2=8.25 $Y2=0.85
r160 40 49 3.2703 $w=2.4e-07 $l=1.85e-07 $layer=LI1_cond $X=8.275 $Y=1.035
+ $X2=8.275 $Y2=1.22
r161 40 42 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=8.275 $Y=1.035
+ $X2=8.275 $Y2=0.85
r162 33 36 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.995 $Y=1.12
+ $X2=7.995 $Y2=1.285
r163 33 35 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.995 $Y=1.12
+ $X2=7.995 $Y2=0.955
r164 33 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.97
+ $Y=1.12 $X2=7.97 $Y2=1.12
r165 28 31 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.695 $Y=0.93
+ $X2=4.695 $Y2=1.095
r166 28 30 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.695 $Y=0.93
+ $X2=4.695 $Y2=0.765
r167 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.67
+ $Y=0.93 $X2=4.67 $Y2=0.93
r168 25 54 0.00119732 $w=5.22e-07 $l=5e-09 $layer=MET1_cond $X=8.05 $Y=1.007
+ $X2=8.055 $Y2=1.007
r169 25 47 0.022749 $w=5.22e-07 $l=9.5e-08 $layer=MET1_cond $X=8.05 $Y=1.007
+ $X2=7.955 $Y2=1.007
r170 23 47 0.11063 $w=5.22e-07 $l=2.17748e-07 $layer=MET1_cond $X=7.81 $Y=0.85
+ $X2=7.955 $Y2=1.007
r171 23 24 3.57054 $w=1.4e-07 $l=2.885e-06 $layer=MET1_cond $X=7.81 $Y=0.85
+ $X2=4.925 $Y2=0.85
r172 20 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.73 $Y=0.85
+ $X2=4.73 $Y2=0.85
r173 18 24 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=4.81 $Y=0.85
+ $X2=4.925 $Y2=0.85
r174 18 20 0.0513283 $w=2.3e-07 $l=8e-08 $layer=MET1_cond $X=4.81 $Y=0.85
+ $X2=4.73 $Y2=0.85
r175 16 35 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.985 $Y=0.445
+ $X2=7.985 $Y2=0.955
r176 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.96 $Y=1.99
+ $X2=7.96 $Y2=2.275
r177 10 11 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.96 $Y=1.89 $X2=7.96
+ $Y2=1.99
r178 10 36 200.604 $w=2e-07 $l=6.05e-07 $layer=POLY_cond $X=7.96 $Y=1.89
+ $X2=7.96 $Y2=1.285
r179 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.69 $Y=1.99
+ $X2=4.69 $Y2=2.275
r180 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.69 $Y=1.89 $X2=4.69
+ $Y2=1.99
r181 5 31 263.604 $w=2e-07 $l=7.95e-07 $layer=POLY_cond $X=4.69 $Y=1.89 $X2=4.69
+ $Y2=1.095
r182 3 30 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.61 $Y=0.445
+ $X2=4.61 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%A_583_47# 1 2 9 11 13 15 16 20 25 27 28 29
+ 34 35
c128 35 0 6.20412e-20 $X=5.2 $Y=1.17
c129 29 0 1.61046e-19 $X=3.85 $Y=1.27
c130 9 0 1.25508e-19 $X=5.37 $Y=0.555
r131 35 40 51.3607 $w=3.05e-07 $l=3.25e-07 $layer=POLY_cond $X=5.255 $Y=1.17
+ $X2=5.255 $Y2=1.495
r132 34 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.2 $Y=1.17 $X2=5.2
+ $Y2=1.27
r133 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.2
+ $Y=1.17 $X2=5.2 $Y2=1.17
r134 30 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.58 $Y=1.27
+ $X2=3.765 $Y2=1.27
r135 29 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=1.27
+ $X2=3.765 $Y2=1.27
r136 28 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=1.27
+ $X2=5.2 $Y2=1.27
r137 28 29 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=5.115 $Y=1.27
+ $X2=3.85 $Y2=1.27
r138 27 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=1.185
+ $X2=3.765 $Y2=1.27
r139 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.765 $Y=0.475
+ $X2=3.765 $Y2=1.185
r140 24 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=1.355
+ $X2=3.58 $Y2=1.27
r141 24 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.58 $Y=1.355
+ $X2=3.58 $Y2=2.135
r142 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.68 $Y=0.39
+ $X2=3.765 $Y2=0.475
r143 20 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.68 $Y=0.39
+ $X2=3.11 $Y2=0.39
r144 16 25 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.495 $Y=2.3
+ $X2=3.58 $Y2=2.135
r145 16 18 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.495 $Y=2.3
+ $X2=3.1 $Y2=2.3
r146 13 15 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=5.775 $Y=1.57
+ $X2=5.775 $Y2=2.065
r147 12 40 19.3576 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.445 $Y=1.495
+ $X2=5.255 $Y2=1.495
r148 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.685 $Y=1.495
+ $X2=5.775 $Y2=1.57
r149 11 12 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.685 $Y=1.495
+ $X2=5.445 $Y2=1.495
r150 7 35 38.5368 $w=3.05e-07 $l=2.14942e-07 $layer=POLY_cond $X=5.37 $Y=1.005
+ $X2=5.255 $Y2=1.17
r151 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.37 $Y=1.005
+ $X2=5.37 $Y2=0.555
r152 2 18 600 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=2.95
+ $Y=2.065 $X2=3.1 $Y2=2.33
r153 1 22 182 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.11 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%A_1403_21# 1 2 9 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 42 46 47 48 51 53 54 55 56 57 58 64 69 75 85
c199 75 0 6.23215e-20 $X=7.37 $Y=0.98
c200 69 0 2.04429e-20 $X=7.85 $Y=0.78
c201 57 0 1.99375e-19 $X=8.875 $Y=1.295
c202 12 0 2.4959e-20 $X=7.37 $Y=1.89
r203 85 86 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=10.865 $Y=1.202
+ $X2=10.89 $Y2=1.202
r204 82 83 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=10.395 $Y=1.202
+ $X2=10.42 $Y2=1.202
r205 81 82 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=9.95 $Y=1.202
+ $X2=10.395 $Y2=1.202
r206 80 81 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=9.925 $Y=1.202
+ $X2=9.95 $Y2=1.202
r207 79 80 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=9.48 $Y=1.202
+ $X2=9.925 $Y2=1.202
r208 65 85 30.6135 $w=3.7e-07 $l=2.35e-07 $layer=POLY_cond $X=10.63 $Y=1.202
+ $X2=10.865 $Y2=1.202
r209 65 83 27.3568 $w=3.7e-07 $l=2.1e-07 $layer=POLY_cond $X=10.63 $Y=1.202
+ $X2=10.42 $Y2=1.202
r210 64 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.63
+ $Y=1.16 $X2=10.63 $Y2=1.16
r211 62 79 2.60541 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=9.46 $Y=1.202
+ $X2=9.48 $Y2=1.202
r212 62 77 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=9.46 $Y=1.202
+ $X2=9.455 $Y2=1.202
r213 61 64 61.7922 $w=2.08e-07 $l=1.17e-06 $layer=LI1_cond $X=9.46 $Y=1.18
+ $X2=10.63 $Y2=1.18
r214 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.46
+ $Y=1.16 $X2=9.46 $Y2=1.16
r215 59 73 3.45218 $w=2.1e-07 $l=1.73e-07 $layer=LI1_cond $X=8.96 $Y=1.18
+ $X2=8.787 $Y2=1.18
r216 59 61 26.4069 $w=2.08e-07 $l=5e-07 $layer=LI1_cond $X=8.96 $Y=1.18 $X2=9.46
+ $Y2=1.18
r217 57 73 7.13508 $w=3.34e-07 $l=1.52791e-07 $layer=LI1_cond $X=8.875 $Y=1.295
+ $X2=8.787 $Y2=1.18
r218 57 58 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.875 $Y=1.295
+ $X2=8.875 $Y2=1.915
r219 56 73 13.1497 $w=3.34e-07 $l=3.65951e-07 $layer=LI1_cond $X=8.775 $Y=0.82
+ $X2=8.787 $Y2=1.18
r220 55 72 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.775 $Y=0.465
+ $X2=8.775 $Y2=0.38
r221 55 56 12.7849 $w=3.18e-07 $l=3.55e-07 $layer=LI1_cond $X=8.775 $Y=0.465
+ $X2=8.775 $Y2=0.82
r222 53 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.79 $Y=2
+ $X2=8.875 $Y2=1.915
r223 53 54 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.79 $Y=2 $X2=8.28
+ $Y2=2
r224 49 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.195 $Y=2.085
+ $X2=8.28 $Y2=2
r225 49 51 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.195 $Y=2.085
+ $X2=8.195 $Y2=2.21
r226 47 72 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.615 $Y=0.38
+ $X2=8.775 $Y2=0.38
r227 47 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.615 $Y=0.38
+ $X2=7.935 $Y2=0.38
r228 46 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.85 $Y=0.695
+ $X2=7.85 $Y2=0.78
r229 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.85 $Y=0.465
+ $X2=7.935 $Y2=0.38
r230 45 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.85 $Y=0.465
+ $X2=7.85 $Y2=0.695
r231 43 75 13.2835 $w=2.54e-07 $l=7e-08 $layer=POLY_cond $X=7.44 $Y=0.98
+ $X2=7.37 $Y2=0.98
r232 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.44
+ $Y=0.98 $X2=7.44 $Y2=0.98
r233 40 69 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.49 $Y=0.78
+ $X2=7.85 $Y2=0.78
r234 40 42 4.90855 $w=2.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.49 $Y=0.865
+ $X2=7.49 $Y2=0.98
r235 37 86 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.89 $Y=0.995
+ $X2=10.89 $Y2=1.202
r236 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.89 $Y=0.995
+ $X2=10.89 $Y2=0.56
r237 34 85 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.865 $Y=1.41
+ $X2=10.865 $Y2=1.202
r238 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.865 $Y=1.41
+ $X2=10.865 $Y2=1.985
r239 31 83 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.42 $Y=0.995
+ $X2=10.42 $Y2=1.202
r240 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.42 $Y=0.995
+ $X2=10.42 $Y2=0.56
r241 28 82 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.395 $Y=1.41
+ $X2=10.395 $Y2=1.202
r242 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.395 $Y=1.41
+ $X2=10.395 $Y2=1.985
r243 25 81 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.95 $Y=0.995
+ $X2=9.95 $Y2=1.202
r244 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.95 $Y=0.995
+ $X2=9.95 $Y2=0.56
r245 22 80 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.925 $Y=1.41
+ $X2=9.925 $Y2=1.202
r246 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.925 $Y=1.41
+ $X2=9.925 $Y2=1.985
r247 19 79 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.48 $Y=0.995
+ $X2=9.48 $Y2=1.202
r248 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.48 $Y=0.995
+ $X2=9.48 $Y2=0.56
r249 16 77 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.455 $Y=1.41
+ $X2=9.455 $Y2=1.202
r250 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.455 $Y=1.41
+ $X2=9.455 $Y2=1.985
r251 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.37 $Y=1.99
+ $X2=7.37 $Y2=2.275
r252 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.37 $Y=1.89 $X2=7.37
+ $Y2=1.99
r253 11 75 8.45288 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.37 $Y=1.145
+ $X2=7.37 $Y2=0.98
r254 11 12 247.025 $w=2e-07 $l=7.45e-07 $layer=POLY_cond $X=7.37 $Y=1.145
+ $X2=7.37 $Y2=1.89
r255 7 75 53.1339 $w=2.54e-07 $l=3.52987e-07 $layer=POLY_cond $X=7.09 $Y=0.815
+ $X2=7.37 $Y2=0.98
r256 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.09 $Y=0.815
+ $X2=7.09 $Y2=0.445
r257 2 51 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=8.05
+ $Y=2.065 $X2=8.195 $Y2=2.21
r258 1 72 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=8.565
+ $Y=0.235 $X2=8.7 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%A_1188_47# 1 2 7 9 12 14 18 23 25 26 28
c100 26 0 2.04429e-20 $X=7.47 $Y=1.66
c101 23 0 1.92806e-19 $X=7.05 $Y=1.315
r102 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.405
+ $Y=1.66 $X2=8.405 $Y2=1.66
r103 26 28 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=7.47 $Y=1.66 $X2=8.405
+ $Y2=1.66
r104 24 26 6.67215 $w=2.83e-07 $l=1.30576e-07 $layer=LI1_cond $X=7.36 $Y=1.615
+ $X2=7.47 $Y2=1.66
r105 24 25 19.9058 $w=2.18e-07 $l=3.8e-07 $layer=LI1_cond $X=7.36 $Y=1.745
+ $X2=7.36 $Y2=2.125
r106 23 24 13.364 $w=2.83e-07 $l=4.34856e-07 $layer=LI1_cond $X=7.05 $Y=1.315
+ $X2=7.36 $Y2=1.615
r107 22 23 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=7.05 $Y=0.535
+ $X2=7.05 $Y2=1.315
r108 18 25 7.23167 $w=3.4e-07 $l=2.18174e-07 $layer=LI1_cond $X=7.25 $Y=2.295
+ $X2=7.36 $Y2=2.125
r109 18 20 23.2183 $w=3.38e-07 $l=6.85e-07 $layer=LI1_cond $X=7.25 $Y=2.295
+ $X2=6.565 $Y2=2.295
r110 14 22 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.965 $Y=0.395
+ $X2=7.05 $Y2=0.535
r111 14 16 31.4864 $w=2.78e-07 $l=7.65e-07 $layer=LI1_cond $X=6.965 $Y=0.395
+ $X2=6.2 $Y2=0.395
r112 10 29 38.7299 $w=2.8e-07 $l=1.92678e-07 $layer=POLY_cond $X=8.49 $Y=1.495
+ $X2=8.43 $Y2=1.66
r113 10 12 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=8.49 $Y=1.495
+ $X2=8.49 $Y2=0.445
r114 7 29 62.9382 $w=2.8e-07 $l=3.3e-07 $layer=POLY_cond $X=8.43 $Y=1.99
+ $X2=8.43 $Y2=1.66
r115 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=8.43 $Y=1.99
+ $X2=8.43 $Y2=2.275
r116 2 20 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=6.41
+ $Y=2.065 $X2=6.565 $Y2=2.335
r117 1 16 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=5.94
+ $Y=0.235 $X2=6.2 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 48
+ 52 56 60 63 64 65 66 68 69 71 72 74 75 76 78 83 88 114 115 118 121 124 127
r171 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r172 127 130 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=8.65 $Y=2.34
+ $X2=8.65 $Y2=2.72
r173 124 125 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r174 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r175 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r176 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r177 112 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r178 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r179 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r180 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r181 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r182 106 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r183 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r184 103 130 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.84 $Y=2.72
+ $X2=8.65 $Y2=2.72
r185 103 105 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=8.84 $Y=2.72
+ $X2=8.97 $Y2=2.72
r186 102 131 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r187 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r188 99 102 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=7.59 $Y2=2.72
r189 98 101 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=7.59 $Y2=2.72
r190 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r191 96 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r192 96 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r193 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r194 93 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=4.455 $Y2=2.72
r195 93 95 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=5.29 $Y2=2.72
r196 92 125 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.37 $Y2=2.72
r197 92 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r198 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r199 89 121 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.2 $Y=2.72
+ $X2=2.075 $Y2=2.72
r200 89 91 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.2 $Y=2.72
+ $X2=2.53 $Y2=2.72
r201 88 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.29 $Y=2.72
+ $X2=4.455 $Y2=2.72
r202 88 91 114.824 $w=1.68e-07 $l=1.76e-06 $layer=LI1_cond $X=4.29 $Y=2.72
+ $X2=2.53 $Y2=2.72
r203 87 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r204 87 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r205 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r206 84 118 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r207 84 86 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r208 83 121 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.95 $Y=2.72
+ $X2=2.075 $Y2=2.72
r209 83 86 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.95 $Y=2.72
+ $X2=1.61 $Y2=2.72
r210 78 118 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r211 78 80 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r212 76 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r213 76 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r214 74 111 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=11.015 $Y=2.72
+ $X2=10.81 $Y2=2.72
r215 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.015 $Y=2.72
+ $X2=11.1 $Y2=2.72
r216 73 114 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=11.185 $Y=2.72
+ $X2=11.27 $Y2=2.72
r217 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.185 $Y=2.72
+ $X2=11.1 $Y2=2.72
r218 71 108 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=10.075 $Y=2.72
+ $X2=9.89 $Y2=2.72
r219 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.075 $Y=2.72
+ $X2=10.16 $Y2=2.72
r220 70 111 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=10.245 $Y=2.72
+ $X2=10.81 $Y2=2.72
r221 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.245 $Y=2.72
+ $X2=10.16 $Y2=2.72
r222 68 105 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.135 $Y=2.72
+ $X2=8.97 $Y2=2.72
r223 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.135 $Y=2.72
+ $X2=9.22 $Y2=2.72
r224 67 108 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=9.305 $Y=2.72
+ $X2=9.89 $Y2=2.72
r225 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.305 $Y=2.72
+ $X2=9.22 $Y2=2.72
r226 65 101 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=7.64 $Y=2.72
+ $X2=7.59 $Y2=2.72
r227 65 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.64 $Y=2.72
+ $X2=7.765 $Y2=2.72
r228 63 95 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.305 $Y=2.72
+ $X2=5.29 $Y2=2.72
r229 63 64 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.305 $Y=2.72
+ $X2=5.515 $Y2=2.72
r230 62 98 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.725 $Y=2.72
+ $X2=5.75 $Y2=2.72
r231 62 64 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.725 $Y=2.72
+ $X2=5.515 $Y2=2.72
r232 58 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.1 $Y=2.635
+ $X2=11.1 $Y2=2.72
r233 58 60 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=11.1 $Y=2.635
+ $X2=11.1 $Y2=1.96
r234 54 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.16 $Y=2.635
+ $X2=10.16 $Y2=2.72
r235 54 56 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=10.16 $Y=2.635
+ $X2=10.16 $Y2=1.96
r236 50 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.22 $Y=2.635
+ $X2=9.22 $Y2=2.72
r237 50 52 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.22 $Y=2.635
+ $X2=9.22 $Y2=2
r238 49 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.89 $Y=2.72
+ $X2=7.765 $Y2=2.72
r239 48 130 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.46 $Y=2.72
+ $X2=8.65 $Y2=2.72
r240 48 49 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.46 $Y=2.72
+ $X2=7.89 $Y2=2.72
r241 44 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.765 $Y=2.635
+ $X2=7.765 $Y2=2.72
r242 44 46 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.765 $Y=2.635
+ $X2=7.765 $Y2=2.34
r243 40 64 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.515 $Y=2.635
+ $X2=5.515 $Y2=2.72
r244 40 42 8.09454 $w=4.18e-07 $l=2.95e-07 $layer=LI1_cond $X=5.515 $Y=2.635
+ $X2=5.515 $Y2=2.34
r245 36 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=2.635
+ $X2=4.455 $Y2=2.72
r246 36 38 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.455 $Y=2.635
+ $X2=4.455 $Y2=2.29
r247 32 121 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=2.635
+ $X2=2.075 $Y2=2.72
r248 32 34 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.075 $Y=2.635
+ $X2=2.075 $Y2=2.34
r249 28 118 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r250 28 30 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r251 9 60 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.955
+ $Y=1.485 $X2=11.1 $Y2=1.96
r252 8 56 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.015
+ $Y=1.485 $X2=10.16 $Y2=1.96
r253 7 52 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=9.095
+ $Y=1.485 $X2=9.22 $Y2=2
r254 6 127 600 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=8.52
+ $Y=2.065 $X2=8.675 $Y2=2.34
r255 5 46 600 $w=1.7e-07 $l=3.85357e-07 $layer=licon1_PDIFF $count=1 $X=7.46
+ $Y=2.065 $X2=7.725 $Y2=2.34
r256 4 42 600 $w=1.7e-07 $l=7.77592e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.645 $X2=5.54 $Y2=2.34
r257 3 38 600 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=2.065 $X2=4.455 $Y2=2.29
r258 2 34 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=2.065 $X2=2.115 $Y2=2.34
r259 1 30 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%A_468_47# 1 2 8 9 11
c35 8 0 6.84282e-20 $X=2.23 $Y=1.835
r36 9 11 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.315 $Y=0.39
+ $X2=2.525 $Y2=0.39
r37 8 14 21.8265 $w=2.86e-07 $l=5.51883e-07 $layer=LI1_cond $X=2.23 $Y=1.835
+ $X2=2.42 $Y2=2.3
r38 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.23 $Y=0.475
+ $X2=2.315 $Y2=0.39
r39 7 8 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.23 $Y=0.475
+ $X2=2.23 $Y2=1.835
r40 2 14 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=2.065 $X2=2.585 $Y2=2.3
r41 1 11 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.34
+ $Y=0.235 $X2=2.525 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%A_699_413# 1 2 9 11 12 15
c37 12 0 1.58851e-19 $X=4.005 $Y=1.95
r38 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.925 $Y=2.035
+ $X2=4.925 $Y2=2.21
r39 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.84 $Y=1.95
+ $X2=4.925 $Y2=2.035
r40 11 12 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.84 $Y=1.95
+ $X2=4.005 $Y2=1.95
r41 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=2.035
+ $X2=4.005 $Y2=1.95
r42 7 9 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.92 $Y=2.035
+ $X2=3.92 $Y2=2.21
r43 2 15 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.78
+ $Y=2.065 $X2=4.925 $Y2=2.21
r44 1 9 600 $w=1.7e-07 $l=4.92189e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=2.065 $X2=3.92 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%Q 1 2 3 4 15 17 19 21 22 23 27 31 33 35 39
+ 41 42 43 44 50 51
r77 44 51 2.47908 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=11.2 $Y=1.54 $X2=11.2
+ $Y2=1.455
r78 44 51 0.140542 $w=4.08e-07 $l=5e-09 $layer=LI1_cond $X=11.2 $Y=1.45 $X2=11.2
+ $Y2=1.455
r79 43 44 7.30818 $w=4.08e-07 $l=2.6e-07 $layer=LI1_cond $X=11.2 $Y=1.19
+ $X2=11.2 $Y2=1.45
r80 42 50 2.47908 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=11.2 $Y=0.82 $X2=11.2
+ $Y2=0.905
r81 42 43 7.58926 $w=4.08e-07 $l=2.7e-07 $layer=LI1_cond $X=11.2 $Y=0.92
+ $X2=11.2 $Y2=1.19
r82 42 50 0.421625 $w=4.08e-07 $l=1.5e-08 $layer=LI1_cond $X=11.2 $Y=0.92
+ $X2=11.2 $Y2=0.905
r83 36 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.795 $Y=0.82
+ $X2=10.605 $Y2=0.82
r84 35 42 5.97895 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=10.995 $Y=0.82
+ $X2=11.2 $Y2=0.82
r85 35 36 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=10.995 $Y=0.82
+ $X2=10.795 $Y2=0.82
r86 34 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.755 $Y=1.54
+ $X2=10.63 $Y2=1.54
r87 33 44 5.97895 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=10.995 $Y=1.54
+ $X2=11.2 $Y2=1.54
r88 33 34 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.995 $Y=1.54
+ $X2=10.755 $Y2=1.54
r89 29 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.63 $Y=1.625
+ $X2=10.63 $Y2=1.54
r90 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=10.63 $Y=1.625
+ $X2=10.63 $Y2=2.3
r91 25 39 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.605 $Y=0.735
+ $X2=10.605 $Y2=0.82
r92 25 27 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=10.605 $Y=0.735
+ $X2=10.605 $Y2=0.39
r93 24 38 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.855 $Y=1.54
+ $X2=9.71 $Y2=1.54
r94 23 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.505 $Y=1.54
+ $X2=10.63 $Y2=1.54
r95 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=10.505 $Y=1.54
+ $X2=9.855 $Y2=1.54
r96 21 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.415 $Y=0.82
+ $X2=10.605 $Y2=0.82
r97 21 22 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=10.415 $Y=0.82
+ $X2=9.855 $Y2=0.82
r98 17 38 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.71 $Y=1.625
+ $X2=9.71 $Y2=1.54
r99 17 19 26.8241 $w=2.88e-07 $l=6.75e-07 $layer=LI1_cond $X=9.71 $Y=1.625
+ $X2=9.71 $Y2=2.3
r100 13 22 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=9.665 $Y=0.735
+ $X2=9.855 $Y2=0.82
r101 13 15 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=9.665 $Y=0.735
+ $X2=9.665 $Y2=0.39
r102 4 41 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.485
+ $Y=1.485 $X2=10.63 $Y2=1.62
r103 4 31 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=10.485
+ $Y=1.485 $X2=10.63 $Y2=2.3
r104 3 38 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.545
+ $Y=1.485 $X2=9.69 $Y2=1.62
r105 3 19 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.545
+ $Y=1.485 $X2=9.69 $Y2=2.3
r106 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=10.495
+ $Y=0.235 $X2=10.63 $Y2=0.39
r107 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.555
+ $Y=0.235 $X2=9.69 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFRTP_4%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 47 48
+ 50 51 53 54 56 57 58 60 69 73 92 93 97 103 106
c169 93 0 2.26487e-19 $X=11.27 $Y=0
r170 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r171 103 104 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r172 97 100 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r173 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r174 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r175 90 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r176 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r177 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r178 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r179 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r180 84 107 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=7.59 $Y2=0
r181 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r182 81 106 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.475 $Y2=0
r183 81 83 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=8.97 $Y2=0
r184 80 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r185 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r186 77 80 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=7.13 $Y2=0
r187 77 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.83 $Y2=0
r188 76 79 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=5.29 $Y=0 $X2=7.13
+ $Y2=0
r189 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r190 74 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=4.99 $Y2=0
r191 74 76 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=5.29 $Y2=0
r192 73 106 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.355 $Y=0
+ $X2=7.475 $Y2=0
r193 73 79 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.355 $Y=0
+ $X2=7.13 $Y2=0
r194 72 104 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=4.83 $Y2=0
r195 71 72 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r196 69 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=4.99 $Y2=0
r197 69 71 179.738 $w=1.68e-07 $l=2.755e-06 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=2.07 $Y2=0
r198 68 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r199 68 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r200 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r201 65 97 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r202 65 67 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.61 $Y2=0
r203 60 97 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r204 60 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r205 58 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r206 58 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r207 56 89 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=11.015 $Y=0
+ $X2=10.81 $Y2=0
r208 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.015 $Y=0 $X2=11.1
+ $Y2=0
r209 55 92 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=11.185 $Y=0
+ $X2=11.27 $Y2=0
r210 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.185 $Y=0 $X2=11.1
+ $Y2=0
r211 53 86 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=10.075 $Y=0
+ $X2=9.89 $Y2=0
r212 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.075 $Y=0
+ $X2=10.16 $Y2=0
r213 52 89 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=10.245 $Y=0
+ $X2=10.81 $Y2=0
r214 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.245 $Y=0
+ $X2=10.16 $Y2=0
r215 50 83 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.135 $Y=0
+ $X2=8.97 $Y2=0
r216 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.135 $Y=0 $X2=9.22
+ $Y2=0
r217 49 86 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=9.305 $Y=0
+ $X2=9.89 $Y2=0
r218 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.305 $Y=0 $X2=9.22
+ $Y2=0
r219 47 67 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.645 $Y=0 $X2=1.61
+ $Y2=0
r220 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=0 $X2=1.81
+ $Y2=0
r221 46 71 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.07
+ $Y2=0
r222 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.81
+ $Y2=0
r223 42 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.1 $Y=0.085
+ $X2=11.1 $Y2=0
r224 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.1 $Y=0.085
+ $X2=11.1 $Y2=0.39
r225 38 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.16 $Y=0.085
+ $X2=10.16 $Y2=0
r226 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.16 $Y=0.085
+ $X2=10.16 $Y2=0.39
r227 34 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.22 $Y=0.085
+ $X2=9.22 $Y2=0
r228 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.22 $Y=0.085
+ $X2=9.22 $Y2=0.39
r229 30 106 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.475 $Y=0.085
+ $X2=7.475 $Y2=0
r230 30 32 13.2051 $w=2.38e-07 $l=2.75e-07 $layer=LI1_cond $X=7.475 $Y=0.085
+ $X2=7.475 $Y2=0.36
r231 26 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0
r232 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0.38
r233 22 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0
r234 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0.36
r235 7 44 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=10.965
+ $Y=0.235 $X2=11.1 $Y2=0.39
r236 6 40 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=10.025
+ $Y=0.235 $X2=10.16 $Y2=0.39
r237 5 36 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=9.095
+ $Y=0.235 $X2=9.22 $Y2=0.39
r238 4 32 182 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_NDIFF $count=1 $X=7.165
+ $Y=0.235 $X2=7.46 $Y2=0.36
r239 3 28 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.235 $X2=4.99 $Y2=0.38
r240 2 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.665
+ $Y=0.235 $X2=1.81 $Y2=0.36
r241 1 100 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

