* File: sky130_fd_sc_hdll__nor3b_2.pex.spice
* Created: Thu Aug 27 19:16:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR3B_2%A 1 3 4 6 7 9 10 12 13 14 22 27
c37 14 0 1.93357e-19 $X=0.66 $Y=1.105
r38 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.01 $Y2=1.202
r39 20 22 43.1263 $w=3.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.645 $Y=1.202
+ $X2=0.985 $Y2=1.202
r40 20 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r41 18 20 16.4895 $w=3.8e-07 $l=1.3e-07 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.645 $Y2=1.202
r42 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r43 14 27 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=0.745 $Y=1.18
+ $X2=0.645 $Y2=1.18
r44 13 27 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.645 $Y2=1.18
r45 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.202
r46 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r47 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r48 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r49 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r50 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r51 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_2%B 1 3 4 6 7 9 10 12 13 20 23
c42 20 0 1.93357e-19 $X=1.925 $Y=1.202
r43 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r44 18 20 31.7105 $w=3.8e-07 $l=2.5e-07 $layer=POLY_cond $X=1.675 $Y=1.202
+ $X2=1.925 $Y2=1.202
r45 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.675
+ $Y=1.16 $X2=1.675 $Y2=1.16
r46 16 18 27.9053 $w=3.8e-07 $l=2.2e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.675 $Y2=1.202
r47 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r48 13 23 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=1.765 $Y=1.18
+ $X2=1.615 $Y2=1.18
r49 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r50 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r51 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r52 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r53 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r54 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r55 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995 $X2=1.43
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_2%A_571_21# 1 2 7 9 10 12 13 15 16 18 19 25
+ 29 32 34 35 40
r62 39 40 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=3.4 $Y=1.202
+ $X2=3.425 $Y2=1.202
r63 38 39 58.9258 $w=3.64e-07 $l=4.45e-07 $layer=POLY_cond $X=2.955 $Y=1.202
+ $X2=3.4 $Y2=1.202
r64 37 38 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=2.93 $Y=1.202
+ $X2=2.955 $Y2=1.202
r65 34 35 11.2584 $w=3.53e-07 $l=2.5e-07 $layer=LI1_cond $X=4.167 $Y=1.705
+ $X2=4.167 $Y2=1.455
r66 29 31 11.0961 $w=3.53e-07 $l=2.45e-07 $layer=LI1_cond $X=4.167 $Y=0.66
+ $X2=4.167 $Y2=0.905
r67 26 32 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.075 $Y=1.285
+ $X2=4.075 $Y2=1.18
r68 26 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.075 $Y=1.285
+ $X2=4.075 $Y2=1.455
r69 25 32 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.075 $Y=1.075
+ $X2=4.075 $Y2=1.18
r70 25 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.075 $Y=1.075
+ $X2=4.075 $Y2=0.905
r71 22 40 36.4148 $w=3.64e-07 $l=2.75e-07 $layer=POLY_cond $X=3.7 $Y=1.202
+ $X2=3.425 $Y2=1.202
r72 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.7
+ $Y=1.16 $X2=3.7 $Y2=1.16
r73 19 32 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.18
+ $X2=4.075 $Y2=1.18
r74 19 21 15.316 $w=2.08e-07 $l=2.9e-07 $layer=LI1_cond $X=3.99 $Y=1.18 $X2=3.7
+ $Y2=1.18
r75 16 40 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.425 $Y2=1.202
r76 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.425 $Y2=1.985
r77 13 39 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.4 $Y=0.995 $X2=3.4
+ $Y2=1.202
r78 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.4 $Y=0.995 $X2=3.4
+ $Y2=0.56
r79 10 38 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.202
r80 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.985
r81 7 37 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=1.202
r82 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.93 $Y=0.995 $X2=2.93
+ $Y2=0.56
r83 2 34 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=4.095
+ $Y=1.485 $X2=4.22 $Y2=1.705
r84 1 29 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.465 $X2=4.22 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_2%C_N 1 3 4 6 7 15
r25 11 15 8.45022 $w=2.08e-07 $l=1.6e-07 $layer=LI1_cond $X=4.495 $Y=1.18
+ $X2=4.655 $Y2=1.18
r26 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.495
+ $Y=1.16 $X2=4.495 $Y2=1.16
r27 7 15 3.4329 $w=2.08e-07 $l=6.5e-08 $layer=LI1_cond $X=4.72 $Y=1.18 $X2=4.655
+ $Y2=1.18
r28 4 10 47.8775 $w=2.99e-07 $l=2.79285e-07 $layer=POLY_cond $X=4.455 $Y=1.41
+ $X2=4.517 $Y2=1.16
r29 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.455 $Y=1.41
+ $X2=4.455 $Y2=1.695
r30 1 10 38.5562 $w=2.99e-07 $l=2.03912e-07 $layer=POLY_cond $X=4.43 $Y=0.995
+ $X2=4.517 $Y2=1.16
r31 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.43 $Y=0.995 $X2=4.43
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_2%A_27_297# 1 2 3 10 12 14 18 20 27 29
r40 21 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=1.54
+ $X2=1.22 $Y2=1.54
r41 20 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=1.54
+ $X2=2.16 $Y2=1.54
r42 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.995 $Y=1.54
+ $X2=1.345 $Y2=1.54
r43 16 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=1.54
r44 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=2.3
r45 15 25 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.247 $Y2=1.54
r46 14 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=1.22 $Y2=1.54
r47 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=0.405 $Y2=1.54
r48 10 25 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=1.625
+ $X2=0.247 $Y2=1.54
r49 10 12 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=0.247 $Y=1.625
+ $X2=0.247 $Y2=2.3
r50 3 29 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.61
r51 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r52 2 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r53 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r54 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_2%VPWR 1 2 11 13 15 17 19 28 32
r45 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r46 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r48 25 26 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r49 23 26 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=4.37 $Y2=2.72
r50 23 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 22 25 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=4.37 $Y2=2.72
r52 22 23 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 20 28 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r54 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 19 31 3.88626 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.812 $Y2=2.72
r56 19 25 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.37 $Y2=2.72
r57 17 29 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r58 13 31 3.2569 $w=2.5e-07 $l=1.58915e-07 $layer=LI1_cond $X=4.69 $Y=2.635
+ $X2=4.812 $Y2=2.72
r59 13 15 42.8709 $w=2.48e-07 $l=9.3e-07 $layer=LI1_cond $X=4.69 $Y=2.635
+ $X2=4.69 $Y2=1.705
r60 9 28 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r61 9 11 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r62 2 15 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=4.545
+ $Y=1.485 $X2=4.69 $Y2=1.705
r63 1 11 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_2%A_309_297# 1 2 3 12 14 15 18 20
r27 18 23 3.04665 $w=2.45e-07 $l=9.5e-08 $layer=LI1_cond $X=3.657 $Y=2.275
+ $X2=3.657 $Y2=2.37
r28 18 20 30.8102 $w=2.43e-07 $l=6.55e-07 $layer=LI1_cond $X=3.657 $Y=2.275
+ $X2=3.657 $Y2=1.62
r29 15 17 52.8278 $w=1.88e-07 $l=9.05e-07 $layer=LI1_cond $X=1.815 $Y=2.37
+ $X2=2.72 $Y2=2.37
r30 14 23 3.91254 $w=1.9e-07 $l=1.22e-07 $layer=LI1_cond $X=3.535 $Y=2.37
+ $X2=3.657 $Y2=2.37
r31 14 17 47.5742 $w=1.88e-07 $l=8.15e-07 $layer=LI1_cond $X=3.535 $Y=2.37
+ $X2=2.72 $Y2=2.37
r32 10 15 6.98266 $w=1.9e-07 $l=1.65831e-07 $layer=LI1_cond $X=1.69 $Y=2.275
+ $X2=1.815 $Y2=2.37
r33 10 12 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=1.69 $Y=2.275
+ $X2=1.69 $Y2=1.96
r34 3 23 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.485 $X2=3.66 $Y2=2.3
r35 3 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.485 $X2=3.66 $Y2=1.62
r36 2 17 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=1.485 $X2=2.72 $Y2=2.36
r37 1 12 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_2%Y 1 2 3 4 15 17 18 21 23 27 29 31 32 35
r68 32 35 3.29269 $w=4.18e-07 $l=1.2e-07 $layer=LI1_cond $X=3.145 $Y=0.51
+ $X2=3.145 $Y2=0.39
r69 30 32 5.89941 $w=4.18e-07 $l=2.15e-07 $layer=LI1_cond $X=3.145 $Y=0.725
+ $X2=3.145 $Y2=0.51
r70 30 31 2.27389 $w=4.52e-07 $l=1.05214e-07 $layer=LI1_cond $X=3.145 $Y=0.725
+ $X2=3.112 $Y2=0.815
r71 25 31 2.27389 $w=4.52e-07 $l=9e-08 $layer=LI1_cond $X=3.112 $Y=0.905
+ $X2=3.112 $Y2=0.815
r72 25 27 17.6329 $w=4.83e-07 $l=7.15e-07 $layer=LI1_cond $X=3.112 $Y=0.905
+ $X2=3.112 $Y2=1.62
r73 24 29 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=0.815
+ $X2=1.665 $Y2=0.815
r74 23 31 4.79675 $w=1.8e-07 $l=2.42e-07 $layer=LI1_cond $X=2.87 $Y=0.815
+ $X2=3.112 $Y2=0.815
r75 23 24 62.5404 $w=1.78e-07 $l=1.015e-06 $layer=LI1_cond $X=2.87 $Y=0.815
+ $X2=1.855 $Y2=0.815
r76 19 29 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.815
r77 19 21 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.39
r78 17 29 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=1.665 $Y2=0.815
r79 17 18 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=0.915 $Y2=0.815
r80 13 18 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.815
r81 13 15 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r82 4 27 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.045
+ $Y=1.485 $X2=3.19 $Y2=1.62
r83 3 35 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.005
+ $Y=0.235 $X2=3.19 $Y2=0.39
r84 2 21 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r85 1 15 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_2%VGND 1 2 3 4 5 6 19 21 23 27 31 33 35 38
+ 39 40 51 59 63 69 72
r72 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r73 68 69 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=0.235
+ $X2=2.765 $Y2=0.235
r74 65 68 2.80331 $w=6.38e-07 $l=1.5e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.68 $Y2=0.235
r75 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r76 62 65 6.91483 $w=6.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=0.235
+ $X2=2.53 $Y2=0.235
r77 62 63 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.235
+ $X2=2.075 $Y2=0.235
r78 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r79 54 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r80 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r81 51 71 4.23306 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=4.565 $Y=0 $X2=4.812
+ $Y2=0
r82 51 53 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.565 $Y=0 $X2=4.37
+ $Y2=0
r83 50 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r84 50 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r85 49 69 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=2.765
+ $Y2=0
r86 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r87 46 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r88 46 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r89 45 63 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.075
+ $Y2=0
r90 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r91 43 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r92 43 45 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=2.07
+ $Y2=0
r93 40 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r94 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r95 38 49 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=0 $X2=3.45
+ $Y2=0
r96 38 39 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=3.575 $Y=0 $X2=3.677
+ $Y2=0
r97 37 53 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=4.37
+ $Y2=0
r98 37 39 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=3.677
+ $Y2=0
r99 33 71 3.20479 $w=2.9e-07 $l=1.38109e-07 $layer=LI1_cond $X=4.71 $Y=0.085
+ $X2=4.812 $Y2=0
r100 33 35 22.8502 $w=2.88e-07 $l=5.75e-07 $layer=LI1_cond $X=4.71 $Y=0.085
+ $X2=4.71 $Y2=0.66
r101 29 39 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.677 $Y=0.085
+ $X2=3.677 $Y2=0
r102 29 31 16.5011 $w=2.03e-07 $l=3.05e-07 $layer=LI1_cond $X=3.677 $Y=0.085
+ $X2=3.677 $Y2=0.39
r103 25 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r104 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r105 24 56 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r106 23 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r107 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=0.365 $Y2=0
r108 19 56 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r109 19 21 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r110 6 35 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=4.505
+ $Y=0.465 $X2=4.69 $Y2=0.66
r111 5 31 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.475
+ $Y=0.235 $X2=3.66 $Y2=0.39
r112 4 68 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.235 $X2=2.68 $Y2=0.39
r113 3 62 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r114 2 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
r115 1 21 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

