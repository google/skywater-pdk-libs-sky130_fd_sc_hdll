* File: sky130_fd_sc_hdll__o221a_2.spice
* Created: Wed Sep  2 08:44:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o221a_2.pex.spice"
.subckt sky130_fd_sc_hdll__o221a_2  VNB VPB C1 B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1002 N_A_151_47#_M1002_d N_C1_M1002_g N_A_38_47#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.26975 PD=0.97 PS=2.13 NRD=0 NRS=23.988 M=1 R=4.33333
+ SA=75000.3 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1001 N_A_245_47#_M1001_d N_B1_M1001_g N_A_151_47#_M1002_d VNB NSHORT L=0.15
+ W=0.65 AD=0.092625 AS=0.104 PD=0.935 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.8 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1003 N_A_151_47#_M1003_d N_B2_M1003_g N_A_245_47#_M1001_d VNB NSHORT L=0.15
+ W=0.65 AD=0.19175 AS=0.092625 PD=1.89 PS=0.935 NRD=5.532 NRS=1.836 M=1
+ R=4.33333 SA=75001.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_245_47#_M1008_d N_A2_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_245_47#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1004_d N_A_38_47#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_38_47#_M1013_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_C1_M1007_g N_A_38_47#_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.335 PD=1.35 PS=2.67 NRD=7.8603 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1000 A_255_297# N_B1_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=1 AD=0.1225
+ AS=0.175 PD=1.245 PS=1.35 NRD=13.2778 NRS=5.8903 M=1 R=5.55556 SA=90000.8
+ SB=90003 A=0.18 P=2.36 MULT=1
MM1010 N_A_38_47#_M1010_d N_B2_M1010_g A_255_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.3975 AS=0.1225 PD=1.795 PS=1.245 NRD=0.9653 NRS=13.2778 M=1 R=5.55556
+ SA=90001.2 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1006 A_535_297# N_A2_M1006_g N_A_38_47#_M1010_d VPB PHIGHVT L=0.18 W=1
+ AD=0.115 AS=0.3975 PD=1.23 PS=1.795 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90002.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g A_535_297# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.115 PD=1.35 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90002.6
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1005_d N_A_38_47#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.145 PD=1.35 PS=1.29 NRD=12.7853 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_38_47#_M1012_g N_X_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX15_noxref noxref_16 A2 A2 PROBETYPE=1
pX16_noxref noxref_17 A2 A2 PROBETYPE=1
pX17_noxref noxref_18 A1 A1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o221a_2.pxi.spice"
*
.ends
*
*
