* File: sky130_fd_sc_hdll__o21ai_1.pxi.spice
* Created: Wed Sep  2 08:43:24 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21AI_1%A1 N_A1_c_36_n N_A1_M1002_g N_A1_c_37_n
+ N_A1_M1005_g A1 N_A1_c_38_n PM_SKY130_FD_SC_HDLL__O21AI_1%A1
x_PM_SKY130_FD_SC_HDLL__O21AI_1%A2 N_A2_c_58_n N_A2_M1001_g N_A2_c_59_n
+ N_A2_M1004_g A2 A2 A2 A2 N_A2_c_60_n PM_SKY130_FD_SC_HDLL__O21AI_1%A2
x_PM_SKY130_FD_SC_HDLL__O21AI_1%B1 N_B1_M1003_g N_B1_c_98_n N_B1_M1000_g B1
+ N_B1_c_97_n PM_SKY130_FD_SC_HDLL__O21AI_1%B1
x_PM_SKY130_FD_SC_HDLL__O21AI_1%VPWR N_VPWR_M1002_s N_VPWR_M1000_d
+ N_VPWR_c_126_n N_VPWR_c_127_n N_VPWR_c_128_n N_VPWR_c_129_n VPWR
+ N_VPWR_c_130_n N_VPWR_c_125_n PM_SKY130_FD_SC_HDLL__O21AI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O21AI_1%Y N_Y_M1003_d N_Y_M1001_d N_Y_c_153_n
+ N_Y_c_154_n N_Y_c_155_n N_Y_c_161_n N_Y_c_156_n Y Y
+ PM_SKY130_FD_SC_HDLL__O21AI_1%Y
x_PM_SKY130_FD_SC_HDLL__O21AI_1%A_27_47# N_A_27_47#_M1005_s N_A_27_47#_M1004_d
+ N_A_27_47#_c_186_n N_A_27_47#_c_188_n N_A_27_47#_c_187_n N_A_27_47#_c_199_n
+ PM_SKY130_FD_SC_HDLL__O21AI_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O21AI_1%VGND N_VGND_M1005_d VGND N_VGND_c_210_n
+ N_VGND_c_211_n N_VGND_c_212_n VGND PM_SKY130_FD_SC_HDLL__O21AI_1%VGND
cc_1 VNB N_A1_c_36_n 0.0316965f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A1_c_37_n 0.0232592f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_A1_c_38_n 0.0116706f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_4 VNB N_A2_c_58_n 0.0246767f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_A2_c_59_n 0.0172928f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_A2_c_60_n 0.00210258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B1_M1003_g 0.0398311f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_8 VNB B1 0.00645283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_97_n 0.0089532f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_10 VNB N_VPWR_c_125_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_153_n 0.0167221f $X=-0.19 $Y=-0.24 $X2=0.392 $Y2=1.16
cc_12 VNB N_Y_c_154_n 0.00272225f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_13 VNB N_Y_c_155_n 0.00435338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_156_n 0.0010487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_186_n 0.013695f $X=-0.19 $Y=-0.24 $X2=0.392 $Y2=1.16
cc_16 VNB N_A_27_47#_c_187_n 0.00894105f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_17 VNB N_VGND_c_210_n 0.0354053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_211_n 0.145639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_212_n 0.0275391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VPB N_A1_c_36_n 0.0332938f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_21 VPB N_A1_c_38_n 0.00110729f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_22 VPB N_A2_c_58_n 0.0266694f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_23 VPB A2 5.99582e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_A2_c_60_n 5.99582e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_B1_c_98_n 0.022107f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_26 VPB B1 0.0243014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_B1_c_97_n 0.0473384f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_28 VPB N_VPWR_c_126_n 0.0101063f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_29 VPB N_VPWR_c_127_n 0.0429248f $X=-0.19 $Y=1.305 $X2=0.392 $Y2=1.16
cc_30 VPB N_VPWR_c_128_n 0.01718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_129_n 0.00638493f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_32 VPB N_VPWR_c_130_n 0.0323231f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_125_n 0.04545f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_Y_c_156_n 0.00147285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB Y 7.333e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 N_A1_c_36_n N_A2_c_58_n 0.0966512f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_37 N_A1_c_38_n N_A2_c_58_n 2.10398e-19 $X=0.325 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_38 N_A1_c_37_n N_A2_c_59_n 0.0184238f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_39 N_A1_c_36_n A2 0.0301195f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_40 N_A1_c_36_n N_A2_c_60_n 0.0084031f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_41 N_A1_c_38_n N_A2_c_60_n 0.0252559f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_42 N_A1_c_36_n N_VPWR_c_127_n 0.0236794f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_43 N_A1_c_38_n N_VPWR_c_127_n 0.0193749f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_44 N_A1_c_36_n N_VPWR_c_130_n 0.00675582f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_45 N_A1_c_36_n N_VPWR_c_125_n 0.011085f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_46 N_A1_c_36_n N_A_27_47#_c_188_n 0.00143789f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_47 N_A1_c_37_n N_A_27_47#_c_188_n 0.0177313f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_48 N_A1_c_38_n N_A_27_47#_c_188_n 0.00116801f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_49 N_A1_c_36_n N_A_27_47#_c_187_n 0.00428914f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_50 N_A1_c_38_n N_A_27_47#_c_187_n 0.0163266f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_51 N_A1_c_37_n N_VGND_c_211_n 0.00686351f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_52 N_A1_c_37_n N_VGND_c_212_n 0.00743718f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_53 N_A2_c_59_n N_B1_M1003_g 0.0194743f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A2_c_60_n N_B1_M1003_g 2.92438e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A2_c_58_n N_B1_c_98_n 0.0126516f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_56 N_A2_c_58_n N_B1_c_97_n 0.0287948f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_57 A2 N_B1_c_97_n 2.76862e-19 $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_58 N_A2_c_58_n N_VPWR_c_127_n 0.00190657f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_59 A2 N_VPWR_c_127_n 0.064605f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_60 N_A2_c_58_n N_VPWR_c_130_n 0.00675913f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_61 A2 N_VPWR_c_130_n 0.00878874f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_62 N_A2_c_58_n N_VPWR_c_125_n 0.0122498f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_63 A2 N_VPWR_c_125_n 0.00917514f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_64 A2 A_117_297# 0.00136507f $X=0.605 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_65 N_A2_c_59_n N_Y_c_154_n 0.00221037f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_66 N_A2_c_60_n N_Y_c_154_n 0.0112424f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A2_c_58_n N_Y_c_161_n 0.00459576f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A2_c_60_n N_Y_c_161_n 0.00347315f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A2_c_58_n N_Y_c_156_n 0.00287984f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_70 A2 N_Y_c_156_n 0.00680409f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_71 N_A2_c_60_n N_Y_c_156_n 0.0154689f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A2_c_58_n N_A_27_47#_c_188_n 0.0044421f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A2_c_59_n N_A_27_47#_c_188_n 0.0131996f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_74 N_A2_c_60_n N_A_27_47#_c_188_n 0.0281481f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A2_c_59_n N_VGND_c_210_n 0.00365831f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A2_c_59_n N_VGND_c_211_n 0.00425872f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A2_c_59_n N_VGND_c_212_n 0.00781489f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B1_c_98_n N_VPWR_c_129_n 0.0177663f $X=1.505 $Y=1.71 $X2=0 $Y2=0
cc_79 B1 N_VPWR_c_129_n 0.0379919f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_80 N_B1_c_97_n N_VPWR_c_129_n 0.0019161f $X=1.505 $Y=1.502 $X2=0 $Y2=0
cc_81 N_B1_c_98_n N_VPWR_c_130_n 0.00702461f $X=1.505 $Y=1.71 $X2=0 $Y2=0
cc_82 N_B1_c_98_n N_VPWR_c_125_n 0.0140015f $X=1.505 $Y=1.71 $X2=0 $Y2=0
cc_83 N_B1_M1003_g N_Y_c_153_n 0.0183527f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_84 B1 N_Y_c_153_n 0.0395414f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_85 N_B1_c_97_n N_Y_c_153_n 0.00933449f $X=1.505 $Y=1.502 $X2=0 $Y2=0
cc_86 N_B1_M1003_g N_Y_c_154_n 0.00194183f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_87 N_B1_M1003_g N_Y_c_155_n 0.0190244f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_88 N_B1_c_97_n N_Y_c_161_n 0.00816564f $X=1.505 $Y=1.502 $X2=0 $Y2=0
cc_89 N_B1_M1003_g N_Y_c_156_n 0.00781833f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_90 B1 N_Y_c_156_n 0.0210024f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_91 N_B1_c_97_n N_Y_c_156_n 0.00563319f $X=1.505 $Y=1.502 $X2=0 $Y2=0
cc_92 N_B1_c_98_n Y 0.00251938f $X=1.505 $Y=1.71 $X2=0 $Y2=0
cc_93 N_B1_M1003_g N_A_27_47#_c_188_n 0.00120957f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_94 N_B1_M1003_g N_VGND_c_210_n 0.00585385f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_95 N_B1_M1003_g N_VGND_c_211_n 0.0122169f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_96 N_B1_M1003_g N_VGND_c_212_n 0.00130665f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_97 N_VPWR_c_125_n A_117_297# 0.00192225f $X=2.07 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_98 N_VPWR_c_125_n N_Y_M1001_d 0.00375648f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_99 N_VPWR_c_130_n Y 0.0251372f $X=1.645 $Y=2.72 $X2=0 $Y2=0
cc_100 N_VPWR_c_125_n Y 0.0157128f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_101 N_Y_c_154_n N_A_27_47#_c_188_n 0.0118985f $X=1.415 $Y=1.04 $X2=0 $Y2=0
cc_102 N_Y_c_155_n N_A_27_47#_c_188_n 0.0112667f $X=1.885 $Y=0.36 $X2=0 $Y2=0
cc_103 N_Y_c_155_n N_A_27_47#_c_199_n 0.0193857f $X=1.885 $Y=0.36 $X2=0 $Y2=0
cc_104 N_Y_c_155_n N_VGND_c_210_n 0.0288485f $X=1.885 $Y=0.36 $X2=0 $Y2=0
cc_105 N_Y_M1003_d N_VGND_c_211_n 0.00901528f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_106 N_Y_c_155_n N_VGND_c_211_n 0.0176597f $X=1.885 $Y=0.36 $X2=0 $Y2=0
cc_107 N_Y_c_155_n N_VGND_c_212_n 9.85286e-19 $X=1.885 $Y=0.36 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_188_n N_VGND_M1005_d 0.00601033f $X=1.175 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_27_47#_c_188_n N_VGND_c_210_n 0.00263539f $X=1.175 $Y=0.7 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_199_n N_VGND_c_210_n 0.00982795f $X=1.27 $Y=0.475 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_M1005_s N_VGND_c_211_n 0.00271326f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_M1004_d N_VGND_c_211_n 0.00231933f $X=1.135 $Y=0.235 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_186_n N_VGND_c_211_n 0.01096f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_188_n N_VGND_c_211_n 0.0121915f $X=1.175 $Y=0.7 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_199_n N_VGND_c_211_n 0.00844509f $X=1.27 $Y=0.475 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_186_n N_VGND_c_212_n 0.0187215f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_188_n N_VGND_c_212_n 0.0258321f $X=1.175 $Y=0.7 $X2=0 $Y2=0
