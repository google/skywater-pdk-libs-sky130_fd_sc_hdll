* File: sky130_fd_sc_hdll__and4b_4.spice
* Created: Wed Sep  2 08:23:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and4b_4.pex.spice"
.subckt sky130_fd_sc_hdll__and4b_4  VNB VPB A_N D C B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* C	C
* D	D
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_N_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1302 PD=0.765421 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1013_d N_A_184_21#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11785 AS=0.104 PD=1.18458 PS=0.97 NRD=9.228 NRS=8.304 M=1 R=4.33333
+ SA=75000.5 SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_184_21#_M1007_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1007_d N_A_184_21#_M1014_g N_X_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.5
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_184_21#_M1015_g N_X_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.15925 AS=0.104 PD=1.14 PS=0.97 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1002 A_624_47# N_D_M1002_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.15925 PD=0.97 PS=1.14 NRD=19.38 NRS=23.988 M=1 R=4.33333 SA=75002.6
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1001 A_718_47# N_C_M1001_g A_624_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.104 PD=0.98 PS=0.97 NRD=20.304 NRS=19.38 M=1 R=4.33333 SA=75003
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1005 A_814_47# N_B_M1005_g A_718_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.10725 PD=1.03 PS=0.98 NRD=24.912 NRS=20.304 M=1 R=4.33333 SA=75003.5
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1000 N_A_184_21#_M1000_d N_A_27_47#_M1000_g A_814_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.1235 PD=1.82 PS=1.03 NRD=0 NRS=24.912 M=1 R=4.33333 SA=75004.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_27_47#_M1003_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0874606 AS=0.1134 PD=0.795634 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90004.2 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1003_d N_A_184_21#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.208239 AS=0.145 PD=1.89437 PS=1.29 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.4 SB=90003.7 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_184_21#_M1010_g N_X_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.9 SB=90003.2 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1010_d N_A_184_21#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.3 SB=90002.8 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1017_d N_A_184_21#_M1017_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.205 AS=0.145 PD=1.41 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.8 SB=90002.3 A=0.18 P=2.36 MULT=1
MM1016 N_A_184_21#_M1016_d N_D_M1016_g N_VPWR_M1017_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.205 PD=1.29 PS=1.41 NRD=0.9653 NRS=24.6053 M=1 R=5.55556
+ SA=90002.4 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_C_M1009_g N_A_184_21#_M1016_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.145 PD=1.35 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.9 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1004 N_A_184_21#_M1004_d N_B_M1004_g N_VPWR_M1009_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=5.8903 NRS=12.7853 M=1 R=5.55556
+ SA=90003.4 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_27_47#_M1012_g N_A_184_21#_M1004_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.175 PD=2.54 PS=1.35 NRD=0.9653 NRS=7.8603 M=1 R=5.55556
+ SA=90003.9 SB=90000.2 A=0.18 P=2.36 MULT=1
DX18_noxref VNB VPB NWDIODE A=8.7312 P=14.09
pX19_noxref noxref_15 X X PROBETYPE=1
pX20_noxref noxref_16 X X PROBETYPE=1
pX21_noxref noxref_17 X X PROBETYPE=1
c_75 VPB 0 1.24891e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__and4b_4.pxi.spice"
*
.ends
*
*
