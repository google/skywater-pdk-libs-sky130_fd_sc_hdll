* File: sky130_fd_sc_hdll__o31ai_4.spice
* Created: Thu Aug 27 19:22:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o31ai_4.pex.spice"
.subckt sky130_fd_sc_hdll__o31ai_4  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_A_31_47#_M1003_d N_A1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75007.9 A=0.0975 P=1.6 MULT=1
MM1014 N_A_31_47#_M1014_d N_A1_M1014_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75007.4 A=0.0975 P=1.6 MULT=1
MM1015 N_A_31_47#_M1014_d N_A1_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75006.9 A=0.0975 P=1.6 MULT=1
MM1026 N_A_31_47#_M1026_d N_A1_M1026_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_31_47#_M1026_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75006 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1008_d N_A2_M1011_g N_A_31_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A2_M1021_g N_A_31_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1029 N_VGND_M1021_d N_A2_M1029_g N_A_31_47#_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A3_M1000_g N_A_31_47#_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.255125 AS=0.08775 PD=1.435 PS=0.92 NRD=22.152 NRS=0 M=1 R=4.33333
+ SA=75003.9 SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1000_d N_A3_M1017_g N_A_31_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.255125 AS=0.104 PD=1.435 PS=0.97 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75004.9 SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1023_d N_A3_M1023_g N_A_31_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.15925 AS=0.104 PD=1.14 PS=0.97 NRD=19.38 NRS=0 M=1 R=4.33333 SA=75005.3
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1023_d N_A3_M1027_g N_A_31_47#_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.15925 AS=0.08775 PD=1.14 PS=0.92 NRD=19.38 NRS=0 M=1 R=4.33333 SA=75006
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1004 N_A_31_47#_M1027_s N_B1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.4
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1009 N_A_31_47#_M1009_d N_B1_M1009_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006.9
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1012 N_A_31_47#_M1009_d N_B1_M1012_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75007.3
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1022 N_A_31_47#_M1022_d N_B1_M1022_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75007.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_27_297#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1002_d N_A1_M1006_g N_A_27_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90003 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A1_M1013_g N_A_27_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1013_d N_A1_M1020_g N_A_27_297#_M1020_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1001 N_A_497_297#_M1001_d N_A2_M1001_g N_A_27_297#_M1020_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1016 N_A_497_297#_M1001_d N_A2_M1016_g N_A_27_297#_M1016_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1024 N_A_497_297#_M1024_d N_A2_M1024_g N_A_27_297#_M1016_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1031 N_A_497_297#_M1024_d N_A2_M1031_g N_A_27_297#_M1031_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_Y_M1005_d N_A3_M1005_g N_A_497_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.295 AS=0.145 PD=2.59 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1007 N_Y_M1007_d N_A3_M1007_g N_A_497_297#_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90003 A=0.18 P=2.36 MULT=1
MM1018 N_Y_M1007_d N_A3_M1018_g N_A_497_297#_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1028 N_Y_M1028_d N_A3_M1028_g N_A_497_297#_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1010 N_Y_M1028_d N_B1_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1019 N_Y_M1019_d N_B1_M1019_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1025 N_Y_M1019_d N_B1_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1030 N_Y_M1030_d N_B1_M1030_g N_VPWR_M1025_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX32_noxref VNB VPB NWDIODE A=14.6376 P=21.45
*
.include "sky130_fd_sc_hdll__o31ai_4.pxi.spice"
*
.ends
*
*
