* File: sky130_fd_sc_hdll__dlxtn_1.pxi.spice
* Created: Thu Aug 27 19:06:13 2020
* 
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%GATE_N N_GATE_N_c_126_n N_GATE_N_c_127_n
+ N_GATE_N_M1001_g N_GATE_N_c_121_n N_GATE_N_M1012_g N_GATE_N_c_122_n GATE_N
+ GATE_N N_GATE_N_c_124_n N_GATE_N_c_125_n PM_SKY130_FD_SC_HDLL__DLXTN_1%GATE_N
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%A_27_47# N_A_27_47#_M1012_s N_A_27_47#_M1001_s
+ N_A_27_47#_c_172_n N_A_27_47#_c_173_n N_A_27_47#_M1015_g N_A_27_47#_M1000_g
+ N_A_27_47#_M1014_g N_A_27_47#_c_174_n N_A_27_47#_M1004_g N_A_27_47#_c_309_p
+ N_A_27_47#_c_163_n N_A_27_47#_c_164_n N_A_27_47#_c_175_n N_A_27_47#_c_176_n
+ N_A_27_47#_c_177_n N_A_27_47#_c_165_n N_A_27_47#_c_166_n N_A_27_47#_c_167_n
+ N_A_27_47#_c_168_n N_A_27_47#_c_179_n N_A_27_47#_c_180_n N_A_27_47#_c_181_n
+ N_A_27_47#_c_182_n N_A_27_47#_c_183_n N_A_27_47#_c_169_n N_A_27_47#_c_170_n
+ N_A_27_47#_c_171_n PM_SKY130_FD_SC_HDLL__DLXTN_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%D N_D_c_325_n N_D_c_330_n N_D_M1011_g
+ N_D_M1008_g D N_D_c_327_n N_D_c_328_n PM_SKY130_FD_SC_HDLL__DLXTN_1%D
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%A_319_47# N_A_319_47#_M1008_s
+ N_A_319_47#_M1011_s N_A_319_47#_c_368_n N_A_319_47#_c_376_n
+ N_A_319_47#_M1007_g N_A_319_47#_M1009_g N_A_319_47#_c_377_n
+ N_A_319_47#_c_369_n N_A_319_47#_c_378_n N_A_319_47#_c_379_n
+ N_A_319_47#_c_370_n N_A_319_47#_c_371_n N_A_319_47#_c_372_n
+ N_A_319_47#_c_373_n N_A_319_47#_c_374_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_1%A_319_47#
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%A_211_363# N_A_211_363#_M1000_d
+ N_A_211_363#_M1015_d N_A_211_363#_c_456_n N_A_211_363#_c_461_n
+ N_A_211_363#_c_462_n N_A_211_363#_M1017_g N_A_211_363#_c_457_n
+ N_A_211_363#_M1010_g N_A_211_363#_c_459_n N_A_211_363#_c_465_n
+ N_A_211_363#_c_466_n N_A_211_363#_c_467_n N_A_211_363#_c_468_n
+ N_A_211_363#_c_469_n N_A_211_363#_c_470_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_1%A_211_363#
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%A_760_21# N_A_760_21#_M1006_s
+ N_A_760_21#_M1002_s N_A_760_21#_M1016_g N_A_760_21#_c_572_n
+ N_A_760_21#_M1005_g N_A_760_21#_c_567_n N_A_760_21#_M1013_g
+ N_A_760_21#_c_568_n N_A_760_21#_M1003_g N_A_760_21#_c_574_n
+ N_A_760_21#_c_625_p N_A_760_21#_c_610_p N_A_760_21#_c_569_n
+ N_A_760_21#_c_575_n N_A_760_21#_c_570_n N_A_760_21#_c_591_p
+ N_A_760_21#_c_592_p N_A_760_21#_c_593_p
+ PM_SKY130_FD_SC_HDLL__DLXTN_1%A_760_21#
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%A_607_47# N_A_607_47#_M1014_d
+ N_A_607_47#_M1017_d N_A_607_47#_c_642_n N_A_607_47#_M1002_g
+ N_A_607_47#_c_636_n N_A_607_47#_M1006_g N_A_607_47#_c_637_n
+ N_A_607_47#_c_638_n N_A_607_47#_c_647_n N_A_607_47#_c_650_n
+ N_A_607_47#_c_639_n N_A_607_47#_c_645_n N_A_607_47#_c_640_n
+ N_A_607_47#_c_641_n PM_SKY130_FD_SC_HDLL__DLXTN_1%A_607_47#
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%VPWR N_VPWR_M1001_d N_VPWR_M1011_d
+ N_VPWR_M1005_d N_VPWR_M1002_d N_VPWR_c_719_n N_VPWR_c_720_n N_VPWR_c_721_n
+ N_VPWR_c_722_n N_VPWR_c_723_n N_VPWR_c_724_n N_VPWR_c_725_n N_VPWR_c_726_n
+ N_VPWR_c_727_n N_VPWR_c_728_n VPWR N_VPWR_c_729_n N_VPWR_c_730_n
+ N_VPWR_c_718_n N_VPWR_c_732_n PM_SKY130_FD_SC_HDLL__DLXTN_1%VPWR
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%Q N_Q_M1003_d N_Q_M1013_d Q Q Q
+ PM_SKY130_FD_SC_HDLL__DLXTN_1%Q
x_PM_SKY130_FD_SC_HDLL__DLXTN_1%VGND N_VGND_M1012_d N_VGND_M1008_d
+ N_VGND_M1016_d N_VGND_M1006_d N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n
+ N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n VGND N_VGND_c_830_n
+ N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n
+ PM_SKY130_FD_SC_HDLL__DLXTN_1%VGND
cc_1 VNB N_GATE_N_c_121_n 0.0173562f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_2 VNB N_GATE_N_c_122_n 0.0272334f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_3 VNB GATE_N 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_124_n 0.0217779f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_125_n 0.0136718f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1000_g 0.0409859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_163_n 0.00233896f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_8 VNB N_A_27_47#_c_164_n 0.00643242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_165_n 0.0013847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_166_n 0.00663785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_167_n 0.027628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_168_n 0.0024484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_169_n 0.0266603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_170_n 0.0177091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_171_n 0.00337398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_c_325_n 0.00677792f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.07
cc_17 VNB N_D_M1008_g 0.0259075f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_18 VNB N_D_c_327_n 0.00715095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_D_c_328_n 0.0452157f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_20 VNB N_A_319_47#_c_368_n 0.014357f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_21 VNB N_A_319_47#_c_369_n 0.00320313f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_22 VNB N_A_319_47#_c_370_n 0.00905692f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_23 VNB N_A_319_47#_c_371_n 0.00340984f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_24 VNB N_A_319_47#_c_372_n 0.00287801f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_25 VNB N_A_319_47#_c_373_n 0.0237537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_319_47#_c_374_n 0.0173868f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_211_363#_c_456_n 0.00586653f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_28 VNB N_A_211_363#_c_457_n 0.0107433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_211_363#_M1010_g 0.0463356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_211_363#_c_459_n 0.01415f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_31 VNB N_A_760_21#_M1016_g 0.0465371f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_32 VNB N_A_760_21#_c_567_n 0.0230716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_760_21#_c_568_n 0.02f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_34 VNB N_A_760_21#_c_569_n 0.00259455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_760_21#_c_570_n 0.00281539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_607_47#_c_636_n 0.0199493f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_37 VNB N_A_607_47#_c_637_n 0.0449172f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_38 VNB N_A_607_47#_c_638_n 0.0124501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_607_47#_c_639_n 0.00272011f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_40 VNB N_A_607_47#_c_640_n 0.00439888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_607_47#_c_641_n 0.00245432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_718_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB Q 0.0417654f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_44 VNB N_VGND_c_824_n 0.0169498f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_45 VNB N_VGND_c_825_n 0.00527913f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_46 VNB N_VGND_c_826_n 0.0450357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_827_n 0.00538573f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_48 VNB N_VGND_c_828_n 0.0213492f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_49 VNB N_VGND_c_829_n 0.00519339f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_50 VNB N_VGND_c_830_n 0.0154125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_831_n 0.0298657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_832_n 0.0221545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_833_n 0.318922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_834_n 0.0085923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_835_n 0.00556536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VPB N_GATE_N_c_126_n 0.0108902f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_57 VPB N_GATE_N_c_127_n 0.0470277f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_58 VPB GATE_N 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_59 VPB N_GATE_N_c_124_n 0.0110489f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_60 VPB N_A_27_47#_c_172_n 0.0196311f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_61 VPB N_A_27_47#_c_173_n 0.0261759f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_62 VPB N_A_27_47#_c_174_n 0.0511882f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_63 VPB N_A_27_47#_c_175_n 0.00146141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_47#_c_176_n 0.0046949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_47#_c_177_n 0.00363222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_165_n 6.22232e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_47#_c_179_n 0.0263712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_c_180_n 0.00387417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_c_181_n 0.00593858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_182_n 0.00279656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_183_n 0.00475048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_169_n 0.0120947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_171_n 2.90663e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_D_c_325_n 0.0240874f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.07
cc_75 VPB N_D_c_330_n 0.0271119f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_76 VPB N_D_c_327_n 0.00340154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_319_47#_c_368_n 0.0191152f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_78 VPB N_A_319_47#_c_376_n 0.0225552f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_79 VPB N_A_319_47#_c_377_n 0.00714124f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_80 VPB N_A_319_47#_c_378_n 0.00424606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_319_47#_c_379_n 0.00286464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_319_47#_c_371_n 0.00369206f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_83 VPB N_A_211_363#_c_456_n 0.0306708f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_84 VPB N_A_211_363#_c_461_n 0.0107952f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_85 VPB N_A_211_363#_c_462_n 0.0237245f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_86 VPB N_A_211_363#_c_457_n 0.0155543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_211_363#_c_459_n 0.00827089f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_88 VPB N_A_211_363#_c_465_n 0.00300202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_211_363#_c_466_n 0.00507872f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_90 VPB N_A_211_363#_c_467_n 0.00241696f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_91 VPB N_A_211_363#_c_468_n 0.0071704f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_92 VPB N_A_211_363#_c_469_n 0.00114173f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_93 VPB N_A_211_363#_c_470_n 0.0123773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_760_21#_M1016_g 0.0157901f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_95 VPB N_A_760_21#_c_572_n 0.0718489f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_96 VPB N_A_760_21#_c_567_n 0.0283374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_760_21#_c_574_n 0.00678594f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_98 VPB N_A_760_21#_c_575_n 0.00378052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_760_21#_c_570_n 0.00281539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_607_47#_c_642_n 0.0193905f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_101 VPB N_A_607_47#_c_637_n 0.0157968f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_102 VPB N_A_607_47#_c_638_n 0.00698873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_607_47#_c_645_n 0.00484721f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_104 VPB N_A_607_47#_c_640_n 0.00221288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_719_n 0.00126291f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_106 VPB N_VPWR_c_720_n 0.00367613f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_107 VPB N_VPWR_c_721_n 0.00980734f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_108 VPB N_VPWR_c_722_n 0.00205463f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_109 VPB N_VPWR_c_723_n 0.0326954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_724_n 0.00446482f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_111 VPB N_VPWR_c_725_n 0.0424754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_726_n 0.00574408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_727_n 0.019323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_728_n 0.0040431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_729_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_730_n 0.0204428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_718_n 0.0598916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_732_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB Q 0.048838f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_120 N_GATE_N_c_127_n N_A_27_47#_c_172_n 0.00641193f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_121 N_GATE_N_c_124_n N_A_27_47#_c_172_n 0.00265145f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_122 N_GATE_N_c_127_n N_A_27_47#_c_173_n 0.0182633f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_123 N_GATE_N_c_121_n N_A_27_47#_M1000_g 0.015454f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_124 N_GATE_N_c_125_n N_A_27_47#_M1000_g 0.00178537f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_125 N_GATE_N_c_121_n N_A_27_47#_c_163_n 0.00633651f $X=0.52 $Y=0.73 $X2=0
+ $Y2=0
cc_126 N_GATE_N_c_122_n N_A_27_47#_c_163_n 0.0136405f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_127 N_GATE_N_c_122_n N_A_27_47#_c_164_n 0.00657185f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_128 GATE_N N_A_27_47#_c_164_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_129 N_GATE_N_c_124_n N_A_27_47#_c_164_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_130 N_GATE_N_c_127_n N_A_27_47#_c_175_n 0.0185787f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_131 N_GATE_N_c_127_n N_A_27_47#_c_177_n 0.00836964f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_132 GATE_N N_A_27_47#_c_177_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_133 N_GATE_N_c_124_n N_A_27_47#_c_177_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_134 N_GATE_N_c_124_n N_A_27_47#_c_165_n 0.00207629f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_135 N_GATE_N_c_122_n N_A_27_47#_c_166_n 0.00186433f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_136 GATE_N N_A_27_47#_c_166_n 0.0250709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_137 N_GATE_N_c_125_n N_A_27_47#_c_166_n 6.20429e-19 $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_138 N_GATE_N_c_126_n N_A_27_47#_c_180_n 0.0015178f $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_139 N_GATE_N_c_127_n N_A_27_47#_c_180_n 0.00103413f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_140 GATE_N N_A_27_47#_c_180_n 0.00630136f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_141 N_GATE_N_c_126_n N_A_27_47#_c_181_n 4.6708e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_142 N_GATE_N_c_127_n N_A_27_47#_c_181_n 0.00432676f $X=0.495 $Y=1.74 $X2=0
+ $Y2=0
cc_143 GATE_N N_A_27_47#_c_169_n 0.00100538f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_144 N_GATE_N_c_124_n N_A_27_47#_c_169_n 0.0129544f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_145 N_GATE_N_c_127_n N_VPWR_c_719_n 0.0125197f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_146 N_GATE_N_c_127_n N_VPWR_c_729_n 0.00304525f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_147 N_GATE_N_c_127_n N_VPWR_c_718_n 0.00454898f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_148 N_GATE_N_c_121_n N_VGND_c_830_n 0.00198377f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_149 N_GATE_N_c_122_n N_VGND_c_830_n 6.41851e-19 $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_150 N_GATE_N_c_121_n N_VGND_c_833_n 0.00367064f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_151 N_GATE_N_c_121_n N_VGND_c_834_n 0.0142867f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_179_n N_D_c_325_n 0.00789696f $X=3.115 $Y=1.53 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_179_n N_D_c_327_n 0.0134197f $X=3.115 $Y=1.53 $X2=0 $Y2=0
cc_154 N_A_27_47#_M1000_g N_D_c_328_n 0.00523969f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_179_n N_A_319_47#_c_368_n 0.00625272f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_171_n N_A_319_47#_c_368_n 0.00364423f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_179_n N_A_319_47#_c_378_n 0.0135374f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_c_179_n N_A_319_47#_c_379_n 0.0114021f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_167_n N_A_319_47#_c_370_n 0.0010551f $X=2.97 $Y=0.87 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_168_n N_A_319_47#_c_370_n 0.0139508f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_179_n N_A_319_47#_c_370_n 0.00840141f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_171_n N_A_319_47#_c_370_n 0.00169583f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_179_n N_A_319_47#_c_371_n 0.0109087f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_167_n N_A_319_47#_c_373_n 0.0109791f $X=2.97 $Y=0.87 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_168_n N_A_319_47#_c_373_n 3.19436e-19 $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_171_n N_A_319_47#_c_373_n 2.98232e-19 $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_167_n N_A_319_47#_c_374_n 0.00201203f $X=2.97 $Y=0.87 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_168_n N_A_319_47#_c_374_n 2.06079e-19 $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_170_n N_A_319_47#_c_374_n 0.0198312f $X=2.97 $Y=0.705 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_174_n N_A_211_363#_c_456_n 0.0163105f $X=3.49 $Y=1.99 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_167_n N_A_211_363#_c_456_n 0.0183306f $X=2.97 $Y=0.87 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_168_n N_A_211_363#_c_456_n 0.00140109f $X=3.255 $Y=0.87
+ $X2=0 $Y2=0
cc_173 N_A_27_47#_c_179_n N_A_211_363#_c_456_n 0.00674363f $X=3.115 $Y=1.53
+ $X2=0 $Y2=0
cc_174 N_A_27_47#_c_182_n N_A_211_363#_c_456_n 0.00206946f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_171_n N_A_211_363#_c_456_n 0.002331f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_174_n N_A_211_363#_c_461_n 0.00360594f $X=3.49 $Y=1.99 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_183_n N_A_211_363#_c_461_n 0.002331f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_174_n N_A_211_363#_c_462_n 0.0169203f $X=3.49 $Y=1.99 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_176_n N_A_211_363#_c_462_n 0.00236706f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_180 N_A_27_47#_c_174_n N_A_211_363#_c_457_n 0.0139799f $X=3.49 $Y=1.99 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_168_n N_A_211_363#_c_457_n 0.00301645f $X=3.255 $Y=0.87
+ $X2=0 $Y2=0
cc_182 N_A_27_47#_c_179_n N_A_211_363#_c_457_n 0.00144279f $X=3.115 $Y=1.53
+ $X2=0 $Y2=0
cc_183 N_A_27_47#_c_182_n N_A_211_363#_c_457_n 0.00140625f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_183_n N_A_211_363#_c_457_n 0.00392485f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_171_n N_A_211_363#_c_457_n 0.0125072f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_167_n N_A_211_363#_M1010_g 0.0201193f $X=2.97 $Y=0.87 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_168_n N_A_211_363#_M1010_g 0.00775335f $X=3.255 $Y=0.87
+ $X2=0 $Y2=0
cc_188 N_A_27_47#_c_170_n N_A_211_363#_M1010_g 0.0123046f $X=2.97 $Y=0.705 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_171_n N_A_211_363#_M1010_g 0.00649688f $X=3.34 $Y=1.415
+ $X2=0 $Y2=0
cc_190 N_A_27_47#_M1000_g N_A_211_363#_c_459_n 0.0112065f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_163_n N_A_211_363#_c_459_n 0.00937011f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_165_n N_A_211_363#_c_459_n 0.0196553f $X=0.805 $Y=1.235
+ $X2=0 $Y2=0
cc_193 N_A_27_47#_c_166_n N_A_211_363#_c_459_n 0.0138555f $X=0.775 $Y=1.07 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_179_n N_A_211_363#_c_459_n 0.0187427f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_180_n N_A_211_363#_c_459_n 0.00220079f $X=0.89 $Y=1.53 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_181_n N_A_211_363#_c_459_n 0.0175551f $X=0.745 $Y=1.53 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_172_n N_A_211_363#_c_465_n 0.0112065f $X=0.965 $Y=1.64 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_173_n N_A_211_363#_c_465_n 0.00723076f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_199 N_A_27_47#_c_175_n N_A_211_363#_c_465_n 0.00387314f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_179_n N_A_211_363#_c_465_n 0.00195186f $X=3.115 $Y=1.53
+ $X2=0 $Y2=0
cc_201 N_A_27_47#_c_179_n N_A_211_363#_c_466_n 0.0950762f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_173_n N_A_211_363#_c_467_n 0.00459592f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_203 N_A_27_47#_c_175_n N_A_211_363#_c_467_n 0.00534864f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_179_n N_A_211_363#_c_467_n 0.0259095f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_181_n N_A_211_363#_c_467_n 0.00107077f $X=0.745 $Y=1.53
+ $X2=0 $Y2=0
cc_206 N_A_27_47#_c_176_n N_A_211_363#_c_469_n 0.00155242f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_207 N_A_27_47#_c_179_n N_A_211_363#_c_469_n 0.0255946f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_174_n N_A_211_363#_c_470_n 3.98959e-19 $X=3.49 $Y=1.99 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_167_n N_A_211_363#_c_470_n 5.31837e-19 $X=2.97 $Y=0.87 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_168_n N_A_211_363#_c_470_n 0.00286407f $X=3.255 $Y=0.87
+ $X2=0 $Y2=0
cc_211 N_A_27_47#_c_179_n N_A_211_363#_c_470_n 0.0237184f $X=3.115 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_182_n N_A_211_363#_c_470_n 0.00264902f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_171_n N_A_211_363#_c_470_n 0.0367681f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_168_n N_A_760_21#_M1016_g 3.00559e-19 $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_183_n N_A_760_21#_M1016_g 5.23954e-19 $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_171_n N_A_760_21#_M1016_g 4.28547e-19 $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_174_n N_A_760_21#_c_572_n 0.0589955f $X=3.49 $Y=1.99 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_176_n N_A_760_21#_c_572_n 8.63256e-19 $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_167_n N_A_607_47#_c_647_n 0.00144439f $X=2.97 $Y=0.87 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_168_n N_A_607_47#_c_647_n 0.0202428f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_170_n N_A_607_47#_c_647_n 0.00433832f $X=2.97 $Y=0.705 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_174_n N_A_607_47#_c_650_n 0.0142229f $X=3.49 $Y=1.99 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_176_n N_A_607_47#_c_650_n 0.0156588f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_182_n N_A_607_47#_c_650_n 0.00267734f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_168_n N_A_607_47#_c_639_n 0.0132672f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_174_n N_A_607_47#_c_645_n 0.00808669f $X=3.49 $Y=1.99 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_182_n N_A_607_47#_c_645_n 0.00129859f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_183_n N_A_607_47#_c_645_n 0.043119f $X=3.26 $Y=1.53 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_171_n N_A_607_47#_c_645_n 0.00387486f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_168_n N_A_607_47#_c_641_n 0.00201058f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_171_n N_A_607_47#_c_641_n 0.0139727f $X=3.34 $Y=1.415 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_175_n N_VPWR_M1001_d 0.0022997f $X=0.66 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_233 N_A_27_47#_c_173_n N_VPWR_c_719_n 0.00977612f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_175_n N_VPWR_c_719_n 0.0196375f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_177_n N_VPWR_c_719_n 0.0246493f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_180_n N_VPWR_c_719_n 0.00314061f $X=0.89 $Y=1.53 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_179_n N_VPWR_c_720_n 0.0018348f $X=3.115 $Y=1.53 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_173_n N_VPWR_c_723_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_174_n N_VPWR_c_725_n 0.00439333f $X=3.49 $Y=1.99 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_175_n N_VPWR_c_729_n 0.00180073f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_177_n N_VPWR_c_729_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_173_n N_VPWR_c_718_n 0.0113647f $X=0.965 $Y=1.74 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_174_n N_VPWR_c_718_n 0.00618212f $X=3.49 $Y=1.99 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_175_n N_VPWR_c_718_n 0.00504362f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_177_n N_VPWR_c_718_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_163_n N_VGND_M1012_d 0.00215196f $X=0.66 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_247 N_A_27_47#_c_167_n N_VGND_c_826_n 9.43262e-19 $X=2.97 $Y=0.87 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_168_n N_VGND_c_826_n 0.00175247f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_170_n N_VGND_c_826_n 0.00424048f $X=2.97 $Y=0.705 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_309_p N_VGND_c_830_n 0.00725596f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_163_n N_VGND_c_830_n 0.00244154f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_252 N_A_27_47#_M1000_g N_VGND_c_831_n 0.00585385f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_M1012_s N_VGND_c_833_n 0.00437169f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_M1000_g N_VGND_c_833_n 0.0120602f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_309_p N_VGND_c_833_n 0.00608739f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_163_n N_VGND_c_833_n 0.00595002f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_167_n N_VGND_c_833_n 0.00121904f $X=2.97 $Y=0.87 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_168_n N_VGND_c_833_n 0.00332341f $X=3.255 $Y=0.87 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_170_n N_VGND_c_833_n 0.00629139f $X=2.97 $Y=0.705 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1000_g N_VGND_c_834_n 0.00317372f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_309_p N_VGND_c_834_n 0.00895866f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_163_n N_VGND_c_834_n 0.0205047f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_165_n N_VGND_c_834_n 0.00148975f $X=0.805 $Y=1.235 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_169_n N_VGND_c_834_n 7.59537e-19 $X=0.99 $Y=1.235 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_170_n N_VGND_c_835_n 0.00168882f $X=2.97 $Y=0.705 $X2=0
+ $Y2=0
cc_266 N_D_c_328_n N_A_319_47#_c_368_n 0.0145035f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_267 N_D_c_325_n N_A_319_47#_c_376_n 0.0145035f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_268 N_D_c_330_n N_A_319_47#_c_376_n 0.00935018f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_269 N_D_c_330_n N_A_319_47#_c_377_n 0.0136011f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_270 N_D_M1008_g N_A_319_47#_c_369_n 0.0152747f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_271 N_D_c_327_n N_A_319_47#_c_369_n 0.00639931f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_272 N_D_c_328_n N_A_319_47#_c_369_n 0.0029398f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_273 N_D_c_325_n N_A_319_47#_c_378_n 0.0106635f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_274 N_D_c_325_n N_A_319_47#_c_379_n 0.00412429f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_275 N_D_c_327_n N_A_319_47#_c_379_n 0.0233961f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_276 N_D_c_328_n N_A_319_47#_c_379_n 0.00131849f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_277 N_D_M1008_g N_A_319_47#_c_370_n 0.00591272f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_278 N_D_c_327_n N_A_319_47#_c_370_n 0.00920968f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_279 N_D_c_327_n N_A_319_47#_c_371_n 0.013986f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_280 N_D_c_328_n N_A_319_47#_c_371_n 0.0057769f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_281 N_D_M1008_g N_A_319_47#_c_372_n 8.59557e-19 $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_282 N_D_c_327_n N_A_319_47#_c_372_n 0.0138491f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_283 N_D_c_328_n N_A_319_47#_c_372_n 0.0042466f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_284 N_D_M1008_g N_A_319_47#_c_373_n 0.0198331f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_285 N_D_M1008_g N_A_319_47#_c_374_n 0.0140113f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_286 N_D_c_325_n N_A_211_363#_c_459_n 0.00463913f $X=1.955 $Y=1.67 $X2=0 $Y2=0
cc_287 N_D_M1008_g N_A_211_363#_c_459_n 0.00193515f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_288 N_D_c_327_n N_A_211_363#_c_459_n 0.0287516f $X=1.725 $Y=1.04 $X2=0 $Y2=0
cc_289 N_D_c_328_n N_A_211_363#_c_459_n 0.00236382f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_290 N_D_c_330_n N_A_211_363#_c_465_n 0.00132248f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_291 N_D_c_330_n N_A_211_363#_c_466_n 0.00420236f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_292 N_D_c_330_n N_VPWR_c_720_n 0.00664063f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_293 N_D_c_330_n N_VPWR_c_723_n 0.00674916f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_294 N_D_c_330_n N_VPWR_c_718_n 0.00848136f $X=1.955 $Y=1.77 $X2=0 $Y2=0
cc_295 N_D_M1008_g N_VGND_c_831_n 0.00196986f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_296 N_D_M1008_g N_VGND_c_833_n 0.00398772f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_297 N_D_c_328_n N_VGND_c_833_n 0.00103829f $X=1.98 $Y=1.04 $X2=0 $Y2=0
cc_298 N_D_M1008_g N_VGND_c_835_n 0.0140914f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_299 N_A_319_47#_c_368_n N_A_211_363#_c_456_n 0.0253115f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_300 N_A_319_47#_c_376_n N_A_211_363#_c_461_n 0.0107827f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_301 N_A_319_47#_c_376_n N_A_211_363#_c_462_n 0.0228578f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_302 N_A_319_47#_c_377_n N_A_211_363#_c_459_n 0.0010921f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_303 N_A_319_47#_c_379_n N_A_211_363#_c_459_n 0.00880329f $X=1.885 $Y=1.58
+ $X2=0 $Y2=0
cc_304 N_A_319_47#_c_372_n N_A_211_363#_c_459_n 0.0191835f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_305 N_A_319_47#_c_377_n N_A_211_363#_c_465_n 0.0471073f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_306 N_A_319_47#_c_376_n N_A_211_363#_c_466_n 0.00505686f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_307 N_A_319_47#_c_377_n N_A_211_363#_c_466_n 0.0230027f $X=1.72 $Y=1.99 $X2=0
+ $Y2=0
cc_308 N_A_319_47#_c_378_n N_A_211_363#_c_466_n 0.00667484f $X=2.12 $Y=1.58
+ $X2=0 $Y2=0
cc_309 N_A_319_47#_c_377_n N_A_211_363#_c_467_n 0.00273055f $X=1.72 $Y=1.99
+ $X2=0 $Y2=0
cc_310 N_A_319_47#_c_376_n N_A_211_363#_c_469_n 0.00149778f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_311 N_A_319_47#_c_368_n N_A_211_363#_c_470_n 0.00472707f $X=2.425 $Y=1.67
+ $X2=0 $Y2=0
cc_312 N_A_319_47#_c_376_n N_A_211_363#_c_470_n 0.00231211f $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_313 N_A_319_47#_c_378_n N_A_211_363#_c_470_n 0.00664087f $X=2.12 $Y=1.58
+ $X2=0 $Y2=0
cc_314 N_A_319_47#_c_371_n N_A_211_363#_c_470_n 0.00578855f $X=2.205 $Y=1.495
+ $X2=0 $Y2=0
cc_315 N_A_319_47#_c_374_n N_A_607_47#_c_647_n 6.60835e-19 $X=2.405 $Y=0.765
+ $X2=0 $Y2=0
cc_316 N_A_319_47#_c_376_n N_A_607_47#_c_650_n 4.97528e-19 $X=2.425 $Y=1.77
+ $X2=0 $Y2=0
cc_317 N_A_319_47#_c_376_n N_VPWR_c_720_n 0.022734f $X=2.425 $Y=1.77 $X2=0 $Y2=0
cc_318 N_A_319_47#_c_377_n N_VPWR_c_720_n 0.0355228f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_319 N_A_319_47#_c_378_n N_VPWR_c_720_n 0.013562f $X=2.12 $Y=1.58 $X2=0 $Y2=0
cc_320 N_A_319_47#_c_377_n N_VPWR_c_723_n 0.0159613f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_321 N_A_319_47#_c_376_n N_VPWR_c_725_n 0.00368966f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_322 N_A_319_47#_M1011_s N_VPWR_c_718_n 0.00181388f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_323 N_A_319_47#_c_376_n N_VPWR_c_718_n 0.00385316f $X=2.425 $Y=1.77 $X2=0
+ $Y2=0
cc_324 N_A_319_47#_c_377_n N_VPWR_c_718_n 0.0057885f $X=1.72 $Y=1.99 $X2=0 $Y2=0
cc_325 N_A_319_47#_c_370_n N_VGND_M1008_d 0.00178147f $X=2.205 $Y=1.095 $X2=0
+ $Y2=0
cc_326 N_A_319_47#_c_373_n N_VGND_c_826_n 3.25575e-19 $X=2.405 $Y=0.93 $X2=0
+ $Y2=0
cc_327 N_A_319_47#_c_374_n N_VGND_c_826_n 0.00546359f $X=2.405 $Y=0.765 $X2=0
+ $Y2=0
cc_328 N_A_319_47#_c_369_n N_VGND_c_831_n 0.00256875f $X=2.12 $Y=0.7 $X2=0 $Y2=0
cc_329 N_A_319_47#_c_372_n N_VGND_c_831_n 0.00723406f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_330 N_A_319_47#_M1008_s N_VGND_c_833_n 0.00343585f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_331 N_A_319_47#_c_369_n N_VGND_c_833_n 0.0051978f $X=2.12 $Y=0.7 $X2=0 $Y2=0
cc_332 N_A_319_47#_c_370_n N_VGND_c_833_n 0.00720854f $X=2.205 $Y=1.095 $X2=0
+ $Y2=0
cc_333 N_A_319_47#_c_372_n N_VGND_c_833_n 0.00607883f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_334 N_A_319_47#_c_374_n N_VGND_c_833_n 0.00516246f $X=2.405 $Y=0.765 $X2=0
+ $Y2=0
cc_335 N_A_319_47#_c_369_n N_VGND_c_835_n 0.00613814f $X=2.12 $Y=0.7 $X2=0 $Y2=0
cc_336 N_A_319_47#_c_370_n N_VGND_c_835_n 0.0153831f $X=2.205 $Y=1.095 $X2=0
+ $Y2=0
cc_337 N_A_319_47#_c_372_n N_VGND_c_835_n 0.00746555f $X=1.72 $Y=0.51 $X2=0
+ $Y2=0
cc_338 N_A_319_47#_c_374_n N_VGND_c_835_n 0.00852549f $X=2.405 $Y=0.765 $X2=0
+ $Y2=0
cc_339 N_A_211_363#_M1010_g N_A_760_21#_M1016_g 0.0463008f $X=3.4 $Y=0.415 $X2=0
+ $Y2=0
cc_340 N_A_211_363#_M1010_g N_A_607_47#_c_647_n 0.0127111f $X=3.4 $Y=0.415 $X2=0
+ $Y2=0
cc_341 N_A_211_363#_c_462_n N_A_607_47#_c_650_n 0.00429541f $X=2.95 $Y=1.99
+ $X2=0 $Y2=0
cc_342 N_A_211_363#_M1010_g N_A_607_47#_c_639_n 0.0055762f $X=3.4 $Y=0.415 $X2=0
+ $Y2=0
cc_343 N_A_211_363#_c_457_n N_A_607_47#_c_645_n 6.15458e-19 $X=3.325 $Y=1.32
+ $X2=0 $Y2=0
cc_344 N_A_211_363#_M1010_g N_A_607_47#_c_641_n 0.00305873f $X=3.4 $Y=0.415
+ $X2=0 $Y2=0
cc_345 N_A_211_363#_c_466_n N_VPWR_M1011_d 8.51638e-19 $X=2.61 $Y=1.87 $X2=0
+ $Y2=0
cc_346 N_A_211_363#_c_468_n N_VPWR_c_719_n 0.0206383f $X=1.255 $Y=1.87 $X2=0
+ $Y2=0
cc_347 N_A_211_363#_c_462_n N_VPWR_c_720_n 0.00315507f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_348 N_A_211_363#_c_466_n N_VPWR_c_720_n 0.017675f $X=2.61 $Y=1.87 $X2=0 $Y2=0
cc_349 N_A_211_363#_c_469_n N_VPWR_c_720_n 0.00130564f $X=2.755 $Y=1.87 $X2=0
+ $Y2=0
cc_350 N_A_211_363#_c_470_n N_VPWR_c_720_n 0.00772079f $X=2.87 $Y=1.52 $X2=0
+ $Y2=0
cc_351 N_A_211_363#_c_468_n N_VPWR_c_723_n 0.015988f $X=1.255 $Y=1.87 $X2=0
+ $Y2=0
cc_352 N_A_211_363#_c_462_n N_VPWR_c_725_n 0.00583292f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_353 N_A_211_363#_c_470_n N_VPWR_c_725_n 0.00457854f $X=2.87 $Y=1.52 $X2=0
+ $Y2=0
cc_354 N_A_211_363#_c_462_n N_VPWR_c_718_n 0.00923621f $X=2.95 $Y=1.99 $X2=0
+ $Y2=0
cc_355 N_A_211_363#_c_466_n N_VPWR_c_718_n 0.0567835f $X=2.61 $Y=1.87 $X2=0
+ $Y2=0
cc_356 N_A_211_363#_c_467_n N_VPWR_c_718_n 0.0152065f $X=1.4 $Y=1.87 $X2=0 $Y2=0
cc_357 N_A_211_363#_c_468_n N_VPWR_c_718_n 0.00389918f $X=1.255 $Y=1.87 $X2=0
+ $Y2=0
cc_358 N_A_211_363#_c_469_n N_VPWR_c_718_n 0.0151073f $X=2.755 $Y=1.87 $X2=0
+ $Y2=0
cc_359 N_A_211_363#_c_470_n N_VPWR_c_718_n 0.00405108f $X=2.87 $Y=1.52 $X2=0
+ $Y2=0
cc_360 N_A_211_363#_c_466_n A_503_369# 0.00150032f $X=2.61 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_361 N_A_211_363#_c_469_n A_503_369# 0.00122092f $X=2.755 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_362 N_A_211_363#_c_470_n A_503_369# 0.0032229f $X=2.87 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_363 N_A_211_363#_M1010_g N_VGND_c_826_n 0.0037981f $X=3.4 $Y=0.415 $X2=0
+ $Y2=0
cc_364 N_A_211_363#_c_459_n N_VGND_c_831_n 0.00732874f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_365 N_A_211_363#_M1000_d N_VGND_c_833_n 0.00535012f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_366 N_A_211_363#_M1010_g N_VGND_c_833_n 0.00558435f $X=3.4 $Y=0.415 $X2=0
+ $Y2=0
cc_367 N_A_211_363#_c_459_n N_VGND_c_833_n 0.00616598f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_368 N_A_760_21#_c_572_n N_A_607_47#_c_642_n 0.00329184f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_369 N_A_760_21#_c_567_n N_A_607_47#_c_642_n 0.0185382f $X=5.37 $Y=1.41 $X2=0
+ $Y2=0
cc_370 N_A_760_21#_c_575_n N_A_607_47#_c_642_n 0.00413095f $X=4.705 $Y=1.535
+ $X2=0 $Y2=0
cc_371 N_A_760_21#_c_568_n N_A_607_47#_c_636_n 0.0169359f $X=5.395 $Y=0.995
+ $X2=0 $Y2=0
cc_372 N_A_760_21#_c_569_n N_A_607_47#_c_636_n 0.00635275f $X=4.705 $Y=0.995
+ $X2=0 $Y2=0
cc_373 N_A_760_21#_M1016_g N_A_607_47#_c_637_n 0.01646f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_374 N_A_760_21#_c_572_n N_A_607_47#_c_637_n 0.00487525f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_375 N_A_760_21#_c_574_n N_A_607_47#_c_637_n 0.00879412f $X=4.57 $Y=1.7 $X2=0
+ $Y2=0
cc_376 N_A_760_21#_c_591_p N_A_607_47#_c_637_n 0.00203472f $X=4.68 $Y=0.825
+ $X2=0 $Y2=0
cc_377 N_A_760_21#_c_592_p N_A_607_47#_c_637_n 0.00212837f $X=4.655 $Y=1.755
+ $X2=0 $Y2=0
cc_378 N_A_760_21#_c_593_p N_A_607_47#_c_637_n 0.0181912f $X=4.705 $Y=1.16 $X2=0
+ $Y2=0
cc_379 N_A_760_21#_c_567_n N_A_607_47#_c_638_n 0.0252983f $X=5.37 $Y=1.41 $X2=0
+ $Y2=0
cc_380 N_A_760_21#_c_575_n N_A_607_47#_c_638_n 0.0036022f $X=4.705 $Y=1.535
+ $X2=0 $Y2=0
cc_381 N_A_760_21#_c_570_n N_A_607_47#_c_638_n 0.0276191f $X=5.335 $Y=1.16 $X2=0
+ $Y2=0
cc_382 N_A_760_21#_M1016_g N_A_607_47#_c_647_n 0.00502711f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_383 N_A_760_21#_c_572_n N_A_607_47#_c_650_n 0.00434287f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_384 N_A_760_21#_M1016_g N_A_607_47#_c_639_n 0.0142483f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_385 N_A_760_21#_M1016_g N_A_607_47#_c_645_n 0.0116647f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_386 N_A_760_21#_c_572_n N_A_607_47#_c_645_n 0.0243839f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_387 N_A_760_21#_c_574_n N_A_607_47#_c_645_n 0.0204069f $X=4.57 $Y=1.7 $X2=0
+ $Y2=0
cc_388 N_A_760_21#_M1016_g N_A_607_47#_c_640_n 0.0161022f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_389 N_A_760_21#_c_572_n N_A_607_47#_c_640_n 0.00820473f $X=3.9 $Y=1.99 $X2=0
+ $Y2=0
cc_390 N_A_760_21#_c_574_n N_A_607_47#_c_640_n 0.02399f $X=4.57 $Y=1.7 $X2=0
+ $Y2=0
cc_391 N_A_760_21#_c_593_p N_A_607_47#_c_640_n 0.0253721f $X=4.705 $Y=1.16 $X2=0
+ $Y2=0
cc_392 N_A_760_21#_M1016_g N_A_607_47#_c_641_n 0.00407241f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_393 N_A_760_21#_c_572_n N_VPWR_c_721_n 0.0124315f $X=3.9 $Y=1.99 $X2=0 $Y2=0
cc_394 N_A_760_21#_c_574_n N_VPWR_c_721_n 0.0154822f $X=4.57 $Y=1.7 $X2=0 $Y2=0
cc_395 N_A_760_21#_c_610_p N_VPWR_c_721_n 0.0196385f $X=4.655 $Y=2.27 $X2=0
+ $Y2=0
cc_396 N_A_760_21#_c_567_n N_VPWR_c_722_n 0.0227159f $X=5.37 $Y=1.41 $X2=0 $Y2=0
cc_397 N_A_760_21#_c_570_n N_VPWR_c_722_n 0.0195663f $X=5.335 $Y=1.16 $X2=0
+ $Y2=0
cc_398 N_A_760_21#_c_572_n N_VPWR_c_725_n 0.00665561f $X=3.9 $Y=1.99 $X2=0 $Y2=0
cc_399 N_A_760_21#_c_610_p N_VPWR_c_727_n 0.0115253f $X=4.655 $Y=2.27 $X2=0
+ $Y2=0
cc_400 N_A_760_21#_c_567_n N_VPWR_c_730_n 0.00661659f $X=5.37 $Y=1.41 $X2=0
+ $Y2=0
cc_401 N_A_760_21#_M1002_s N_VPWR_c_718_n 0.00284579f $X=4.53 $Y=1.485 $X2=0
+ $Y2=0
cc_402 N_A_760_21#_c_572_n N_VPWR_c_718_n 0.0136422f $X=3.9 $Y=1.99 $X2=0 $Y2=0
cc_403 N_A_760_21#_c_567_n N_VPWR_c_718_n 0.0121339f $X=5.37 $Y=1.41 $X2=0 $Y2=0
cc_404 N_A_760_21#_c_574_n N_VPWR_c_718_n 0.00898578f $X=4.57 $Y=1.7 $X2=0 $Y2=0
cc_405 N_A_760_21#_c_610_p N_VPWR_c_718_n 0.00827281f $X=4.655 $Y=2.27 $X2=0
+ $Y2=0
cc_406 N_A_760_21#_c_567_n Q 0.0252263f $X=5.37 $Y=1.41 $X2=0 $Y2=0
cc_407 N_A_760_21#_c_568_n Q 0.0267384f $X=5.395 $Y=0.995 $X2=0 $Y2=0
cc_408 N_A_760_21#_c_570_n Q 0.0272217f $X=5.335 $Y=1.16 $X2=0 $Y2=0
cc_409 N_A_760_21#_M1016_g N_VGND_c_824_n 0.0122754f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_410 N_A_760_21#_c_625_p N_VGND_c_824_n 0.0230546f $X=4.655 $Y=0.58 $X2=0
+ $Y2=0
cc_411 N_A_760_21#_c_567_n N_VGND_c_825_n 0.00204045f $X=5.37 $Y=1.41 $X2=0
+ $Y2=0
cc_412 N_A_760_21#_c_568_n N_VGND_c_825_n 0.00404192f $X=5.395 $Y=0.995 $X2=0
+ $Y2=0
cc_413 N_A_760_21#_c_570_n N_VGND_c_825_n 0.0205335f $X=5.335 $Y=1.16 $X2=0
+ $Y2=0
cc_414 N_A_760_21#_M1016_g N_VGND_c_826_n 0.00516796f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_415 N_A_760_21#_c_625_p N_VGND_c_828_n 0.00732441f $X=4.655 $Y=0.58 $X2=0
+ $Y2=0
cc_416 N_A_760_21#_c_568_n N_VGND_c_832_n 0.00585385f $X=5.395 $Y=0.995 $X2=0
+ $Y2=0
cc_417 N_A_760_21#_M1006_s N_VGND_c_833_n 0.00589711f $X=4.53 $Y=0.235 $X2=0
+ $Y2=0
cc_418 N_A_760_21#_M1016_g N_VGND_c_833_n 0.0104553f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_760_21#_c_568_n N_VGND_c_833_n 0.0119007f $X=5.395 $Y=0.995 $X2=0
+ $Y2=0
cc_420 N_A_760_21#_c_625_p N_VGND_c_833_n 0.00762661f $X=4.655 $Y=0.58 $X2=0
+ $Y2=0
cc_421 N_A_607_47#_c_650_n N_VPWR_c_720_n 0.00469266f $X=3.68 $Y=2.34 $X2=0
+ $Y2=0
cc_422 N_A_607_47#_c_642_n N_VPWR_c_721_n 0.00253117f $X=4.89 $Y=1.41 $X2=0
+ $Y2=0
cc_423 N_A_607_47#_c_650_n N_VPWR_c_721_n 0.0122631f $X=3.68 $Y=2.34 $X2=0 $Y2=0
cc_424 N_A_607_47#_c_645_n N_VPWR_c_721_n 0.00774669f $X=3.765 $Y=2.255 $X2=0
+ $Y2=0
cc_425 N_A_607_47#_c_642_n N_VPWR_c_722_n 0.00284809f $X=4.89 $Y=1.41 $X2=0
+ $Y2=0
cc_426 N_A_607_47#_c_650_n N_VPWR_c_725_n 0.0370617f $X=3.68 $Y=2.34 $X2=0 $Y2=0
cc_427 N_A_607_47#_c_642_n N_VPWR_c_727_n 0.00702461f $X=4.89 $Y=1.41 $X2=0
+ $Y2=0
cc_428 N_A_607_47#_M1017_d N_VPWR_c_718_n 0.00291507f $X=3.04 $Y=2.065 $X2=0
+ $Y2=0
cc_429 N_A_607_47#_c_642_n N_VPWR_c_718_n 0.0139178f $X=4.89 $Y=1.41 $X2=0 $Y2=0
cc_430 N_A_607_47#_c_650_n N_VPWR_c_718_n 0.0292009f $X=3.68 $Y=2.34 $X2=0 $Y2=0
cc_431 N_A_607_47#_c_650_n A_716_413# 0.00279977f $X=3.68 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_432 N_A_607_47#_c_645_n A_716_413# 0.00210862f $X=3.765 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_433 N_A_607_47#_c_636_n N_VGND_c_824_n 0.00673308f $X=4.915 $Y=0.995 $X2=0
+ $Y2=0
cc_434 N_A_607_47#_c_637_n N_VGND_c_824_n 0.00207331f $X=4.79 $Y=1.16 $X2=0
+ $Y2=0
cc_435 N_A_607_47#_c_647_n N_VGND_c_824_n 0.0138426f $X=3.68 $Y=0.45 $X2=0 $Y2=0
cc_436 N_A_607_47#_c_639_n N_VGND_c_824_n 0.0213894f $X=3.765 $Y=0.995 $X2=0
+ $Y2=0
cc_437 N_A_607_47#_c_640_n N_VGND_c_824_n 0.0242249f $X=4.345 $Y=1.16 $X2=0
+ $Y2=0
cc_438 N_A_607_47#_c_636_n N_VGND_c_825_n 0.00404192f $X=4.915 $Y=0.995 $X2=0
+ $Y2=0
cc_439 N_A_607_47#_c_647_n N_VGND_c_826_n 0.027917f $X=3.68 $Y=0.45 $X2=0 $Y2=0
cc_440 N_A_607_47#_c_636_n N_VGND_c_828_n 0.00585385f $X=4.915 $Y=0.995 $X2=0
+ $Y2=0
cc_441 N_A_607_47#_M1014_d N_VGND_c_833_n 0.00246479f $X=3.035 $Y=0.235 $X2=0
+ $Y2=0
cc_442 N_A_607_47#_c_636_n N_VGND_c_833_n 0.0121898f $X=4.915 $Y=0.995 $X2=0
+ $Y2=0
cc_443 N_A_607_47#_c_647_n N_VGND_c_833_n 0.0284427f $X=3.68 $Y=0.45 $X2=0 $Y2=0
cc_444 N_A_607_47#_c_647_n N_VGND_c_835_n 0.00207581f $X=3.68 $Y=0.45 $X2=0
+ $Y2=0
cc_445 N_A_607_47#_c_647_n A_695_47# 0.00809944f $X=3.68 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_446 N_A_607_47#_c_639_n A_695_47# 0.00141478f $X=3.765 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_447 N_VPWR_c_718_n A_503_369# 0.00393797f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_448 N_VPWR_c_718_n A_716_413# 0.00186715f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_449 N_VPWR_c_718_n N_Q_M1013_d 0.00730742f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_450 N_VPWR_c_722_n Q 0.046975f $X=5.125 $Y=1.735 $X2=0 $Y2=0
cc_451 N_VPWR_c_730_n Q 0.018801f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_452 N_VPWR_c_718_n Q 0.0108473f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_453 Q N_VGND_c_832_n 0.0097883f $X=5.645 $Y=0.425 $X2=0 $Y2=0
cc_454 N_Q_M1003_d N_VGND_c_833_n 0.00705989f $X=5.47 $Y=0.235 $X2=0 $Y2=0
cc_455 Q N_VGND_c_833_n 0.00994173f $X=5.645 $Y=0.425 $X2=0 $Y2=0
cc_456 N_VGND_c_833_n A_499_47# 0.0141891f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_457 N_VGND_c_833_n A_695_47# 0.00276139f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
