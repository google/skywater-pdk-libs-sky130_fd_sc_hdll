# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand2_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  15.64000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.440000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.505000 1.055000 14.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  4.440000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.055000 7.525000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  6.499000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.565000 1.495000 14.995000 1.665000 ;
        RECT  0.565000 1.665000  0.895000 2.465000 ;
        RECT  1.505000 1.665000  1.835000 2.465000 ;
        RECT  2.445000 1.665000  2.775000 2.465000 ;
        RECT  3.385000 1.665000  3.715000 2.465000 ;
        RECT  4.325000 1.665000  4.655000 2.465000 ;
        RECT  5.265000 1.665000  5.595000 2.465000 ;
        RECT  6.205000 1.665000  6.535000 2.465000 ;
        RECT  7.145000 1.665000  7.475000 2.465000 ;
        RECT  7.925000 1.055000  8.335000 1.495000 ;
        RECT  8.035000 0.635000 14.995000 0.885000 ;
        RECT  8.035000 0.885000  8.335000 1.055000 ;
        RECT  8.085000 1.665000  8.415000 2.465000 ;
        RECT  9.025000 1.665000  9.355000 2.465000 ;
        RECT  9.965000 1.665000 10.295000 2.465000 ;
        RECT 10.905000 1.665000 11.235000 2.465000 ;
        RECT 11.845000 1.665000 12.175000 2.465000 ;
        RECT 12.785000 1.665000 13.115000 2.465000 ;
        RECT 13.725000 1.665000 14.055000 2.465000 ;
        RECT 14.665000 1.665000 14.995000 2.465000 ;
        RECT 14.725000 0.885000 14.995000 1.055000 ;
        RECT 14.725000 1.055000 15.115000 1.325000 ;
        RECT 14.725000 1.325000 14.995000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.640000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.640000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.640000 0.085000 ;
      RECT  0.000000  2.635000 15.640000 2.805000 ;
      RECT  0.095000  0.255000  0.425000 0.715000 ;
      RECT  0.095000  0.715000  7.865000 0.885000 ;
      RECT  0.125000  1.495000  0.395000 2.635000 ;
      RECT  0.595000  0.085000  0.865000 0.545000 ;
      RECT  1.035000  0.255000  1.365000 0.715000 ;
      RECT  1.065000  1.835000  1.335000 2.635000 ;
      RECT  1.535000  0.085000  1.805000 0.545000 ;
      RECT  1.975000  0.255000  2.305000 0.715000 ;
      RECT  2.005000  1.835000  2.275000 2.635000 ;
      RECT  2.475000  0.085000  2.745000 0.545000 ;
      RECT  2.915000  0.255000  3.245000 0.715000 ;
      RECT  2.945000  1.835000  3.215000 2.635000 ;
      RECT  3.415000  0.085000  3.685000 0.545000 ;
      RECT  3.855000  0.255000  4.185000 0.715000 ;
      RECT  3.885000  1.835000  4.155000 2.635000 ;
      RECT  4.355000  0.085000  4.625000 0.545000 ;
      RECT  4.795000  0.255000  5.125000 0.715000 ;
      RECT  4.825000  1.835000  5.095000 2.635000 ;
      RECT  5.295000  0.085000  5.565000 0.545000 ;
      RECT  5.735000  0.255000  6.065000 0.715000 ;
      RECT  5.765000  1.835000  6.035000 2.635000 ;
      RECT  6.235000  0.085000  6.505000 0.545000 ;
      RECT  6.675000  0.255000  7.005000 0.715000 ;
      RECT  6.705000  1.835000  6.975000 2.635000 ;
      RECT  7.175000  0.085000  7.445000 0.545000 ;
      RECT  7.615000  0.255000 15.465000 0.465000 ;
      RECT  7.615000  0.465000  7.865000 0.715000 ;
      RECT  7.645000  1.835000  7.915000 2.635000 ;
      RECT  8.585000  1.835000  8.855000 2.635000 ;
      RECT  9.525000  1.835000  9.795000 2.635000 ;
      RECT 10.465000  1.835000 10.735000 2.635000 ;
      RECT 11.405000  1.835000 11.675000 2.635000 ;
      RECT 12.345000  1.835000 12.615000 2.635000 ;
      RECT 13.285000  1.835000 13.555000 2.635000 ;
      RECT 14.225000  1.835000 14.495000 2.635000 ;
      RECT 15.165000  1.495000 15.435000 2.635000 ;
      RECT 15.215000  0.465000 15.465000 0.885000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_16
