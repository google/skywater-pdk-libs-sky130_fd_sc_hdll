* NGSPICE file created from sky130_fd_sc_hdll__buf_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__buf_1 A VGND VNB VPB VPWR X
M1000 VPWR A a_27_47# VPB phighvt w=790000u l=180000u
+  ad=2.449e+11p pd=2.2e+06u as=2.133e+11p ps=2.12e+06u
M1001 X a_27_47# VPWR VPB phighvt w=790000u l=180000u
+  ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 VGND A a_27_47# VNB nshort w=520000u l=150000u
+  ad=1.768e+11p pd=1.72e+06u as=1.612e+11p ps=1.66e+06u
M1003 X a_27_47# VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
.ends

