* File: sky130_fd_sc_hdll__sdfrtp_2.pex.spice
* Created: Wed Sep  2 08:51:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%CLK 1 3 4 6 7 8 14
r31 14 15 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r32 12 14 32.6888 $w=3.76e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=1.202
+ $X2=0.495 $Y2=1.202
r33 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r34 7 8 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.315 $Y=1.53 $X2=0.315
+ $Y2=1.16
r35 4 15 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r37 1 14 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%A_27_47# 1 2 7 9 10 12 15 16 17 19 21 23
+ 24 26 28 29 31 34 38 39 45 47 48 49 54 56 57 58 59 60 67 69 73 74 77 79 81 91
c268 77 0 1.2887e-19 $X=0.94 $Y=1.16
c269 74 0 9.11424e-20 $X=9.32 $Y=1.11
c270 69 0 6.17614e-20 $X=9.32 $Y=1.19
c271 49 0 5.54695e-20 $X=0.71 $Y=1.88
c272 28 0 5.91276e-20 $X=9.185 $Y=1.89
c273 17 0 1.63397e-19 $X=6.43 $Y=1.32
c274 16 0 1.28412e-19 $X=5.72 $Y=0.745
r275 79 82 16.4869 $w=3.15e-07 $l=9e-08 $layer=POLY_cond $X=5.562 $Y=1.23
+ $X2=5.562 $Y2=1.32
r276 79 81 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=5.562 $Y=1.23
+ $X2=5.562 $Y2=1.065
r277 77 92 7.44021 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.867 $Y=1.16
+ $X2=0.867 $Y2=1.325
r278 77 91 8.29536 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.867 $Y=1.16
+ $X2=0.867 $Y2=0.995
r279 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r280 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.32
+ $Y=1.11 $X2=9.32 $Y2=1.11
r281 69 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.32 $Y=1.19
+ $X2=9.32 $Y2=1.19
r282 67 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.565
+ $Y=1.23 $X2=5.565 $Y2=1.23
r283 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.565 $Y=1.19
+ $X2=5.565 $Y2=1.19
r284 62 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.94 $Y=1.19
+ $X2=0.94 $Y2=1.19
r285 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.71 $Y=1.19
+ $X2=5.565 $Y2=1.19
r286 59 69 0.128299 $w=2.3e-07 $l=1.65e-07 $layer=MET1_cond $X=9.155 $Y=1.19
+ $X2=9.32 $Y2=1.19
r287 59 60 4.26361 $w=1.4e-07 $l=3.445e-06 $layer=MET1_cond $X=9.155 $Y=1.19
+ $X2=5.71 $Y2=1.19
r288 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.085 $Y=1.19
+ $X2=0.94 $Y2=1.19
r289 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.42 $Y=1.19
+ $X2=5.565 $Y2=1.19
r290 57 58 5.36509 $w=1.4e-07 $l=4.335e-06 $layer=MET1_cond $X=5.42 $Y=1.19
+ $X2=1.085 $Y2=1.19
r291 54 92 25.4279 $w=2.03e-07 $l=4.7e-07 $layer=LI1_cond $X=0.812 $Y=1.795
+ $X2=0.812 $Y2=1.325
r292 51 91 12.0416 $w=1.73e-07 $l=1.9e-07 $layer=LI1_cond $X=0.797 $Y=0.805
+ $X2=0.797 $Y2=0.995
r293 50 56 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.217 $Y2=1.88
r294 49 54 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=0.71 $Y=1.88
+ $X2=0.812 $Y2=1.795
r295 49 50 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.71 $Y=1.88
+ $X2=0.345 $Y2=1.88
r296 47 51 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=0.71 $Y=0.72
+ $X2=0.797 $Y2=0.805
r297 47 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.71 $Y=0.72
+ $X2=0.345 $Y2=0.72
r298 43 48 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=0.635
+ $X2=0.345 $Y2=0.72
r299 43 45 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.22 $Y=0.635
+ $X2=0.22 $Y2=0.51
r300 39 73 6.10776 $w=2.75e-07 $l=2.8e-08 $layer=POLY_cond $X=9.317 $Y=1.082
+ $X2=9.317 $Y2=1.11
r301 39 40 42.1909 $w=2.75e-07 $l=1.37e-07 $layer=POLY_cond $X=9.317 $Y=1.082
+ $X2=9.317 $Y2=0.945
r302 37 73 32.7201 $w=2.75e-07 $l=1.5e-07 $layer=POLY_cond $X=9.317 $Y=1.26
+ $X2=9.317 $Y2=1.11
r303 37 38 28.5635 $w=2.75e-07 $l=1.1e-07 $layer=POLY_cond $X=9.27 $Y=1.26
+ $X2=9.27 $Y2=1.37
r304 34 40 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.255 $Y=0.415
+ $X2=9.255 $Y2=0.945
r305 29 31 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.185 $Y=1.99
+ $X2=9.185 $Y2=2.275
r306 28 29 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=9.185 $Y=1.89 $X2=9.185
+ $Y2=1.99
r307 28 38 172.42 $w=2e-07 $l=5.2e-07 $layer=POLY_cond $X=9.185 $Y=1.89
+ $X2=9.185 $Y2=1.37
r308 24 26 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.53 $Y=1.99
+ $X2=6.53 $Y2=2.275
r309 23 24 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.53 $Y=1.89 $X2=6.53
+ $Y2=1.99
r310 22 23 164.131 $w=2e-07 $l=4.95e-07 $layer=POLY_cond $X=6.53 $Y=1.395
+ $X2=6.53 $Y2=1.89
r311 19 21 81.94 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.985 $Y=0.67
+ $X2=5.985 $Y2=0.415
r312 18 82 20.1192 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=5.72 $Y=1.32
+ $X2=5.562 $Y2=1.32
r313 17 22 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=6.43 $Y=1.32
+ $X2=6.53 $Y2=1.395
r314 17 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.43 $Y=1.32
+ $X2=5.72 $Y2=1.32
r315 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.91 $Y=0.745
+ $X2=5.985 $Y2=0.67
r316 15 16 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.91 $Y=0.745
+ $X2=5.72 $Y2=0.745
r317 13 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.645 $Y=0.82
+ $X2=5.72 $Y2=0.745
r318 13 81 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=5.645 $Y=0.82
+ $X2=5.645 $Y2=1.065
r319 10 76 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.965 $Y2=1.16
r320 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r321 7 76 48.1208 $w=2.95e-07 $l=2.57391e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.965 $Y2=1.16
r322 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.985
r323 2 56 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r324 1 45 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%A_331_66# 1 2 7 9 11 12 14 17 19 20 23 26
+ 28 30 31 33 34 35 38 46
c142 46 0 1.12841e-19 $X=2.62 $Y=1.165
c143 31 0 8.29887e-20 $X=2.73 $Y=1.09
r144 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.35
+ $Y=1.52 $X2=4.35 $Y2=1.52
r145 36 38 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=4.35 $Y=0.425
+ $X2=4.35 $Y2=1.52
r146 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.265 $Y=0.34
+ $X2=4.35 $Y2=0.425
r147 34 35 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=4.265 $Y=0.34
+ $X2=3.445 $Y2=0.34
r148 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.36 $Y=0.425
+ $X2=3.445 $Y2=0.34
r149 32 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.36 $Y=0.425
+ $X2=3.36 $Y2=0.995
r150 31 45 6.85038 $w=2.77e-07 $l=1.6895e-07 $layer=LI1_cond $X=2.73 $Y=1.09
+ $X2=2.602 $Y2=0.995
r151 30 33 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.275 $Y=1.09
+ $X2=3.36 $Y2=0.995
r152 30 31 31.8134 $w=1.88e-07 $l=5.45e-07 $layer=LI1_cond $X=3.275 $Y=1.09
+ $X2=2.73 $Y2=1.09
r153 29 46 18.2945 $w=3.8e-07 $l=1.25e-07 $layer=POLY_cond $X=2.62 $Y=1.29
+ $X2=2.62 $Y2=1.165
r154 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.29 $X2=2.645 $Y2=1.29
r155 26 28 28.2462 $w=2.53e-07 $l=6.25e-07 $layer=LI1_cond $X=2.602 $Y=1.915
+ $X2=2.602 $Y2=1.29
r156 25 45 1.23816 $w=2.55e-07 $l=1.9e-07 $layer=LI1_cond $X=2.602 $Y=1.185
+ $X2=2.602 $Y2=0.995
r157 25 28 4.74535 $w=2.53e-07 $l=1.05e-07 $layer=LI1_cond $X=2.602 $Y=1.185
+ $X2=2.602 $Y2=1.29
r158 21 26 23.2909 $w=1.68e-07 $l=3.57e-07 $layer=LI1_cond $X=2.245 $Y=2
+ $X2=2.602 $Y2=2
r159 21 23 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.245 $Y=2.085
+ $X2=2.245 $Y2=2.22
r160 19 45 16.6508 $w=2.77e-07 $l=4.17407e-07 $layer=LI1_cond $X=2.265 $Y=0.815
+ $X2=2.602 $Y2=0.995
r161 19 20 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.265 $Y=0.815
+ $X2=1.865 $Y2=0.815
r162 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.78 $Y=0.73
+ $X2=1.865 $Y2=0.815
r163 15 17 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.78 $Y=0.73
+ $X2=1.78 $Y2=0.56
r164 12 39 65.191 $w=2.89e-07 $l=3.82034e-07 $layer=POLY_cond $X=4.26 $Y=1.87
+ $X2=4.327 $Y2=1.52
r165 12 14 92.3833 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=4.26 $Y=1.87
+ $X2=4.26 $Y2=2.215
r166 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.08 $Y=1.09 $X2=3.08
+ $Y2=0.805
r167 8 46 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.81 $Y=1.165
+ $X2=2.62 $Y2=1.165
r168 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.005 $Y=1.165
+ $X2=3.08 $Y2=1.09
r169 7 8 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.005 $Y=1.165
+ $X2=2.81 $Y2=1.165
r170 2 23 600 $w=1.7e-07 $l=3.85357e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.945 $X2=2.295 $Y2=2.22
r171 1 17 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.33 $X2=1.78 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%D 1 3 6 8
r45 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.62 $X2=3.445 $Y2=1.62
r46 8 12 2.01209 $w=5.33e-07 $l=9e-08 $layer=LI1_cond $X=3.387 $Y=1.53 $X2=3.387
+ $Y2=1.62
r47 4 11 38.6899 $w=2.83e-07 $l=2.00237e-07 $layer=POLY_cond $X=3.54 $Y=1.455
+ $X2=3.462 $Y2=1.62
r48 4 6 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.54 $Y=1.455 $X2=3.54
+ $Y2=0.805
r49 1 11 48.9395 $w=2.83e-07 $l=2.74773e-07 $layer=POLY_cond $X=3.41 $Y=1.87
+ $X2=3.462 $Y2=1.62
r50 1 3 92.3833 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=3.41 $Y=1.87 $X2=3.41
+ $Y2=2.215
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%SCE 4 6 7 8 9 10 11 13 14 16 18 19 21 22
+ 23 24 26
c103 23 0 8.29887e-20 $X=2.04 $Y=1.31
c104 14 0 5.48891e-20 $X=2.9 $Y=1.71
r105 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.805
+ $Y=1.31 $X2=1.805 $Y2=1.31
r106 26 30 5.58377 $w=5.79e-07 $l=2.65e-07 $layer=LI1_cond $X=2.07 $Y=1.407
+ $X2=1.805 $Y2=1.407
r107 22 29 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.965 $Y=1.31
+ $X2=1.805 $Y2=1.31
r108 22 23 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.965 $Y=1.31
+ $X2=2.04 $Y2=1.31
r109 19 21 27.474 $w=5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.245 $Y=0.255
+ $X2=4.245 $Y2=0.54
r110 16 18 92.3833 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=3 $Y=1.87 $X2=3
+ $Y2=2.215
r111 15 24 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=2.63 $Y=1.71 $X2=2.53
+ $Y2=1.71
r112 14 16 27.2212 $w=1.5e-07 $l=2.03961e-07 $layer=POLY_cond $X=2.9 $Y=1.71
+ $X2=3 $Y2=1.87
r113 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.9 $Y=1.71
+ $X2=2.63 $Y2=1.71
r114 11 24 53.8601 $w=2e-07 $l=1.6e-07 $layer=POLY_cond $X=2.53 $Y=1.87 $X2=2.53
+ $Y2=1.71
r115 11 13 92.3833 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=2.53 $Y=1.87
+ $X2=2.53 $Y2=2.215
r116 9 24 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=2.43 $Y=1.71 $X2=2.53
+ $Y2=1.71
r117 9 10 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.43 $Y=1.71
+ $X2=2.115 $Y2=1.71
r118 7 19 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.995 $Y=0.18
+ $X2=4.245 $Y2=0.255
r119 7 8 964 $w=1.5e-07 $l=1.88e-06 $layer=POLY_cond $X=3.995 $Y=0.18 $X2=2.115
+ $Y2=0.18
r120 6 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.04 $Y=1.635
+ $X2=2.115 $Y2=1.71
r121 5 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.475
+ $X2=2.04 $Y2=1.31
r122 5 6 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.04 $Y=1.475
+ $X2=2.04 $Y2=1.635
r123 2 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.145
+ $X2=2.04 $Y2=1.31
r124 2 4 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=2.04 $Y=1.145
+ $X2=2.04 $Y2=0.54
r125 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.04 $Y=0.255
+ $X2=2.115 $Y2=0.18
r126 1 4 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.04 $Y=0.255
+ $X2=2.04 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%SCD 1 3 6 8 14
c39 8 0 1.28412e-19 $X=4.745 $Y=1.445
r40 8 14 0.0616162 $w=9.88e-07 $l=5e-09 $layer=LI1_cond $X=4.835 $Y=1.205
+ $X2=4.83 $Y2=1.205
r41 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.87
+ $Y=1.535 $X2=4.87 $Y2=1.535
r42 4 11 34.2818 $w=2.92e-07 $l=2.0106e-07 $layer=POLY_cond $X=4.955 $Y=1.37
+ $X2=4.875 $Y2=1.535
r43 4 6 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=4.955 $Y=1.37
+ $X2=4.955 $Y2=0.54
r44 1 11 62.3435 $w=2.92e-07 $l=3.68341e-07 $layer=POLY_cond $X=4.805 $Y=1.87
+ $X2=4.875 $Y2=1.535
r45 1 3 92.3833 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=4.805 $Y=1.87
+ $X2=4.805 $Y2=2.215
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%A_213_47# 1 2 7 9 10 12 13 15 16 18 23 25
+ 30 31 33 34 36 39 40 41 46 47 48 49 52 58 63 66 74 81
c253 66 0 3.82543e-21 $X=6.535 $Y=0.87
c254 46 0 2.76238e-19 $X=5.89 $Y=1.87
c255 41 0 5.99032e-20 $X=9.315 $Y=1.58
r256 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.63
+ $Y=1.745 $X2=9.63 $Y2=1.745
r257 63 81 7.18001 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.97 $Y=1.74
+ $X2=5.97 $Y2=1.575
r258 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.905
+ $Y=1.74 $X2=5.905 $Y2=1.74
r259 58 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.65 $Y=1.87
+ $X2=9.65 $Y2=1.87
r260 55 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.035 $Y=1.87
+ $X2=6.035 $Y2=1.87
r261 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.22 $Y=1.87
+ $X2=1.22 $Y2=1.87
r262 49 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.18 $Y=1.87
+ $X2=6.035 $Y2=1.87
r263 48 58 0.118675 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=9.5 $Y=1.87
+ $X2=9.65 $Y2=1.87
r264 48 49 4.1089 $w=1.4e-07 $l=3.32e-06 $layer=MET1_cond $X=9.5 $Y=1.87
+ $X2=6.18 $Y2=1.87
r265 47 51 0.118675 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=1.37 $Y=1.87
+ $X2=1.22 $Y2=1.87
r266 46 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.89 $Y=1.87
+ $X2=6.035 $Y2=1.87
r267 46 47 5.59405 $w=1.4e-07 $l=4.52e-06 $layer=MET1_cond $X=5.89 $Y=1.87
+ $X2=1.37 $Y2=1.87
r268 44 74 7.22718 $w=2.93e-07 $l=1.85e-07 $layer=LI1_cond $X=9.445 $Y=1.807
+ $X2=9.63 $Y2=1.807
r269 41 44 10.0617 $w=2.58e-07 $l=2.27e-07 $layer=LI1_cond $X=9.315 $Y=1.58
+ $X2=9.315 $Y2=1.807
r270 39 52 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.25 $Y=1.845
+ $X2=1.25 $Y2=1.87
r271 39 40 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.25 $Y=1.845
+ $X2=1.25 $Y2=1.73
r272 38 40 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=1.28 $Y=0.675
+ $X2=1.28 $Y2=1.73
r273 36 38 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=0.51
+ $X2=1.24 $Y2=0.675
r274 33 41 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.185 $Y=1.58
+ $X2=9.315 $Y2=1.58
r275 33 34 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.185 $Y=1.58
+ $X2=8.97 $Y2=1.58
r276 31 68 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=8.835 $Y=0.87
+ $X2=8.71 $Y2=0.87
r277 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.835
+ $Y=0.87 $X2=8.835 $Y2=0.87
r278 28 34 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=8.84 $Y=1.495
+ $X2=8.97 $Y2=1.58
r279 28 30 27.703 $w=2.58e-07 $l=6.25e-07 $layer=LI1_cond $X=8.84 $Y=1.495
+ $X2=8.84 $Y2=0.87
r280 26 66 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=6.425 $Y=0.87
+ $X2=6.535 $Y2=0.87
r281 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.425
+ $Y=0.87 $X2=6.425 $Y2=0.87
r282 23 25 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.12 $Y=0.87
+ $X2=6.425 $Y2=0.87
r283 21 23 7.17723 $w=3.3e-07 $l=2.13014e-07 $layer=LI1_cond $X=6.01 $Y=1.035
+ $X2=6.12 $Y2=0.87
r284 21 81 28.2872 $w=2.18e-07 $l=5.4e-07 $layer=LI1_cond $X=6.01 $Y=1.035
+ $X2=6.01 $Y2=1.575
r285 16 73 47.186 $w=2.97e-07 $l=2.4995e-07 $layer=POLY_cond $X=9.665 $Y=1.99
+ $X2=9.655 $Y2=1.745
r286 16 18 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.665 $Y=1.99
+ $X2=9.665 $Y2=2.275
r287 13 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.71 $Y=0.705
+ $X2=8.71 $Y2=0.87
r288 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.71 $Y=0.705
+ $X2=8.71 $Y2=0.415
r289 10 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.535 $Y=0.705
+ $X2=6.535 $Y2=0.87
r290 10 12 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.535 $Y=0.705
+ $X2=6.535 $Y2=0.415
r291 7 62 46.5577 $w=3.26e-07 $l=2.54951e-07 $layer=POLY_cond $X=5.92 $Y=1.99
+ $X2=5.93 $Y2=1.74
r292 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.92 $Y=1.99
+ $X2=5.92 $Y2=2.275
r293 2 52 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.485 $X2=1.22 $Y2=1.96
r294 1 36 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%A_1380_303# 1 2 7 9 12 14 20 23 27 30 33
+ 34 35
c108 35 0 5.91276e-20 $X=8.385 $Y=1.595
c109 33 0 1.46876e-19 $X=8.385 $Y=0.835
c110 1 0 1.64006e-19 $X=8.31 $Y=0.235
r111 34 36 8.92214 $w=3.08e-07 $l=2.4e-07 $layer=LI1_cond $X=8.385 $Y=1.68
+ $X2=8.385 $Y2=1.92
r112 34 35 5.49324 $w=3.08e-07 $l=8.5e-08 $layer=LI1_cond $X=8.385 $Y=1.68
+ $X2=8.385 $Y2=1.595
r113 33 35 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=8.455 $Y=0.835
+ $X2=8.455 $Y2=1.595
r114 30 32 3.00288 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=0.36
+ $X2=8.42 $Y2=0.445
r115 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.9 $Y=2.005
+ $X2=8.9 $Y2=2.3
r116 24 36 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.54 $Y=1.92
+ $X2=8.385 $Y2=1.92
r117 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.815 $Y=1.92
+ $X2=8.9 $Y2=2.005
r118 23 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.815 $Y=1.92
+ $X2=8.54 $Y2=1.92
r119 20 33 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=8.385 $Y=0.68
+ $X2=8.385 $Y2=0.835
r120 20 32 8.73626 $w=3.08e-07 $l=2.35e-07 $layer=LI1_cond $X=8.385 $Y=0.68
+ $X2=8.385 $Y2=0.445
r121 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.125
+ $Y=1.68 $X2=7.125 $Y2=1.68
r122 14 34 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.23 $Y=1.68
+ $X2=8.385 $Y2=1.68
r123 14 16 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=8.23 $Y=1.68
+ $X2=7.125 $Y2=1.68
r124 10 17 38.7839 $w=3.5e-07 $l=1.83916e-07 $layer=POLY_cond $X=7.065 $Y=1.515
+ $X2=7.105 $Y2=1.68
r125 10 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=7.065 $Y=1.515
+ $X2=7.065 $Y2=0.445
r126 7 17 54.0257 $w=3.5e-07 $l=3.58678e-07 $layer=POLY_cond $X=7 $Y=1.99
+ $X2=7.105 $Y2=1.68
r127 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7 $Y=1.99 $X2=7
+ $Y2=2.275
r128 2 27 600 $w=1.7e-07 $l=7.26137e-07 $layer=licon1_PDIFF $count=1 $X=8.75
+ $Y=1.645 $X2=8.9 $Y2=2.3
r129 1 30 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=8.31
+ $Y=0.235 $X2=8.445 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%RESET_B 3 5 6 8 11 14 15 17 18 21 24 27
+ 29 30 31 34 36 45
c157 45 0 4.8947e-20 $X=11.225 $Y=0.85
c158 34 0 1.46876e-19 $X=7.535 $Y=0.96
c159 29 0 1.64006e-19 $X=11.08 $Y=0.85
c160 21 0 8.70495e-20 $X=10.77 $Y=1.15
c161 18 0 1.48828e-19 $X=11.065 $Y=1.17
c162 5 0 1.10071e-19 $X=7.62 $Y=1.89
r163 34 37 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.56 $Y=0.96
+ $X2=7.56 $Y2=1.125
r164 34 36 53.3639 $w=3.2e-07 $l=2.05e-07 $layer=POLY_cond $X=7.56 $Y=0.96
+ $X2=7.56 $Y2=0.755
r165 31 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.225 $Y=0.85
+ $X2=11.225 $Y2=0.85
r166 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.08 $Y=0.85
+ $X2=11.225 $Y2=0.85
r167 29 30 3.93564 $w=1.4e-07 $l=3.18e-06 $layer=MET1_cond $X=11.08 $Y=0.85
+ $X2=7.9 $Y2=0.85
r168 27 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.535
+ $Y=0.96 $X2=7.535 $Y2=0.96
r169 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.7 $Y=0.85
+ $X2=7.7 $Y2=0.85
r170 24 30 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=7.785 $Y=0.85
+ $X2=7.9 $Y2=0.85
r171 24 26 0.0545364 $w=2.3e-07 $l=8.5e-08 $layer=MET1_cond $X=7.785 $Y=0.85
+ $X2=7.7 $Y2=0.85
r172 23 45 8.12378 $w=3.03e-07 $l=2.15e-07 $layer=LI1_cond $X=11.217 $Y=1.065
+ $X2=11.217 $Y2=0.85
r173 21 40 39.5599 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=10.787 $Y=1.15
+ $X2=10.787 $Y2=1.315
r174 21 39 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=10.787 $Y=1.15
+ $X2=10.787 $Y2=0.985
r175 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.77
+ $Y=1.15 $X2=10.77 $Y2=1.15
r176 18 23 7.12258 $w=2.1e-07 $l=1.97646e-07 $layer=LI1_cond $X=11.065 $Y=1.17
+ $X2=11.217 $Y2=1.065
r177 18 20 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=11.065 $Y=1.17
+ $X2=10.77 $Y2=1.17
r178 15 17 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.735 $Y=1.99
+ $X2=10.735 $Y2=2.275
r179 14 15 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=10.735 $Y=1.89
+ $X2=10.735 $Y2=1.99
r180 14 40 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=10.735 $Y=1.89
+ $X2=10.735 $Y2=1.315
r181 11 39 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=10.71 $Y=0.445
+ $X2=10.71 $Y2=0.985
r182 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.62 $Y=1.99
+ $X2=7.62 $Y2=2.275
r183 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.62 $Y=1.89 $X2=7.62
+ $Y2=1.99
r184 5 37 253.657 $w=2e-07 $l=7.65e-07 $layer=POLY_cond $X=7.62 $Y=1.89 $X2=7.62
+ $Y2=1.125
r185 3 36 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.475 $Y=0.445
+ $X2=7.475 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%A_1202_413# 1 2 9 11 13 15 16 22 23 25 26
+ 29 30 32 34 35
c139 34 0 1.10071e-19 $X=8.065 $Y=1.17
c140 32 0 1.87801e-19 $X=6.925 $Y=1.3
c141 11 0 3.66493e-20 $X=8.57 $Y=1.495
r142 35 40 51.3607 $w=3.05e-07 $l=3.25e-07 $layer=POLY_cond $X=8.12 $Y=1.17
+ $X2=8.12 $Y2=1.495
r143 34 37 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=8.065 $Y=1.17
+ $X2=8.065 $Y2=1.3
r144 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.065
+ $Y=1.17 $X2=8.065 $Y2=1.17
r145 29 30 9.47152 $w=3.63e-07 $l=1.95e-07 $layer=LI1_cond $X=6.277 $Y=2.33
+ $X2=6.277 $Y2=2.135
r146 27 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=1.3
+ $X2=6.925 $Y2=1.3
r147 26 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=1.3
+ $X2=8.065 $Y2=1.3
r148 26 27 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=7.98 $Y=1.3
+ $X2=7.01 $Y2=1.3
r149 25 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=1.215
+ $X2=6.925 $Y2=1.3
r150 24 25 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.925 $Y=0.475
+ $X2=6.925 $Y2=1.215
r151 22 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=1.3
+ $X2=6.925 $Y2=1.3
r152 22 23 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.84 $Y=1.3
+ $X2=6.46 $Y2=1.3
r153 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=1.385
+ $X2=6.46 $Y2=1.3
r154 20 30 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=6.375 $Y=1.385
+ $X2=6.375 $Y2=2.135
r155 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.84 $Y=0.39
+ $X2=6.925 $Y2=0.475
r156 16 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.84 $Y=0.39
+ $X2=6.275 $Y2=0.39
r157 13 15 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.66 $Y=1.57
+ $X2=8.66 $Y2=2.065
r158 12 40 19.3576 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.31 $Y=1.495
+ $X2=8.12 $Y2=1.495
r159 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.57 $Y=1.495
+ $X2=8.66 $Y2=1.57
r160 11 12 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=8.57 $Y=1.495
+ $X2=8.31 $Y2=1.495
r161 7 35 38.5368 $w=3.05e-07 $l=2.14942e-07 $layer=POLY_cond $X=8.235 $Y=1.005
+ $X2=8.12 $Y2=1.17
r162 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=8.235 $Y=1.005
+ $X2=8.235 $Y2=0.555
r163 2 29 600 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=1 $X=6.01
+ $Y=2.065 $X2=6.295 $Y2=2.33
r164 1 18 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=6.06
+ $Y=0.235 $X2=6.275 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%A_1972_21# 1 2 9 12 13 15 16 18 19 21 22
+ 24 25 27 30 33 34 36 37 38 43 45 46 48 50 53 56 58 63
c155 63 0 1.97775e-19 $X=12.845 $Y=1.202
c156 58 0 8.39514e-20 $X=10.175 $Y=0.98
c157 33 0 2.50234e-20 $X=10.56 $Y=0.78
c158 30 0 8.70495e-20 $X=10.235 $Y=0.98
c159 12 0 7.19093e-21 $X=10.175 $Y=1.89
r160 63 64 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=12.845 $Y=1.202
+ $X2=12.87 $Y2=1.202
r161 62 63 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=12.4 $Y=1.202
+ $X2=12.845 $Y2=1.202
r162 61 62 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=12.375 $Y=1.202
+ $X2=12.4 $Y2=1.202
r163 54 61 29.7123 $w=3.65e-07 $l=2.25e-07 $layer=POLY_cond $X=12.15 $Y=1.202
+ $X2=12.375 $Y2=1.202
r164 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.15
+ $Y=1.16 $X2=12.15 $Y2=1.16
r165 51 56 0.850971 $w=3.3e-07 $l=8.8e-08 $layer=LI1_cond $X=11.735 $Y=1.16
+ $X2=11.647 $Y2=1.16
r166 51 53 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=11.735 $Y=1.16
+ $X2=12.15 $Y2=1.16
r167 49 56 8.52281 $w=1.72e-07 $l=1.65997e-07 $layer=LI1_cond $X=11.645 $Y=1.325
+ $X2=11.647 $Y2=1.16
r168 49 50 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.645 $Y=1.325
+ $X2=11.645 $Y2=1.915
r169 48 56 8.52281 $w=1.72e-07 $l=1.65e-07 $layer=LI1_cond $X=11.647 $Y=0.995
+ $X2=11.647 $Y2=1.16
r170 47 48 33.5896 $w=1.73e-07 $l=5.3e-07 $layer=LI1_cond $X=11.647 $Y=0.465
+ $X2=11.647 $Y2=0.995
r171 45 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.56 $Y=2
+ $X2=11.645 $Y2=1.915
r172 45 46 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=11.56 $Y=2
+ $X2=11.08 $Y2=2
r173 41 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.995 $Y=2.085
+ $X2=11.08 $Y2=2
r174 41 43 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.995 $Y=2.085
+ $X2=10.995 $Y2=2.21
r175 38 40 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=10.73 $Y=0.38
+ $X2=11.445 $Y2=0.38
r176 37 47 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=11.56 $Y=0.38
+ $X2=11.647 $Y2=0.465
r177 37 40 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=11.56 $Y=0.38
+ $X2=11.445 $Y2=0.38
r178 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.645 $Y=0.465
+ $X2=10.73 $Y2=0.38
r179 35 36 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=10.645 $Y=0.465
+ $X2=10.645 $Y2=0.695
r180 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.56 $Y=0.78
+ $X2=10.645 $Y2=0.695
r181 33 34 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.56 $Y=0.78
+ $X2=10.37 $Y2=0.78
r182 31 58 11.1231 $w=2.6e-07 $l=6e-08 $layer=POLY_cond $X=10.235 $Y=0.98
+ $X2=10.175 $Y2=0.98
r183 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.235
+ $Y=0.98 $X2=10.235 $Y2=0.98
r184 28 34 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=10.26 $Y=0.865
+ $X2=10.37 $Y2=0.78
r185 28 30 6.02413 $w=2.18e-07 $l=1.15e-07 $layer=LI1_cond $X=10.26 $Y=0.865
+ $X2=10.26 $Y2=0.98
r186 25 64 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.87 $Y=0.995
+ $X2=12.87 $Y2=1.202
r187 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.87 $Y=0.995
+ $X2=12.87 $Y2=0.56
r188 22 63 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.845 $Y=1.41
+ $X2=12.845 $Y2=1.202
r189 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.845 $Y=1.41
+ $X2=12.845 $Y2=1.985
r190 19 62 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.4 $Y=0.995
+ $X2=12.4 $Y2=1.202
r191 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.4 $Y=0.995
+ $X2=12.4 $Y2=0.56
r192 16 61 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.375 $Y=1.41
+ $X2=12.375 $Y2=1.202
r193 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.375 $Y=1.41
+ $X2=12.375 $Y2=1.985
r194 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.175 $Y=1.99
+ $X2=10.175 $Y2=2.275
r195 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=10.175 $Y=1.89
+ $X2=10.175 $Y2=1.99
r196 11 58 8.99251 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.175 $Y=1.145
+ $X2=10.175 $Y2=0.98
r197 11 12 247.025 $w=2e-07 $l=7.45e-07 $layer=POLY_cond $X=10.175 $Y=1.145
+ $X2=10.175 $Y2=1.89
r198 7 58 44.4923 $w=2.6e-07 $l=3.11769e-07 $layer=POLY_cond $X=9.935 $Y=0.815
+ $X2=10.175 $Y2=0.98
r199 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.935 $Y=0.815
+ $X2=9.935 $Y2=0.445
r200 2 43 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=10.825
+ $Y=2.065 $X2=10.995 $Y2=2.21
r201 1 40 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=11.265
+ $Y=0.235 $X2=11.445 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%A_1757_47# 1 2 9 10 12 14 15 16 17 21 26
+ 28 29 31
c112 28 0 2.32539e-20 $X=10.127 $Y=2.125
c113 14 0 2.50234e-20 $X=11.275 $Y=1.495
r114 34 35 15.507 $w=2.73e-07 $l=3.47e-07 $layer=LI1_cond $X=9.78 $Y=1.485
+ $X2=10.127 $Y2=1.485
r115 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.18
+ $Y=1.66 $X2=11.18 $Y2=1.66
r116 29 35 8.78748 $w=2.73e-07 $l=2.41402e-07 $layer=LI1_cond $X=10.285 $Y=1.66
+ $X2=10.127 $Y2=1.485
r117 29 31 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=10.285 $Y=1.66
+ $X2=11.18 $Y2=1.66
r118 27 35 3.3616 $w=1.75e-07 $l=2.6e-07 $layer=LI1_cond $X=10.127 $Y=1.745
+ $X2=10.127 $Y2=1.485
r119 27 28 24.0831 $w=1.73e-07 $l=3.8e-07 $layer=LI1_cond $X=10.127 $Y=1.745
+ $X2=10.127 $Y2=2.125
r120 26 34 2.00371 $w=2.2e-07 $l=1.7e-07 $layer=LI1_cond $X=9.78 $Y=1.315
+ $X2=9.78 $Y2=1.485
r121 25 26 40.8593 $w=2.18e-07 $l=7.8e-07 $layer=LI1_cond $X=9.78 $Y=0.535
+ $X2=9.78 $Y2=1.315
r122 21 28 7.76859 $w=3.4e-07 $l=2.09022e-07 $layer=LI1_cond $X=10.04 $Y=2.295
+ $X2=10.127 $Y2=2.125
r123 21 23 20.6762 $w=3.38e-07 $l=6.1e-07 $layer=LI1_cond $X=10.04 $Y=2.295
+ $X2=9.43 $Y2=2.295
r124 17 25 6.94494 $w=2.8e-07 $l=1.87083e-07 $layer=LI1_cond $X=9.67 $Y=0.395
+ $X2=9.78 $Y2=0.535
r125 17 19 29.84 $w=2.78e-07 $l=7.25e-07 $layer=LI1_cond $X=9.67 $Y=0.395
+ $X2=8.945 $Y2=0.395
r126 15 16 44.0828 $w=2e-07 $l=1.2e-07 $layer=POLY_cond $X=11.245 $Y=0.73
+ $X2=11.245 $Y2=0.85
r127 14 32 32.2196 $w=2.86e-07 $l=1.94808e-07 $layer=POLY_cond $X=11.275
+ $Y=1.495 $X2=11.21 $Y2=1.66
r128 14 16 213.867 $w=2e-07 $l=6.45e-07 $layer=POLY_cond $X=11.275 $Y=1.495
+ $X2=11.275 $Y2=0.85
r129 10 32 62.2041 $w=2.86e-07 $l=3.42272e-07 $layer=POLY_cond $X=11.235 $Y=1.99
+ $X2=11.21 $Y2=1.66
r130 10 12 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=11.235 $Y=1.99
+ $X2=11.235 $Y2=2.275
r131 9 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.19 $Y=0.445
+ $X2=11.19 $Y2=0.73
r132 2 23 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=9.275
+ $Y=2.065 $X2=9.43 $Y2=2.335
r133 1 19 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=8.785
+ $Y=0.235 $X2=8.945 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 48
+ 52 56 58 63 64 66 67 69 72 75 76 77 79 103 111 116 122 125 128 135 139 142
c189 139 0 1.26055e-19 $X=13.11 $Y=2.72
c190 66 0 1.00946e-19 $X=4.855 $Y=2.72
c191 63 0 5.54695e-20 $X=2.6 $Y=2.72
r192 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r193 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r194 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r195 128 131 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=11.445 $Y=2.34
+ $X2=11.445 $Y2=2.72
r196 125 126 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r197 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r198 120 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r199 120 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r200 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r201 117 135 10.2049 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=12.33 $Y=2.72
+ $X2=12.117 $Y2=2.72
r202 117 119 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.33 $Y=2.72
+ $X2=12.65 $Y2=2.72
r203 116 138 4.04153 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=12.995 $Y=2.72
+ $X2=13.167 $Y2=2.72
r204 116 119 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.995 $Y=2.72
+ $X2=12.65 $Y2=2.72
r205 115 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r206 115 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=11.27 $Y2=2.72
r207 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r208 112 131 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.635 $Y=2.72
+ $X2=11.445 $Y2=2.72
r209 112 114 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=11.635 $Y=2.72
+ $X2=11.73 $Y2=2.72
r210 111 135 10.2049 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=11.905 $Y=2.72
+ $X2=12.117 $Y2=2.72
r211 111 114 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=11.905 $Y=2.72
+ $X2=11.73 $Y2=2.72
r212 110 132 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r213 110 126 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=8.51 $Y2=2.72
r214 109 110 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r215 107 125 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.57 $Y=2.72
+ $X2=8.36 $Y2=2.72
r216 107 109 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=8.57 $Y=2.72
+ $X2=10.35 $Y2=2.72
r217 106 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r218 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r219 103 125 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.15 $Y=2.72
+ $X2=8.36 $Y2=2.72
r220 103 105 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=8.15 $Y=2.72
+ $X2=8.05 $Y2=2.72
r221 102 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r222 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r223 99 102 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=7.13 $Y2=2.72
r224 98 101 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=7.13 $Y2=2.72
r225 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r226 96 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r227 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r228 93 96 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.83 $Y2=2.72
r229 92 95 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=4.83 $Y2=2.72
r230 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r231 90 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r232 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r233 87 90 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r234 87 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r235 86 89 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r236 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r237 84 122 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=2.72
+ $X2=0.72 $Y2=2.72
r238 84 86 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.91 $Y=2.72
+ $X2=1.15 $Y2=2.72
r239 81 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r240 79 122 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.53 $Y=2.72
+ $X2=0.72 $Y2=2.72
r241 79 81 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.53 $Y=2.72 $X2=0.23
+ $Y2=2.72
r242 77 123 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r243 77 142 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r244 75 109 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.35 $Y2=2.72
r245 75 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.54 $Y2=2.72
r246 73 105 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=7.465 $Y=2.72
+ $X2=8.05 $Y2=2.72
r247 72 101 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=7.135 $Y=2.72
+ $X2=7.13 $Y2=2.72
r248 71 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.3 $Y=2.72
+ $X2=7.465 $Y2=2.72
r249 71 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.3 $Y=2.72
+ $X2=7.135 $Y2=2.72
r250 69 71 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=7.3 $Y=2.44 $X2=7.3
+ $Y2=2.72
r251 66 95 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.855 $Y=2.72
+ $X2=4.83 $Y2=2.72
r252 66 67 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.855 $Y=2.72
+ $X2=5.03 $Y2=2.72
r253 65 98 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=2.72
+ $X2=5.29 $Y2=2.72
r254 65 67 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.205 $Y=2.72
+ $X2=5.03 $Y2=2.72
r255 63 89 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.6 $Y=2.72 $X2=2.53
+ $Y2=2.72
r256 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=2.72
+ $X2=2.765 $Y2=2.72
r257 62 92 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.93 $Y=2.72 $X2=2.99
+ $Y2=2.72
r258 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=2.72
+ $X2=2.765 $Y2=2.72
r259 58 61 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=13.12 $Y=1.66
+ $X2=13.12 $Y2=2.34
r260 56 138 3.10164 $w=2.5e-07 $l=1.05924e-07 $layer=LI1_cond $X=13.12 $Y=2.635
+ $X2=13.167 $Y2=2.72
r261 56 61 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=13.12 $Y=2.635
+ $X2=13.12 $Y2=2.34
r262 52 55 18.4391 $w=4.23e-07 $l=6.8e-07 $layer=LI1_cond $X=12.117 $Y=1.66
+ $X2=12.117 $Y2=2.34
r263 50 135 1.63918 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=12.117 $Y=2.635
+ $X2=12.117 $Y2=2.72
r264 50 55 7.99931 $w=4.23e-07 $l=2.95e-07 $layer=LI1_cond $X=12.117 $Y=2.635
+ $X2=12.117 $Y2=2.34
r265 49 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.665 $Y=2.72
+ $X2=10.54 $Y2=2.72
r266 48 131 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.255 $Y=2.72
+ $X2=11.445 $Y2=2.72
r267 48 49 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.255 $Y=2.72
+ $X2=10.665 $Y2=2.72
r268 44 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.54 $Y=2.635
+ $X2=10.54 $Y2=2.72
r269 44 46 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=10.54 $Y=2.635
+ $X2=10.54 $Y2=2.36
r270 40 125 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=2.635
+ $X2=8.36 $Y2=2.72
r271 40 42 8.09454 $w=4.18e-07 $l=2.95e-07 $layer=LI1_cond $X=8.36 $Y=2.635
+ $X2=8.36 $Y2=2.34
r272 36 67 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=2.635
+ $X2=5.03 $Y2=2.72
r273 36 38 9.05491 $w=3.48e-07 $l=2.75e-07 $layer=LI1_cond $X=5.03 $Y=2.635
+ $X2=5.03 $Y2=2.36
r274 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=2.635
+ $X2=2.765 $Y2=2.72
r275 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.765 $Y=2.635
+ $X2=2.765 $Y2=2.34
r276 28 122 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.72
r277 28 30 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.22
r278 9 61 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.935
+ $Y=1.485 $X2=13.08 $Y2=2.34
r279 9 58 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.935
+ $Y=1.485 $X2=13.08 $Y2=1.66
r280 8 55 400 $w=1.7e-07 $l=9.63159e-07 $layer=licon1_PDIFF $count=1 $X=11.865
+ $Y=1.485 $X2=12.095 $Y2=2.34
r281 8 52 400 $w=1.7e-07 $l=3.05205e-07 $layer=licon1_PDIFF $count=1 $X=11.865
+ $Y=1.485 $X2=12.095 $Y2=1.66
r282 7 128 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=11.325
+ $Y=2.065 $X2=11.47 $Y2=2.34
r283 6 46 600 $w=1.7e-07 $l=3.95411e-07 $layer=licon1_PDIFF $count=1 $X=10.265
+ $Y=2.065 $X2=10.5 $Y2=2.36
r284 5 42 600 $w=1.7e-07 $l=7.77592e-07 $layer=licon1_PDIFF $count=1 $X=8.25
+ $Y=1.645 $X2=8.425 $Y2=2.34
r285 4 69 600 $w=1.7e-07 $l=4.68375e-07 $layer=licon1_PDIFF $count=1 $X=7.09
+ $Y=2.065 $X2=7.3 $Y2=2.44
r286 3 38 600 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.945 $X2=5.04 $Y2=2.36
r287 2 34 600 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=1 $X=2.62
+ $Y=1.945 $X2=2.765 $Y2=2.34
r288 1 30 600 $w=1.7e-07 $l=8.11064e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.745 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%A_700_389# 1 2 3 4 14 17 19 22 23 24 26
+ 30 32 39
c97 32 0 2.74431e-19 $X=3.957 $Y=2.02
c98 26 0 3.82543e-21 $X=5.635 $Y=0.715
r99 36 39 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.635 $Y=0.42
+ $X2=5.725 $Y2=0.42
r100 28 30 5.96389 $w=3.98e-07 $l=2.07e-07 $layer=LI1_cond $X=3.75 $Y=0.875
+ $X2=3.957 $Y2=0.875
r101 25 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=0.505
+ $X2=5.635 $Y2=0.42
r102 25 26 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.635 $Y=0.505
+ $X2=5.635 $Y2=0.715
r103 23 26 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.55 $Y=0.805
+ $X2=5.635 $Y2=0.715
r104 23 24 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=5.55 $Y=0.805
+ $X2=5.31 $Y2=0.805
r105 22 35 20.7085 $w=2.71e-07 $l=5.71489e-07 $layer=LI1_cond $X=5.225 $Y=1.935
+ $X2=5.685 $Y2=2.185
r106 21 24 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.225 $Y=0.895
+ $X2=5.31 $Y2=0.805
r107 21 22 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=5.225 $Y=0.895
+ $X2=5.225 $Y2=1.935
r108 20 32 1.39518 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=4.045 $Y=2.02
+ $X2=3.957 $Y2=2.02
r109 19 22 5.51241 $w=2.71e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.14 $Y=2.02
+ $X2=5.225 $Y2=1.935
r110 19 20 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=5.14 $Y=2.02
+ $X2=4.045 $Y2=2.02
r111 15 32 5.10356 $w=1.72e-07 $l=8.59942e-08 $layer=LI1_cond $X=3.955 $Y=2.105
+ $X2=3.957 $Y2=2.02
r112 15 17 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.955 $Y=2.105
+ $X2=3.955 $Y2=2.3
r113 14 32 5.10356 $w=1.72e-07 $l=8.5e-08 $layer=LI1_cond $X=3.957 $Y=1.935
+ $X2=3.957 $Y2=2.02
r114 13 30 5.61783 $w=1.75e-07 $l=2e-07 $layer=LI1_cond $X=3.957 $Y=1.075
+ $X2=3.957 $Y2=0.875
r115 13 14 54.5039 $w=1.73e-07 $l=8.6e-07 $layer=LI1_cond $X=3.957 $Y=1.075
+ $X2=3.957 $Y2=1.935
r116 4 35 600 $w=1.7e-07 $l=3.16307e-07 $layer=licon1_PDIFF $count=1 $X=5.455
+ $Y=2.065 $X2=5.685 $Y2=2.27
r117 3 17 600 $w=1.7e-07 $l=6.07083e-07 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.945 $X2=3.955 $Y2=2.3
r118 2 39 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=5.6
+ $Y=0.235 $X2=5.725 $Y2=0.42
r119 1 28 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.595 $X2=3.75 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%A_1324_413# 1 2 7 9 14
c31 9 0 1.87801e-19 $X=6.765 $Y=2.02
r32 14 17 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.855 $Y=2.02
+ $X2=7.855 $Y2=2.21
r33 9 12 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.765 $Y=2.02
+ $X2=6.765 $Y2=2.21
r34 8 9 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.85 $Y=2.02 $X2=6.765
+ $Y2=2.02
r35 7 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.77 $Y=2.02
+ $X2=7.855 $Y2=2.02
r36 7 8 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=7.77 $Y=2.02 $X2=6.85
+ $Y2=2.02
r37 2 17 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.71
+ $Y=2.065 $X2=7.855 $Y2=2.21
r38 1 12 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.62
+ $Y=2.065 $X2=6.765 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%Q 1 2 7 8 9 10
r15 9 10 15.7703 $w=2.83e-07 $l=3.9e-07 $layer=LI1_cond $X=12.642 $Y=1.82
+ $X2=12.642 $Y2=2.21
r16 8 9 11.7266 $w=2.83e-07 $l=2.9e-07 $layer=LI1_cond $X=12.642 $Y=1.53
+ $X2=12.642 $Y2=1.82
r17 8 19 36.3929 $w=2.83e-07 $l=9e-07 $layer=LI1_cond $X=12.642 $Y=1.53
+ $X2=12.642 $Y2=0.63
r18 7 19 4.85239 $w=2.83e-07 $l=1.2e-07 $layer=LI1_cond $X=12.642 $Y=0.51
+ $X2=12.642 $Y2=0.63
r19 2 9 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=12.465
+ $Y=1.485 $X2=12.61 $Y2=1.82
r20 1 19 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=12.475
+ $Y=0.235 $X2=12.61 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFRTP_2%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49
+ 51 54 55 57 58 59 61 66 71 76 91 98 105 111 114 117 120 124 127
r195 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r196 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r197 117 118 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r198 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r199 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r200 105 108 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r201 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r202 102 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r203 102 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r204 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r205 99 120 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=12.325 $Y=0
+ $X2=12.115 $Y2=0
r206 99 101 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.325 $Y=0
+ $X2=12.65 $Y2=0
r207 98 123 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=12.995 $Y=0
+ $X2=13.167 $Y2=0
r208 98 101 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.995 $Y=0
+ $X2=12.65 $Y2=0
r209 97 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r210 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r211 94 97 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.73 $Y2=0
r212 93 96 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=10.35 $Y=0
+ $X2=11.73 $Y2=0
r213 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r214 91 120 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=11.905 $Y=0
+ $X2=12.115 $Y2=0
r215 91 96 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=11.905 $Y=0
+ $X2=11.73 $Y2=0
r216 90 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r217 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r218 87 90 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=9.89 $Y2=0
r219 86 89 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=8.05 $Y=0 $X2=9.89
+ $Y2=0
r220 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r221 84 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.05
+ $Y2=0
r222 84 118 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=5.29 $Y2=0
r223 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r224 81 117 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.35 $Y=0
+ $X2=5.177 $Y2=0
r225 81 83 146.139 $w=1.68e-07 $l=2.24e-06 $layer=LI1_cond $X=5.35 $Y=0 $X2=7.59
+ $Y2=0
r226 80 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.29 $Y2=0
r227 80 115 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=2.99 $Y2=0
r228 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r229 77 114 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.035 $Y=0
+ $X2=2.845 $Y2=0
r230 77 79 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=3.035 $Y=0
+ $X2=4.83 $Y2=0
r231 76 117 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=5.005 $Y=0
+ $X2=5.177 $Y2=0
r232 76 79 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.005 $Y=0
+ $X2=4.83 $Y2=0
r233 75 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.99 $Y2=0
r234 75 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.07 $Y2=0
r235 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r236 72 111 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.225 $Y2=0
r237 72 74 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.53 $Y2=0
r238 71 114 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.655 $Y=0
+ $X2=2.845 $Y2=0
r239 71 74 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=0
+ $X2=2.53 $Y2=0
r240 70 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r241 70 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r242 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r243 67 105 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.705 $Y2=0
r244 67 69 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r245 66 111 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.035 $Y=0
+ $X2=2.225 $Y2=0
r246 66 69 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.15
+ $Y2=0
r247 63 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r248 61 105 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.705 $Y2=0
r249 61 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r250 59 106 0.128044 $w=4.8e-07 $l=4.5e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.69 $Y2=0
r251 59 127 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.23 $Y2=0
r252 57 89 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=10.11 $Y=0 $X2=9.89
+ $Y2=0
r253 57 58 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=10.11 $Y=0 $X2=10.22
+ $Y2=0
r254 56 93 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=10.33 $Y=0 $X2=10.35
+ $Y2=0
r255 56 58 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=10.33 $Y=0 $X2=10.22
+ $Y2=0
r256 54 83 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=7.69 $Y=0 $X2=7.59
+ $Y2=0
r257 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.69 $Y=0 $X2=7.855
+ $Y2=0
r258 53 86 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=8.02 $Y=0 $X2=8.05
+ $Y2=0
r259 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.02 $Y=0 $X2=7.855
+ $Y2=0
r260 49 123 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=13.08 $Y=0.085
+ $X2=13.167 $Y2=0
r261 49 51 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.08 $Y=0.085
+ $X2=13.08 $Y2=0.38
r262 45 120 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=12.115 $Y=0.085
+ $X2=12.115 $Y2=0
r263 45 47 10.7013 $w=4.18e-07 $l=3.9e-07 $layer=LI1_cond $X=12.115 $Y=0.085
+ $X2=12.115 $Y2=0.475
r264 41 58 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=10.22 $Y=0.085
+ $X2=10.22 $Y2=0
r265 41 43 14.4055 $w=2.18e-07 $l=2.75e-07 $layer=LI1_cond $X=10.22 $Y=0.085
+ $X2=10.22 $Y2=0.36
r266 37 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=0.085
+ $X2=7.855 $Y2=0
r267 37 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.855 $Y=0.085
+ $X2=7.855 $Y2=0.38
r268 33 117 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.177 $Y=0.085
+ $X2=5.177 $Y2=0
r269 33 35 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=5.177 $Y=0.085
+ $X2=5.177 $Y2=0.455
r270 29 114 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0
r271 29 31 19.8645 $w=3.78e-07 $l=6.55e-07 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0.74
r272 25 111 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0
r273 25 27 11.8277 $w=3.78e-07 $l=3.9e-07 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0.475
r274 8 51 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=12.945
+ $Y=0.235 $X2=13.08 $Y2=0.38
r275 7 47 182 $w=1.7e-07 $l=3.35857e-07 $layer=licon1_NDIFF $count=1 $X=11.865
+ $Y=0.235 $X2=12.095 $Y2=0.475
r276 6 43 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=10.01
+ $Y=0.235 $X2=10.195 $Y2=0.36
r277 5 39 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=7.55
+ $Y=0.235 $X2=7.855 $Y2=0.38
r278 4 35 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.33 $X2=5.185 $Y2=0.455
r279 3 31 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.595 $X2=2.82 $Y2=0.74
r280 2 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.33 $X2=2.25 $Y2=0.475
r281 1 108 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

