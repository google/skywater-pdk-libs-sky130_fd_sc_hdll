# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__and2b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.445000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.630000 1.645000 2.275000 1.955000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.505000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.580000 3.080000 2.365000 ;
        RECT 2.705000 0.255000 3.080000 0.775000 ;
        RECT 2.770000 0.775000 3.080000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.900000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.895000 2.635000 ;
      RECT 0.645000  0.280000 0.885000 0.655000 ;
      RECT 0.665000  0.655000 0.885000 0.805000 ;
      RECT 0.665000  0.805000 1.250000 1.135000 ;
      RECT 0.665000  1.135000 0.900000 1.785000 ;
      RECT 1.070000  1.305000 2.505000 1.325000 ;
      RECT 1.070000  1.325000 2.080000 1.475000 ;
      RECT 1.070000  1.475000 1.405000 2.420000 ;
      RECT 1.215000  0.270000 1.385000 0.415000 ;
      RECT 1.215000  0.415000 1.640000 0.610000 ;
      RECT 1.420000  0.610000 1.640000 0.945000 ;
      RECT 1.420000  0.945000 2.505000 1.305000 ;
      RECT 1.635000  2.165000 2.275000 2.635000 ;
      RECT 2.000000  0.085000 2.445000 0.580000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2b_1
