* File: sky130_fd_sc_hdll__a31oi_2.spice
* Created: Wed Sep  2 08:20:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a31oi_2.pex.spice"
.subckt sky130_fd_sc_hdll__a31oi_2  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1002 N_A_27_47#_M1002_d N_A3_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1012 N_A_27_47#_M1012_d N_A3_M1012_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_A_297_47#_M1005_d N_A2_M1005_g N_A_27_47#_M1012_d VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_A_297_47#_M1005_d N_A2_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g N_A_297_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.11375 PD=1.92 PS=1 NRD=8.304 NRS=4.608 M=1 R=4.33333 SA=75000.2
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_A1_M1004_g N_A_297_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.117 AS=0.11375 PD=1.01 PS=1 NRD=0.912 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.65 AD=0.13
+ AS=0.117 PD=1.05 PS=1.01 NRD=8.304 NRS=13.836 M=1 R=4.33333 SA=75001.2
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1003_d N_B1_M1014_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.65 AD=0.13
+ AS=0.2015 PD=1.05 PS=1.92 NRD=13.836 NRS=8.304 M=1 R=4.33333 SA=75001.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_297#_M1001_d N_A3_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90004.2 A=0.18 P=2.36 MULT=1
MM1006 N_A_27_297#_M1006_d N_A3_M1006_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.8 A=0.18 P=2.36 MULT=1
MM1011 N_A_27_297#_M1006_d N_A2_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90003.3 A=0.18 P=2.36 MULT=1
MM1015 N_A_27_297#_M1015_d N_A2_M1015_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.8 A=0.18 P=2.36 MULT=1
MM1007 N_A_27_297#_M1015_d N_A1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.445 PD=1.29 PS=1.89 NRD=0.9653 NRS=23.6203 M=1 R=5.55556
+ SA=90002.1 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1009_d N_A1_M1009_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.19 AS=0.445 PD=1.38 PS=1.89 NRD=18.715 NRS=29.55 M=1 R=5.55556 SA=90003.1
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1008 N_Y_M1008_d N_B1_M1008_g N_A_27_297#_M1009_d VPB PHIGHVT L=0.18 W=1
+ AD=0.185 AS=0.19 PD=1.37 PS=1.38 NRD=16.7253 NRS=0.9653 M=1 R=5.55556
+ SA=90003.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_Y_M1008_d N_B1_M1010_g N_A_27_297#_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.185 AS=0.27 PD=1.37 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.2 SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
*
.include "sky130_fd_sc_hdll__a31oi_2.pxi.spice"
*
.ends
*
*
