* File: sky130_fd_sc_hdll__clkbuf_6.pxi.spice
* Created: Wed Sep  2 08:25:47 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKBUF_6%A N_A_c_70_n N_A_M1001_g N_A_M1004_g
+ N_A_M1010_g N_A_c_71_n N_A_M1006_g A A N_A_c_69_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_6%A
x_PM_SKY130_FD_SC_HDLL__CLKBUF_6%A_117_297# N_A_117_297#_M1004_s
+ N_A_117_297#_M1001_s N_A_117_297#_c_115_n N_A_117_297#_M1000_g
+ N_A_117_297#_M1005_g N_A_117_297#_M1007_g N_A_117_297#_c_116_n
+ N_A_117_297#_M1002_g N_A_117_297#_c_117_n N_A_117_297#_M1003_g
+ N_A_117_297#_M1011_g N_A_117_297#_M1013_g N_A_117_297#_c_118_n
+ N_A_117_297#_M1008_g N_A_117_297#_c_119_n N_A_117_297#_M1009_g
+ N_A_117_297#_M1014_g N_A_117_297#_M1015_g N_A_117_297#_c_120_n
+ N_A_117_297#_M1012_g N_A_117_297#_c_125_n N_A_117_297#_c_129_n
+ N_A_117_297#_c_113_n N_A_117_297#_c_133_n N_A_117_297#_c_114_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_6%A_117_297#
x_PM_SKY130_FD_SC_HDLL__CLKBUF_6%VPWR N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_M1002_d N_VPWR_M1008_d N_VPWR_M1012_d N_VPWR_c_247_n N_VPWR_c_248_n
+ N_VPWR_c_249_n N_VPWR_c_250_n N_VPWR_c_251_n N_VPWR_c_252_n N_VPWR_c_253_n
+ N_VPWR_c_254_n N_VPWR_c_255_n VPWR N_VPWR_c_256_n N_VPWR_c_257_n
+ N_VPWR_c_246_n N_VPWR_c_259_n N_VPWR_c_260_n N_VPWR_c_261_n N_VPWR_c_262_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_6%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKBUF_6%X N_X_M1005_d N_X_M1011_d N_X_M1014_d
+ N_X_M1000_s N_X_M1003_s N_X_M1009_s N_X_c_317_n N_X_c_323_n N_X_c_327_n
+ N_X_c_309_n N_X_c_310_n N_X_c_339_n N_X_c_343_n N_X_c_347_n N_X_c_311_n
+ N_X_c_355_n N_X_c_312_n N_X_c_362_n N_X_c_313_n N_X_c_369_n N_X_c_314_n
+ N_X_c_376_n X PM_SKY130_FD_SC_HDLL__CLKBUF_6%X
x_PM_SKY130_FD_SC_HDLL__CLKBUF_6%VGND N_VGND_M1004_d N_VGND_M1010_d
+ N_VGND_M1007_s N_VGND_M1013_s N_VGND_M1015_s N_VGND_c_420_n N_VGND_c_421_n
+ N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n N_VGND_c_425_n N_VGND_c_426_n
+ N_VGND_c_427_n N_VGND_c_428_n VGND N_VGND_c_429_n N_VGND_c_430_n
+ N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_6%VGND
cc_1 VNB N_A_M1004_g 0.0317505f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB N_A_M1010_g 0.0284049f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.445
cc_3 VNB A 0.0275664f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_A_c_69_n 0.0612752f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.202
cc_5 VNB N_A_117_297#_M1005_g 0.0287565f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_6 VNB N_A_117_297#_M1007_g 0.0274258f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_7 VNB N_A_117_297#_M1011_g 0.0275253f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=0.85
cc_8 VNB N_A_117_297#_M1013_g 0.0276064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_117_297#_M1014_g 0.027485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_117_297#_M1015_g 0.0345344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_117_297#_c_113_n 0.0037749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_117_297#_c_114_n 0.116556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_246_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_X_c_309_n 0.00641718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_X_c_310_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_X_c_311_n 0.00654821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_X_c_312_n 6.96043e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_X_c_313_n 0.00225504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_314_n 0.0140003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB X 0.015723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_420_n 0.0113827f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_22 VNB N_VGND_c_421_n 0.00461203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_422_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_24 VNB N_VGND_c_423_n 0.0173211f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.202
cc_25 VNB N_VGND_c_424_n 0.00414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_425_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_426_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_427_n 0.0167116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_428_n 0.0170801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_429_n 0.0182311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_430_n 0.0163041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_431_n 0.251742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_432_n 0.00516476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_433_n 0.00515959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_434_n 0.00515959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_435_n 0.00516292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VPB N_A_c_70_n 0.0207627f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_38 VPB N_A_c_71_n 0.0161199f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_39 VPB A 0.00392926f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_40 VPB N_A_c_69_n 0.031942f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.202
cc_41 VPB N_A_117_297#_c_115_n 0.0164402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_117_297#_c_116_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_117_297#_c_117_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_44 VPB N_A_117_297#_c_118_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_117_297#_c_119_n 0.0162548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_117_297#_c_120_n 0.0196139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_117_297#_c_113_n 0.00247361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_117_297#_c_114_n 0.0728182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_247_n 0.0109725f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_50 VPB N_VPWR_c_248_n 0.0429185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_249_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.202
cc_52 VPB N_VPWR_c_250_n 0.0181025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_251_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_252_n 0.0181025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_253_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_254_n 0.0181025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_255_n 0.0288235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_256_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_257_n 0.0163041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_246_n 0.0576986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_259_n 0.0051625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_260_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_261_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_262_n 0.00516583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB X 0.00676826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 N_A_c_71_n N_A_117_297#_c_115_n 0.00970081f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_M1010_g N_A_117_297#_M1005_g 0.0159253f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_M1004_g N_A_117_297#_c_125_n 0.0179655f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_69 N_A_M1010_g N_A_117_297#_c_125_n 0.0155719f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_70 A N_A_117_297#_c_125_n 0.0279461f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_71 N_A_c_69_n N_A_117_297#_c_125_n 0.00709871f $X=0.94 $Y=1.202 $X2=0 $Y2=0
cc_72 N_A_c_70_n N_A_117_297#_c_129_n 0.0154055f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A_c_71_n N_A_117_297#_c_129_n 0.0128277f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_69_n N_A_117_297#_c_129_n 0.00782694f $X=0.94 $Y=1.202 $X2=0 $Y2=0
cc_75 N_A_c_69_n N_A_117_297#_c_113_n 0.0220352f $X=0.94 $Y=1.202 $X2=0 $Y2=0
cc_76 A N_A_117_297#_c_133_n 0.0198664f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_77 N_A_c_69_n N_A_117_297#_c_133_n 0.0181323f $X=0.94 $Y=1.202 $X2=0 $Y2=0
cc_78 N_A_c_69_n N_A_117_297#_c_114_n 0.0210988f $X=0.94 $Y=1.202 $X2=0 $Y2=0
cc_79 N_A_c_70_n N_VPWR_c_248_n 0.00356412f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_80 A N_VPWR_c_248_n 0.0238747f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_81 N_A_c_69_n N_VPWR_c_248_n 0.00214796f $X=0.94 $Y=1.202 $X2=0 $Y2=0
cc_82 N_A_c_71_n N_VPWR_c_249_n 0.00173895f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_c_70_n N_VPWR_c_256_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_71_n N_VPWR_c_256_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_c_70_n N_VPWR_c_246_n 0.0126298f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_c_71_n N_VPWR_c_246_n 0.0117436f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_M1010_g N_X_c_317_n 3.97035e-19 $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_M1010_g N_X_c_310_n 5.27691e-19 $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_89 A N_VGND_c_420_n 0.00101698f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_90 N_A_M1004_g N_VGND_c_421_n 0.00321269f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_91 A N_VGND_c_421_n 0.0213551f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_92 N_A_c_69_n N_VGND_c_421_n 0.00104104f $X=0.94 $Y=1.202 $X2=0 $Y2=0
cc_93 N_A_M1010_g N_VGND_c_422_n 0.00174597f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_M1004_g N_VGND_c_429_n 0.00541763f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_M1010_g N_VGND_c_429_n 0.00541763f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_M1004_g N_VGND_c_431_n 0.0105397f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_M1010_g N_VGND_c_431_n 0.00987959f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_98 A N_VGND_c_431_n 0.00278503f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_99 N_A_117_297#_c_115_n N_VPWR_c_249_n 0.00173895f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_100 N_A_117_297#_c_113_n N_VPWR_c_249_n 0.0186428f $X=3.225 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_117_297#_c_115_n N_VPWR_c_250_n 0.0067375f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_102 N_A_117_297#_c_116_n N_VPWR_c_250_n 0.0067375f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_103 N_A_117_297#_c_116_n N_VPWR_c_251_n 0.00173895f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_104 N_A_117_297#_c_117_n N_VPWR_c_251_n 0.00173895f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_105 N_A_117_297#_c_117_n N_VPWR_c_252_n 0.0067375f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_106 N_A_117_297#_c_118_n N_VPWR_c_252_n 0.0067375f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_107 N_A_117_297#_c_118_n N_VPWR_c_253_n 0.00173895f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_108 N_A_117_297#_c_119_n N_VPWR_c_253_n 0.00173895f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_109 N_A_117_297#_c_119_n N_VPWR_c_254_n 0.0067375f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_110 N_A_117_297#_c_120_n N_VPWR_c_254_n 0.0067375f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_111 N_A_117_297#_c_120_n N_VPWR_c_255_n 0.00354866f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_112 N_A_117_297#_c_129_n N_VPWR_c_256_n 0.0189467f $X=0.73 $Y=1.66 $X2=0
+ $Y2=0
cc_113 N_A_117_297#_M1001_s N_VPWR_c_246_n 0.00231261f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_114 N_A_117_297#_c_115_n N_VPWR_c_246_n 0.0117437f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_115 N_A_117_297#_c_116_n N_VPWR_c_246_n 0.0117185f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_116 N_A_117_297#_c_117_n N_VPWR_c_246_n 0.0117185f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_117 N_A_117_297#_c_118_n N_VPWR_c_246_n 0.0117185f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_118 N_A_117_297#_c_119_n N_VPWR_c_246_n 0.0117185f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_117_297#_c_120_n N_VPWR_c_246_n 0.0130008f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_A_117_297#_c_129_n N_VPWR_c_246_n 0.0123132f $X=0.73 $Y=1.66 $X2=0
+ $Y2=0
cc_121 N_A_117_297#_M1005_g N_X_c_317_n 0.00751737f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_117_297#_M1007_g N_X_c_317_n 0.00791318f $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_123 N_A_117_297#_M1011_g N_X_c_317_n 5.27977e-19 $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_124 N_A_117_297#_c_125_n N_X_c_317_n 0.00324116f $X=0.73 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_117_297#_c_115_n N_X_c_323_n 0.00207151f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_117_297#_c_116_n N_X_c_323_n 5.79575e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_117_297#_c_113_n N_X_c_323_n 0.0214226f $X=3.225 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_117_297#_c_114_n N_X_c_323_n 0.00671335f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_129 N_A_117_297#_c_115_n N_X_c_327_n 0.00850971f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_117_297#_c_116_n N_X_c_327_n 0.00997478f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_117_297#_c_117_n N_X_c_327_n 5.90677e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_117_297#_M1007_g N_X_c_309_n 0.00903265f $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_133 N_A_117_297#_M1011_g N_X_c_309_n 0.00930819f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_134 N_A_117_297#_c_113_n N_X_c_309_n 0.0439086f $X=3.225 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_117_297#_c_114_n N_X_c_309_n 0.00455973f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_136 N_A_117_297#_M1005_g N_X_c_310_n 0.00573192f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A_117_297#_M1007_g N_X_c_310_n 0.00286709f $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_138 N_A_117_297#_c_125_n N_X_c_310_n 0.00469245f $X=0.73 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A_117_297#_c_113_n N_X_c_310_n 0.0269421f $X=3.225 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_117_297#_c_114_n N_X_c_310_n 0.00230339f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_141 N_A_117_297#_c_116_n N_X_c_339_n 0.0137916f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_117_297#_c_117_n N_X_c_339_n 0.0137916f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_117_297#_c_113_n N_X_c_339_n 0.0391038f $X=3.225 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_117_297#_c_114_n N_X_c_339_n 0.00618222f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_145 N_A_117_297#_M1007_g N_X_c_343_n 5.22844e-19 $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_117_297#_M1011_g N_X_c_343_n 0.00772497f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_147 N_A_117_297#_M1013_g N_X_c_343_n 0.00793735f $X=2.82 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A_117_297#_M1014_g N_X_c_343_n 5.26907e-19 $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_117_297#_c_116_n N_X_c_347_n 5.90677e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_117_297#_c_117_n N_X_c_347_n 0.00997478f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_117_297#_c_118_n N_X_c_347_n 0.00997478f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_117_297#_c_119_n N_X_c_347_n 5.90677e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_117_297#_M1013_g N_X_c_311_n 0.00905701f $X=2.82 $Y=0.445 $X2=0 $Y2=0
cc_154 N_A_117_297#_M1014_g N_X_c_311_n 0.00905701f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_155 N_A_117_297#_c_113_n N_X_c_311_n 0.0442765f $X=3.225 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_117_297#_c_114_n N_X_c_311_n 0.00468297f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_157 N_A_117_297#_c_118_n N_X_c_355_n 0.0137916f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_117_297#_c_119_n N_X_c_355_n 0.0137916f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_117_297#_c_113_n N_X_c_355_n 0.039453f $X=3.225 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_117_297#_c_114_n N_X_c_355_n 0.00616252f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_161 N_A_117_297#_M1013_g N_X_c_312_n 5.2762e-19 $X=2.82 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_117_297#_M1014_g N_X_c_312_n 0.00807172f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_117_297#_M1015_g N_X_c_312_n 0.0123142f $X=3.76 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A_117_297#_c_118_n N_X_c_362_n 5.91462e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_117_297#_c_119_n N_X_c_362_n 0.0100507f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_117_297#_c_120_n N_X_c_362_n 0.0144777f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_117_297#_M1011_g N_X_c_313_n 0.00274652f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_168 N_A_117_297#_M1013_g N_X_c_313_n 0.0028989f $X=2.82 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_117_297#_c_113_n N_X_c_313_n 0.0269645f $X=3.225 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_117_297#_c_114_n N_X_c_313_n 0.00243135f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_171 N_A_117_297#_c_117_n N_X_c_369_n 5.79575e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_117_297#_c_118_n N_X_c_369_n 5.79575e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_117_297#_c_113_n N_X_c_369_n 0.0214226f $X=3.225 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_117_297#_c_114_n N_X_c_369_n 0.00669363f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_175 N_A_117_297#_M1014_g N_X_c_314_n 0.0032531f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_176 N_A_117_297#_M1015_g N_X_c_314_n 0.0126708f $X=3.76 $Y=0.445 $X2=0 $Y2=0
cc_177 N_A_117_297#_c_114_n N_X_c_314_n 0.00299987f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_178 N_A_117_297#_c_119_n N_X_c_376_n 7.96011e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_117_297#_c_120_n N_X_c_376_n 0.0148268f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_117_297#_c_114_n N_X_c_376_n 0.00730638f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_181 N_A_117_297#_c_119_n X 4.53853e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_117_297#_M1014_g X 4.94959e-19 $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_183 N_A_117_297#_M1015_g X 0.00403861f $X=3.76 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_117_297#_c_120_n X 0.00421396f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_117_297#_c_113_n X 0.0109381f $X=3.225 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_117_297#_c_114_n X 0.0247582f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_187 N_A_117_297#_M1005_g N_VGND_c_422_n 0.00174597f $X=1.46 $Y=0.445 $X2=0
+ $Y2=0
cc_188 N_A_117_297#_c_113_n N_VGND_c_422_n 0.0108116f $X=3.225 $Y=1.16 $X2=0
+ $Y2=0
cc_189 N_A_117_297#_M1005_g N_VGND_c_423_n 0.00541359f $X=1.46 $Y=0.445 $X2=0
+ $Y2=0
cc_190 N_A_117_297#_M1007_g N_VGND_c_423_n 0.00424416f $X=1.88 $Y=0.445 $X2=0
+ $Y2=0
cc_191 N_A_117_297#_M1007_g N_VGND_c_424_n 0.0016616f $X=1.88 $Y=0.445 $X2=0
+ $Y2=0
cc_192 N_A_117_297#_M1011_g N_VGND_c_424_n 0.0016835f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_193 N_A_117_297#_M1011_g N_VGND_c_425_n 0.00427134f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_A_117_297#_M1013_g N_VGND_c_425_n 0.00424416f $X=2.82 $Y=0.445 $X2=0
+ $Y2=0
cc_195 N_A_117_297#_M1013_g N_VGND_c_426_n 0.00166854f $X=2.82 $Y=0.445 $X2=0
+ $Y2=0
cc_196 N_A_117_297#_M1014_g N_VGND_c_426_n 0.00166854f $X=3.34 $Y=0.445 $X2=0
+ $Y2=0
cc_197 N_A_117_297#_M1014_g N_VGND_c_427_n 0.00423442f $X=3.34 $Y=0.445 $X2=0
+ $Y2=0
cc_198 N_A_117_297#_M1015_g N_VGND_c_427_n 0.00423442f $X=3.76 $Y=0.445 $X2=0
+ $Y2=0
cc_199 N_A_117_297#_M1015_g N_VGND_c_428_n 0.00322276f $X=3.76 $Y=0.445 $X2=0
+ $Y2=0
cc_200 N_A_117_297#_c_125_n N_VGND_c_429_n 0.0177771f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_201 N_A_117_297#_M1004_s N_VGND_c_431_n 0.00217143f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_202 N_A_117_297#_M1005_g N_VGND_c_431_n 0.00987918f $X=1.46 $Y=0.445 $X2=0
+ $Y2=0
cc_203 N_A_117_297#_M1007_g N_VGND_c_431_n 0.00600622f $X=1.88 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_117_297#_M1011_g N_VGND_c_431_n 0.00603609f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_A_117_297#_M1013_g N_VGND_c_431_n 0.00603103f $X=2.82 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A_117_297#_M1014_g N_VGND_c_431_n 0.00603207f $X=3.34 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_117_297#_M1015_g N_VGND_c_431_n 0.00711583f $X=3.76 $Y=0.445 $X2=0
+ $Y2=0
cc_208 N_A_117_297#_c_125_n N_VGND_c_431_n 0.0122848f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_246_n N_X_M1000_s 0.00231418f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_210 N_VPWR_c_246_n N_X_M1003_s 0.00231418f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_211 N_VPWR_c_246_n N_X_M1009_s 0.00231418f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_212 N_VPWR_c_250_n N_X_c_327_n 0.0183657f $X=2.005 $Y=2.72 $X2=0 $Y2=0
cc_213 N_VPWR_c_246_n N_X_c_327_n 0.0122834f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_M1002_d N_X_c_339_n 0.00334388f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_215 N_VPWR_c_251_n N_X_c_339_n 0.0143191f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_216 N_VPWR_c_252_n N_X_c_347_n 0.0183657f $X=2.945 $Y=2.72 $X2=0 $Y2=0
cc_217 N_VPWR_c_246_n N_X_c_347_n 0.0122834f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_M1008_d N_X_c_355_n 0.00334388f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_219 N_VPWR_c_253_n N_X_c_355_n 0.0143191f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_220 N_VPWR_c_254_n N_X_c_362_n 0.0183657f $X=3.885 $Y=2.72 $X2=0 $Y2=0
cc_221 N_VPWR_c_246_n N_X_c_362_n 0.0122834f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_M1012_d N_X_c_376_n 0.00964188f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_223 N_VPWR_c_255_n N_X_c_376_n 0.0115978f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_224 N_VPWR_M1012_d X 8.33267e-19 $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_225 N_X_c_317_n N_VGND_c_423_n 0.0188551f $X=1.67 $Y=0.445 $X2=0 $Y2=0
cc_226 N_X_c_309_n N_VGND_c_423_n 0.00230723f $X=2.445 $Y=0.82 $X2=0 $Y2=0
cc_227 N_X_c_309_n N_VGND_c_424_n 0.0206036f $X=2.445 $Y=0.82 $X2=0 $Y2=0
cc_228 N_X_c_309_n N_VGND_c_425_n 0.00229799f $X=2.445 $Y=0.82 $X2=0 $Y2=0
cc_229 N_X_c_343_n N_VGND_c_425_n 0.0188658f $X=2.61 $Y=0.445 $X2=0 $Y2=0
cc_230 N_X_c_311_n N_VGND_c_425_n 0.00230723f $X=3.385 $Y=0.82 $X2=0 $Y2=0
cc_231 N_X_c_311_n N_VGND_c_426_n 0.0208265f $X=3.385 $Y=0.82 $X2=0 $Y2=0
cc_232 N_X_c_311_n N_VGND_c_427_n 0.00464621f $X=3.385 $Y=0.82 $X2=0 $Y2=0
cc_233 N_X_c_312_n N_VGND_c_427_n 0.0185358f $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_234 N_X_c_314_n N_VGND_c_428_n 0.0147971f $X=3.91 $Y=0.905 $X2=0 $Y2=0
cc_235 N_X_M1005_d N_VGND_c_431_n 0.00216807f $X=1.535 $Y=0.235 $X2=0 $Y2=0
cc_236 N_X_M1011_d N_VGND_c_431_n 0.00220822f $X=2.47 $Y=0.235 $X2=0 $Y2=0
cc_237 N_X_M1014_d N_VGND_c_431_n 0.00216807f $X=3.415 $Y=0.235 $X2=0 $Y2=0
cc_238 N_X_c_317_n N_VGND_c_431_n 0.0123321f $X=1.67 $Y=0.445 $X2=0 $Y2=0
cc_239 N_X_c_309_n N_VGND_c_431_n 0.00860694f $X=2.445 $Y=0.82 $X2=0 $Y2=0
cc_240 N_X_c_343_n N_VGND_c_431_n 0.012355f $X=2.61 $Y=0.445 $X2=0 $Y2=0
cc_241 N_X_c_311_n N_VGND_c_431_n 0.0124963f $X=3.385 $Y=0.82 $X2=0 $Y2=0
cc_242 N_X_c_312_n N_VGND_c_431_n 0.0122362f $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_243 N_X_c_314_n N_VGND_c_431_n 7.07317e-19 $X=3.91 $Y=0.905 $X2=0 $Y2=0
