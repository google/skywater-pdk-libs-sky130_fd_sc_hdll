* File: sky130_fd_sc_hdll__o211ai_4.pex.spice
* Created: Wed Sep  2 08:42:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 30 34 37 45 46
c116 34 0 1.15388e-19 $X=3.855 $Y=1.16
c117 22 0 1.81301e-19 $X=3.895 $Y=0.995
c118 19 0 2.62618e-20 $X=3.86 $Y=1.41
r119 46 47 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.485 $Y2=1.202
r120 44 46 14.8606 $w=3.73e-07 $l=1.15e-07 $layer=POLY_cond $X=1.345 $Y=1.202
+ $X2=1.46 $Y2=1.202
r121 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.345
+ $Y=1.16 $X2=1.345 $Y2=1.16
r122 42 44 47.1662 $w=3.73e-07 $l=3.65e-07 $layer=POLY_cond $X=0.98 $Y=1.202
+ $X2=1.345 $Y2=1.202
r123 39 40 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.475 $Y=1.202
+ $X2=0.5 $Y2=1.202
r124 37 54 1.53625 $w=5.43e-07 $l=7e-08 $layer=LI1_cond $X=1.287 $Y=1.53
+ $X2=1.287 $Y2=1.6
r125 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.855
+ $Y=1.16 $X2=3.855 $Y2=1.16
r126 32 34 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.865 $Y=1.515
+ $X2=3.865 $Y2=1.16
r127 31 54 7.70116 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=1.56 $Y=1.6
+ $X2=1.287 $Y2=1.6
r128 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.7 $Y=1.6
+ $X2=3.865 $Y2=1.515
r129 30 31 139.615 $w=1.68e-07 $l=2.14e-06 $layer=LI1_cond $X=3.7 $Y=1.6
+ $X2=1.56 $Y2=1.6
r130 28 42 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.955 $Y=1.202
+ $X2=0.98 $Y2=1.202
r131 28 40 58.7962 $w=3.73e-07 $l=4.55e-07 $layer=POLY_cond $X=0.955 $Y=1.202
+ $X2=0.5 $Y2=1.202
r132 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=1.16 $X2=0.955 $Y2=1.16
r133 25 37 7.19842 $w=5.43e-07 $l=3.28e-07 $layer=LI1_cond $X=1.287 $Y=1.202
+ $X2=1.287 $Y2=1.53
r134 25 45 0.921749 $w=5.43e-07 $l=4.2e-08 $layer=LI1_cond $X=1.287 $Y=1.202
+ $X2=1.287 $Y2=1.16
r135 25 27 2.71163 $w=2.53e-07 $l=6e-08 $layer=LI1_cond $X=1.015 $Y=1.202
+ $X2=0.955 $Y2=1.202
r136 22 35 38.7084 $w=3.43e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.895 $Y=0.995
+ $X2=3.88 $Y2=1.16
r137 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.895 $Y=0.995
+ $X2=3.895 $Y2=0.56
r138 19 35 45.964 $w=3.43e-07 $l=2.59808e-07 $layer=POLY_cond $X=3.86 $Y=1.41
+ $X2=3.88 $Y2=1.16
r139 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.86 $Y=1.41
+ $X2=3.86 $Y2=1.985
r140 16 47 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.485 $Y2=1.202
r141 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.485 $Y2=0.56
r142 13 46 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.46 $Y=1.41
+ $X2=1.46 $Y2=1.202
r143 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.46 $Y=1.41
+ $X2=1.46 $Y2=1.985
r144 10 42 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.202
r145 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.985
r146 7 28 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=1.202
r147 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r148 4 40 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.202
r149 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
r150 1 39 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.202
r151 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 43
r76 39 40 3.03526 $w=3.97e-07 $l=2.5e-08 $layer=POLY_cond $X=3.38 $Y=1.202
+ $X2=3.405 $Y2=1.202
r77 37 39 23.068 $w=3.97e-07 $l=1.9e-07 $layer=POLY_cond $X=3.19 $Y=1.202
+ $X2=3.38 $Y2=1.202
r78 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.19
+ $Y=1.16 $X2=3.19 $Y2=1.16
r79 35 37 35.2091 $w=3.97e-07 $l=2.9e-07 $layer=POLY_cond $X=2.9 $Y=1.202
+ $X2=3.19 $Y2=1.202
r80 34 35 3.03526 $w=3.97e-07 $l=2.5e-08 $layer=POLY_cond $X=2.875 $Y=1.202
+ $X2=2.9 $Y2=1.202
r81 33 34 55.2418 $w=3.97e-07 $l=4.55e-07 $layer=POLY_cond $X=2.42 $Y=1.202
+ $X2=2.875 $Y2=1.202
r82 32 33 3.03526 $w=3.97e-07 $l=2.5e-08 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.42 $Y2=1.202
r83 30 32 45.529 $w=3.97e-07 $l=3.75e-07 $layer=POLY_cond $X=2.02 $Y=1.202
+ $X2=2.395 $Y2=1.202
r84 30 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.02
+ $Y=1.16 $X2=2.02 $Y2=1.16
r85 28 30 9.71285 $w=3.97e-07 $l=8e-08 $layer=POLY_cond $X=1.94 $Y=1.202
+ $X2=2.02 $Y2=1.202
r86 27 28 3.03526 $w=3.97e-07 $l=2.5e-08 $layer=POLY_cond $X=1.915 $Y=1.202
+ $X2=1.94 $Y2=1.202
r87 25 38 28.1708 $w=2.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.53 $Y=1.21
+ $X2=3.19 $Y2=1.21
r88 25 43 21.7684 $w=2.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.53 $Y=1.21
+ $X2=2.02 $Y2=1.21
r89 22 40 25.678 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.405 $Y=0.995
+ $X2=3.405 $Y2=1.202
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.405 $Y=0.995
+ $X2=3.405 $Y2=0.56
r91 19 39 21.283 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.202
r92 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.985
r93 16 35 21.283 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.9 $Y=1.41 $X2=2.9
+ $Y2=1.202
r94 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.9 $Y=1.41 $X2=2.9
+ $Y2=1.985
r95 13 34 25.678 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.875 $Y=0.995
+ $X2=2.875 $Y2=1.202
r96 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.875 $Y=0.995
+ $X2=2.875 $Y2=0.56
r97 10 33 21.283 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.42 $Y=1.41
+ $X2=2.42 $Y2=1.202
r98 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.42 $Y=1.41
+ $X2=2.42 $Y2=1.985
r99 7 32 25.678 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.395 $Y=0.995
+ $X2=2.395 $Y2=1.202
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.395 $Y=0.995
+ $X2=2.395 $Y2=0.56
r101 4 28 21.283 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.94 $Y=1.41
+ $X2=1.94 $Y2=1.202
r102 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.94 $Y=1.41
+ $X2=1.94 $Y2=1.985
r103 1 27 25.678 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.915 $Y=0.995
+ $X2=1.915 $Y2=1.202
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.915 $Y=0.995
+ $X2=1.915 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 30 34 37 47 51 52 56
c113 47 0 1.97811e-19 $X=5.34 $Y=1.202
c114 16 0 1.91217e-19 $X=5.365 $Y=0.995
r115 51 52 4.05212 $w=6.88e-07 $l=1.25e-07 $layer=LI1_cond $X=4.835 $Y=1.34
+ $X2=4.71 $Y2=1.34
r116 47 48 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=5.34 $Y=1.202
+ $X2=5.365 $Y2=1.202
r117 46 51 6.76044 $w=6.88e-07 $l=3.9e-07 $layer=LI1_cond $X=5.225 $Y=1.34
+ $X2=4.835 $Y2=1.34
r118 45 47 14.8606 $w=3.73e-07 $l=1.15e-07 $layer=POLY_cond $X=5.225 $Y=1.202
+ $X2=5.34 $Y2=1.202
r119 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.225
+ $Y=1.16 $X2=5.225 $Y2=1.16
r120 43 45 47.1662 $w=3.73e-07 $l=3.65e-07 $layer=POLY_cond $X=4.86 $Y=1.202
+ $X2=5.225 $Y2=1.202
r121 42 43 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=4.835 $Y=1.202
+ $X2=4.86 $Y2=1.202
r122 39 40 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=4.355 $Y=1.202
+ $X2=4.38 $Y2=1.202
r123 37 56 11.8676 $w=6.88e-07 $l=2.3e-07 $layer=LI1_cond $X=5.295 $Y=1.34
+ $X2=5.525 $Y2=1.34
r124 37 46 1.21341 $w=6.88e-07 $l=7e-08 $layer=LI1_cond $X=5.295 $Y=1.34
+ $X2=5.225 $Y2=1.34
r125 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.665
+ $Y=1.16 $X2=7.665 $Y2=1.16
r126 32 34 18.5962 $w=2.18e-07 $l=3.55e-07 $layer=LI1_cond $X=7.69 $Y=1.515
+ $X2=7.69 $Y2=1.16
r127 30 32 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.58 $Y=1.6
+ $X2=7.69 $Y2=1.515
r128 30 56 134.07 $w=1.68e-07 $l=2.055e-06 $layer=LI1_cond $X=7.58 $Y=1.6
+ $X2=5.525 $Y2=1.6
r129 28 42 50.3968 $w=3.73e-07 $l=3.9e-07 $layer=POLY_cond $X=4.445 $Y=1.202
+ $X2=4.835 $Y2=1.202
r130 28 40 8.39946 $w=3.73e-07 $l=6.5e-08 $layer=POLY_cond $X=4.445 $Y=1.202
+ $X2=4.38 $Y2=1.202
r131 27 52 7.35897 $w=4.13e-07 $l=2.65e-07 $layer=LI1_cond $X=4.445 $Y=1.202
+ $X2=4.71 $Y2=1.202
r132 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.445
+ $Y=1.16 $X2=4.445 $Y2=1.16
r133 22 35 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=7.775 $Y=0.995
+ $X2=7.69 $Y2=1.16
r134 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.775 $Y=0.995
+ $X2=7.775 $Y2=0.56
r135 19 35 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=7.69 $Y=1.41
+ $X2=7.69 $Y2=1.16
r136 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.69 $Y=1.41
+ $X2=7.69 $Y2=1.985
r137 16 48 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.365 $Y=0.995
+ $X2=5.365 $Y2=1.202
r138 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.365 $Y=0.995
+ $X2=5.365 $Y2=0.56
r139 13 47 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.34 $Y=1.41
+ $X2=5.34 $Y2=1.202
r140 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.34 $Y=1.41
+ $X2=5.34 $Y2=1.985
r141 10 43 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.86 $Y=1.41
+ $X2=4.86 $Y2=1.202
r142 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.86 $Y=1.41
+ $X2=4.86 $Y2=1.985
r143 7 42 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.835 $Y=0.995
+ $X2=4.835 $Y2=1.202
r144 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.835 $Y=0.995
+ $X2=4.835 $Y2=0.56
r145 4 40 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.38 $Y=1.41
+ $X2=4.38 $Y2=1.202
r146 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.38 $Y=1.41
+ $X2=4.38 $Y2=1.985
r147 1 39 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.355 $Y=0.995
+ $X2=4.355 $Y2=1.202
r148 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.355 $Y=0.995
+ $X2=4.355 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%C1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 41 42 46
c80 41 0 1.97811e-19 $X=6.975 $Y=1.16
c81 22 0 1.88158e-19 $X=7.245 $Y=0.995
r82 42 43 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.22 $Y=1.202
+ $X2=7.245 $Y2=1.202
r83 40 42 31.7446 $w=3.72e-07 $l=2.45e-07 $layer=POLY_cond $X=6.975 $Y=1.202
+ $X2=7.22 $Y2=1.202
r84 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.975
+ $Y=1.16 $X2=6.975 $Y2=1.16
r85 38 40 29.1532 $w=3.72e-07 $l=2.25e-07 $layer=POLY_cond $X=6.75 $Y=1.202
+ $X2=6.975 $Y2=1.202
r86 37 38 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.725 $Y=1.202
+ $X2=6.75 $Y2=1.202
r87 35 37 18.1398 $w=3.72e-07 $l=1.4e-07 $layer=POLY_cond $X=6.585 $Y=1.202
+ $X2=6.725 $Y2=1.202
r88 33 35 39.5188 $w=3.72e-07 $l=3.05e-07 $layer=POLY_cond $X=6.28 $Y=1.202
+ $X2=6.585 $Y2=1.202
r89 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.255 $Y=1.202
+ $X2=6.28 $Y2=1.202
r90 30 32 7.77419 $w=3.72e-07 $l=6e-08 $layer=POLY_cond $X=6.195 $Y=1.202
+ $X2=6.255 $Y2=1.202
r91 30 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.195
+ $Y=1.16 $X2=6.195 $Y2=1.16
r92 28 30 49.8844 $w=3.72e-07 $l=3.85e-07 $layer=POLY_cond $X=5.81 $Y=1.202
+ $X2=6.195 $Y2=1.202
r93 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.785 $Y=1.202
+ $X2=5.81 $Y2=1.202
r94 25 41 16.6464 $w=2.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.585 $Y=1.21
+ $X2=6.975 $Y2=1.21
r95 25 46 16.6464 $w=2.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.585 $Y=1.21
+ $X2=6.195 $Y2=1.21
r96 25 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.585
+ $Y=1.16 $X2=6.585 $Y2=1.16
r97 22 43 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.245 $Y=0.995
+ $X2=7.245 $Y2=1.202
r98 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.245 $Y=0.995
+ $X2=7.245 $Y2=0.56
r99 19 42 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.22 $Y=1.41
+ $X2=7.22 $Y2=1.202
r100 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.22 $Y=1.41
+ $X2=7.22 $Y2=1.985
r101 16 38 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.75 $Y=1.41
+ $X2=6.75 $Y2=1.202
r102 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.75 $Y=1.41
+ $X2=6.75 $Y2=1.985
r103 13 37 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.725 $Y=0.995
+ $X2=6.725 $Y2=1.202
r104 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.725 $Y=0.995
+ $X2=6.725 $Y2=0.56
r105 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.28 $Y=1.41
+ $X2=6.28 $Y2=1.202
r106 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.28 $Y=1.41
+ $X2=6.28 $Y2=1.985
r107 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.255 $Y=0.995
+ $X2=6.255 $Y2=1.202
r108 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.255 $Y=0.995
+ $X2=6.255 $Y2=0.56
r109 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.81 $Y=1.41
+ $X2=5.81 $Y2=1.202
r110 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.81 $Y=1.41
+ $X2=5.81 $Y2=1.985
r111 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.785 $Y=0.995
+ $X2=5.785 $Y2=1.202
r112 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.785 $Y=0.995
+ $X2=5.785 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%VPWR 1 2 3 4 5 6 7 22 24 28 30 32 35 36
+ 38 41 45 48 51 53 71 75 84 91 99
r120 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r121 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r122 84 87 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.195 $Y=2.36
+ $X2=1.195 $Y2=2.72
r123 79 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r124 79 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.13 $Y2=2.72
r125 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r126 76 78 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=7.155 $Y=2.72
+ $X2=8.05 $Y2=2.72
r127 75 98 4.49945 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=8.155 $Y=2.72
+ $X2=8.447 $Y2=2.72
r128 75 78 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.155 $Y=2.72
+ $X2=8.05 $Y2=2.72
r129 74 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r130 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r131 71 76 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=6.962 $Y=2.72
+ $X2=7.155 $Y2=2.72
r132 71 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r133 71 91 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=6.962 $Y=2.72
+ $X2=6.962 $Y2=2.36
r134 71 73 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.77 $Y=2.72 $X2=6.67
+ $Y2=2.72
r135 70 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r136 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r137 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r138 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r139 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r140 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r141 61 64 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r142 61 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 60 63 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r144 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r145 58 87 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.385 $Y=2.72
+ $X2=1.195 $Y2=2.72
r146 58 60 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.385 $Y=2.72
+ $X2=1.61 $Y2=2.72
r147 57 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r149 54 81 4.46799 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r150 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r151 53 87 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=1.195 $Y2=2.72
r152 53 56 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=0.69 $Y2=2.72
r153 51 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r154 51 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r155 49 73 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r156 48 69 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=5.83 $Y=2.72 $X2=5.75
+ $Y2=2.72
r157 47 49 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.02 $Y=2.72
+ $X2=6.21 $Y2=2.72
r158 47 48 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.02 $Y=2.72
+ $X2=5.83 $Y2=2.72
r159 45 47 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=6.02 $Y=2.36
+ $X2=6.02 $Y2=2.72
r160 42 69 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.265 $Y=2.72
+ $X2=5.75 $Y2=2.72
r161 41 66 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.885 $Y=2.72
+ $X2=4.83 $Y2=2.72
r162 40 42 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.075 $Y=2.72
+ $X2=5.265 $Y2=2.72
r163 40 41 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.075 $Y=2.72
+ $X2=4.885 $Y2=2.72
r164 38 40 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.075 $Y=2.36
+ $X2=5.075 $Y2=2.72
r165 35 63 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=3.91 $Y2=2.72
r166 35 36 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=4.15 $Y2=2.72
r167 34 66 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.285 $Y=2.72
+ $X2=4.83 $Y2=2.72
r168 34 36 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.285 $Y=2.72
+ $X2=4.15 $Y2=2.72
r169 30 98 3.26672 $w=3.3e-07 $l=1.64085e-07 $layer=LI1_cond $X=8.32 $Y=2.635
+ $X2=8.447 $Y2=2.72
r170 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.32 $Y=2.635
+ $X2=8.32 $Y2=2.36
r171 26 36 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.15 $Y=2.635
+ $X2=4.15 $Y2=2.72
r172 26 28 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.15 $Y=2.635
+ $X2=4.15 $Y2=2.36
r173 22 81 3.00953 $w=2.95e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.192 $Y2=2.72
r174 22 24 31.448 $w=2.93e-07 $l=8.05e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.237 $Y2=1.83
r175 7 32 600 $w=1.7e-07 $l=1.11271e-06 $layer=licon1_PDIFF $count=1 $X=7.78
+ $Y=1.485 $X2=8.32 $Y2=2.36
r176 6 91 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.485 $X2=6.985 $Y2=2.36
r177 5 45 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=5.9
+ $Y=1.485 $X2=6.045 $Y2=2.36
r178 4 38 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.485 $X2=5.1 $Y2=2.36
r179 3 28 600 $w=1.7e-07 $l=9.5623e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.485 $X2=4.12 $Y2=2.36
r180 2 84 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.485 $X2=1.22 $Y2=2.36
r181 1 24 300 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%A_118_297# 1 2 3 4 13 19 23 27
r42 21 23 56.0383 $w=1.88e-07 $l=9.6e-07 $layer=LI1_cond $X=2.66 $Y=2.37
+ $X2=3.62 $Y2=2.37
r43 19 21 51.0766 $w=1.88e-07 $l=8.75e-07 $layer=LI1_cond $X=1.785 $Y=2.37
+ $X2=2.66 $Y2=2.37
r44 16 19 6.82297 $w=1.9e-07 $l=1.32571e-07 $layer=LI1_cond $X=1.695 $Y=2.275
+ $X2=1.785 $Y2=2.37
r45 16 18 7.08586 $w=1.78e-07 $l=1.15e-07 $layer=LI1_cond $X=1.695 $Y=2.275
+ $X2=1.695 $Y2=2.16
r46 15 18 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=1.695 $Y=2.105
+ $X2=1.695 $Y2=2.16
r47 14 27 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.825 $Y=2.02
+ $X2=0.715 $Y2=2.02
r48 13 15 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.605 $Y=2.02
+ $X2=1.695 $Y2=2.105
r49 13 14 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.605 $Y=2.02
+ $X2=0.825 $Y2=2.02
r50 4 23 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.485 $X2=3.62 $Y2=2.36
r51 3 21 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.51
+ $Y=1.485 $X2=2.66 $Y2=2.36
r52 2 18 600 $w=1.7e-07 $l=7.46241e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.485 $X2=1.7 $Y2=2.16
r53 1 27 600 $w=1.7e-07 $l=6.1041e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=2.025
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%Y 1 2 3 4 5 6 7 8 25 33 40 41 42 45 46 47
+ 48 51 55 64
c115 33 0 1.91217e-19 $X=7.265 $Y=0.36
c116 25 0 2.62618e-20 $X=3.695 $Y=1.98
r117 59 61 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=6.515 $Y=1.98
+ $X2=7.455 $Y2=1.98
r118 57 59 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.575 $Y=1.98
+ $X2=6.515 $Y2=1.98
r119 54 57 44.0233 $w=2.48e-07 $l=9.55e-07 $layer=LI1_cond $X=4.62 $Y=1.98
+ $X2=5.575 $Y2=1.98
r120 54 55 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4.62 $Y=1.98
+ $X2=4.495 $Y2=1.98
r121 51 64 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=8.23 $Y=1.98
+ $X2=8.125 $Y2=1.98
r122 48 64 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=8.08 $Y=1.98
+ $X2=8.125 $Y2=1.98
r123 48 61 28.8111 $w=2.48e-07 $l=6.25e-07 $layer=LI1_cond $X=8.08 $Y=1.98
+ $X2=7.455 $Y2=1.98
r124 48 51 0.837255 $w=4.98e-07 $l=3.5e-08 $layer=LI1_cond $X=8.23 $Y=1.82
+ $X2=8.23 $Y2=1.855
r125 46 48 5.50196 $w=4.98e-07 $l=2.3e-07 $layer=LI1_cond $X=8.23 $Y=1.59
+ $X2=8.23 $Y2=1.82
r126 46 47 11.1517 $w=4.98e-07 $l=2.5e-07 $layer=LI1_cond $X=8.23 $Y=1.59
+ $X2=8.23 $Y2=1.34
r127 45 55 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.82 $Y=1.94
+ $X2=4.495 $Y2=1.94
r128 43 47 31.7323 $w=1.78e-07 $l=5.15e-07 $layer=LI1_cond $X=8.07 $Y=0.825
+ $X2=8.07 $Y2=1.34
r129 41 43 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.98 $Y=0.74
+ $X2=8.07 $Y2=0.825
r130 41 42 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.98 $Y=0.74
+ $X2=7.485 $Y2=0.74
r131 40 42 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.375 $Y=0.655
+ $X2=7.485 $Y2=0.74
r132 39 40 10.7387 $w=2.18e-07 $l=2.05e-07 $layer=LI1_cond $X=7.375 $Y=0.45
+ $X2=7.375 $Y2=0.655
r133 35 38 57.9192 $w=1.78e-07 $l=9.4e-07 $layer=LI1_cond $X=6.045 $Y=0.36
+ $X2=6.985 $Y2=0.36
r134 33 39 6.90553 $w=1.8e-07 $l=1.48324e-07 $layer=LI1_cond $X=7.265 $Y=0.36
+ $X2=7.375 $Y2=0.45
r135 33 38 17.2525 $w=1.78e-07 $l=2.8e-07 $layer=LI1_cond $X=7.265 $Y=0.36
+ $X2=6.985 $Y2=0.36
r136 27 30 44.2538 $w=2.48e-07 $l=9.6e-07 $layer=LI1_cond $X=2.18 $Y=1.98
+ $X2=3.14 $Y2=1.98
r137 25 45 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.695 $Y=1.98
+ $X2=3.82 $Y2=1.98
r138 25 30 25.5842 $w=2.48e-07 $l=5.55e-07 $layer=LI1_cond $X=3.695 $Y=1.98
+ $X2=3.14 $Y2=1.98
r139 8 61 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=7.31
+ $Y=1.485 $X2=7.455 $Y2=1.94
r140 7 59 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=6.37
+ $Y=1.485 $X2=6.515 $Y2=1.94
r141 6 57 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=1.485 $X2=5.575 $Y2=1.94
r142 5 54 600 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.485 $X2=4.62 $Y2=1.94
r143 4 30 600 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.485 $X2=3.14 $Y2=1.94
r144 3 27 600 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.485 $X2=2.18 $Y2=1.94
r145 2 38 182 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_NDIFF $count=1 $X=6.8
+ $Y=0.235 $X2=6.985 $Y2=0.365
r146 1 35 182 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_NDIFF $count=1 $X=5.86
+ $Y=0.235 $X2=6.045 $Y2=0.365
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%A_27_47# 1 2 3 4 5 6 7 22 24 25 30 32 34
+ 41 42 43 49 59
c128 42 0 1.15388e-19 $X=8.26 $Y=0.51
c129 34 0 1.88158e-19 $X=8.32 $Y=0.395
c130 30 0 1.4234e-19 $X=4.235 $Y=0.355
r131 56 58 39.302 $w=2.98e-07 $l=9.6e-07 $layer=LI1_cond $X=2.18 $Y=0.665
+ $X2=3.14 $Y2=0.665
r132 50 59 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.405 $Y=0.51
+ $X2=8.405 $Y2=0.395
r133 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.405 $Y=0.51
+ $X2=8.405 $Y2=0.51
r134 46 56 37.8691 $w=2.98e-07 $l=9.25e-07 $layer=LI1_cond $X=1.255 $Y=0.665
+ $X2=2.18 $Y2=0.665
r135 46 53 1.43289 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.255 $Y=0.665
+ $X2=1.22 $Y2=0.665
r136 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.255 $Y=0.51
+ $X2=1.255 $Y2=0.51
r137 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.4 $Y=0.51
+ $X2=1.255 $Y2=0.51
r138 42 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.26 $Y=0.51
+ $X2=8.405 $Y2=0.51
r139 42 43 8.49008 $w=1.4e-07 $l=6.86e-06 $layer=MET1_cond $X=8.26 $Y=0.51
+ $X2=1.4 $Y2=0.51
r140 39 41 3.66807 $w=3.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.26 $Y=0.72
+ $X2=0.355 $Y2=0.72
r141 34 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.32 $Y=0.395
+ $X2=8.405 $Y2=0.395
r142 34 36 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.32 $Y=0.395
+ $X2=7.99 $Y2=0.395
r143 30 32 47.9682 $w=1.98e-07 $l=8.65e-07 $layer=LI1_cond $X=4.235 $Y=0.355
+ $X2=5.1 $Y2=0.355
r144 27 29 6.51381 $w=2.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.12 $Y=0.625
+ $X2=4.12 $Y2=0.495
r145 26 30 6.85974 $w=2e-07 $l=1.57242e-07 $layer=LI1_cond $X=4.12 $Y=0.455
+ $X2=4.235 $Y2=0.355
r146 26 29 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=4.12 $Y=0.455
+ $X2=4.12 $Y2=0.495
r147 25 58 16.1516 $w=2.98e-07 $l=3.61801e-07 $layer=LI1_cond $X=3.48 $Y=0.71
+ $X2=3.14 $Y2=0.665
r148 24 27 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.005 $Y=0.71
+ $X2=4.12 $Y2=0.625
r149 24 25 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.005 $Y=0.71
+ $X2=3.48 $Y2=0.71
r150 22 53 3.94911 $w=2.98e-07 $l=1.39642e-07 $layer=LI1_cond $X=1.125 $Y=0.765
+ $X2=1.22 $Y2=0.665
r151 22 41 31.6922 $w=2.78e-07 $l=7.7e-07 $layer=LI1_cond $X=1.125 $Y=0.765
+ $X2=0.355 $Y2=0.765
r152 7 36 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.85
+ $Y=0.235 $X2=7.99 $Y2=0.395
r153 6 32 182 $w=1.7e-07 $l=2.46577e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.235 $X2=5.1 $Y2=0.365
r154 5 29 182 $w=1.7e-07 $l=3.26497e-07 $layer=licon1_NDIFF $count=1 $X=3.97
+ $Y=0.235 $X2=4.12 $Y2=0.495
r155 4 58 182 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_NDIFF $count=1 $X=2.95
+ $Y=0.235 $X2=3.14 $Y2=0.71
r156 3 56 182 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.235 $X2=2.18 $Y2=0.71
r157 2 53 182 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.22 $Y2=0.71
r158 1 39 182 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%VGND 1 2 3 4 13 17 19 21 23 28 38 39 43
+ 49 53 60
c119 60 0 1.4234e-19 $X=3.45 $Y=0
r120 60 63 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=3.595 $Y2=0.36
r121 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r122 54 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r123 53 56 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.635 $Y=0
+ $X2=2.635 $Y2=0.36
r124 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r125 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r126 44 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r127 43 46 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.715 $Y=0
+ $X2=0.715 $Y2=0.36
r128 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r129 38 39 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r130 36 39 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=3.91 $Y=0 $X2=8.51
+ $Y2=0
r131 36 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r132 35 38 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=8.51
+ $Y2=0
r133 35 36 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r134 33 60 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.595
+ $Y2=0
r135 33 35 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.785 $Y=0
+ $X2=3.91 $Y2=0
r136 32 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r137 32 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r138 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r139 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.7
+ $Y2=0
r140 29 31 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=2.07 $Y2=0
r141 28 53 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.635
+ $Y2=0
r142 28 31 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.07 $Y2=0
r143 23 43 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.715
+ $Y2=0
r144 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.23
+ $Y2=0
r145 21 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r146 21 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r147 20 53 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.635
+ $Y2=0
r148 19 60 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.595
+ $Y2=0
r149 19 20 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.405 $Y=0
+ $X2=2.825 $Y2=0
r150 15 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r151 15 17 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.7 $Y=0.085
+ $X2=1.7 $Y2=0.36
r152 14 43 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.715
+ $Y2=0
r153 13 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.7
+ $Y2=0
r154 13 14 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=0.905 $Y2=0
r155 4 63 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.48
+ $Y=0.235 $X2=3.62 $Y2=0.36
r156 3 56 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.235 $X2=2.66 $Y2=0.36
r157 2 17 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.7 $Y2=0.36
r158 1 46 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.74 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_4%A_886_47# 1 2 11
c27 11 0 1.81301e-19 $X=6.515 $Y=0.725
r28 8 11 116.763 $w=1.78e-07 $l=1.895e-06 $layer=LI1_cond $X=4.62 $Y=0.725
+ $X2=6.515 $Y2=0.725
r29 2 11 182 $w=1.7e-07 $l=5.75109e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.235 $X2=6.515 $Y2=0.725
r30 1 8 182 $w=1.7e-07 $l=5.82301e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.235 $X2=4.62 $Y2=0.73
.ends

