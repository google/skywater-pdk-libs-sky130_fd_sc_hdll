* File: sky130_fd_sc_hdll__a31oi_2.pex.spice
* Created: Wed Sep  2 08:20:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%A3 1 3 4 6 7 9 10 12 13 15 26 34
r40 26 27 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r41 25 34 1.73624 $w=6.18e-07 $l=9e-08 $layer=LI1_cond $X=0.605 $Y=1.305
+ $X2=0.695 $Y2=1.305
r42 24 26 47.5397 $w=3.65e-07 $l=3.6e-07 $layer=POLY_cond $X=0.605 $Y=1.202
+ $X2=0.965 $Y2=1.202
r43 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.16 $X2=0.605 $Y2=1.16
r44 22 24 11.2247 $w=3.65e-07 $l=8.5e-08 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.605 $Y2=1.202
r45 21 22 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r46 15 34 0.964579 $w=6.18e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.305
+ $X2=0.695 $Y2=1.305
r47 13 25 7.13789 $w=6.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.305
+ $X2=0.605 $Y2=1.305
r48 10 27 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r49 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r50 7 26 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r51 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r52 4 22 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r53 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r54 1 21 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r55 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%A2 1 3 4 6 7 9 10 12 13 15 26 32 35 37
r46 35 37 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=1.77 $Y=1.305
+ $X2=1.775 $Y2=1.305
r47 26 27 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r48 24 26 10.7816 $w=3.8e-07 $l=8.5e-08 $layer=POLY_cond $X=1.82 $Y=1.202
+ $X2=1.905 $Y2=1.202
r49 24 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.82
+ $Y=1.16 $X2=1.82 $Y2=1.16
r50 22 24 48.8342 $w=3.8e-07 $l=3.85e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.82 $Y2=1.202
r51 21 22 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r52 15 35 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=1.765 $Y=1.305
+ $X2=1.77 $Y2=1.305
r53 15 32 9.54934 $w=6.18e-07 $l=4.95e-07 $layer=LI1_cond $X=1.765 $Y=1.305
+ $X2=1.27 $Y2=1.305
r54 13 32 0.289374 $w=6.18e-07 $l=1.5e-08 $layer=LI1_cond $X=1.255 $Y=1.305
+ $X2=1.27 $Y2=1.305
r55 10 27 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r56 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r57 7 26 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r58 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r59 4 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r60 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r61 1 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%A1 1 3 4 5 6 8 9 11 12 14 15 17 27 30 34
+ 37 39
c58 27 0 1.44908e-19 $X=3.445 $Y=1.202
r59 37 39 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=2.985 $Y=1.305
+ $X2=2.99 $Y2=1.305
r60 27 28 3.38483 $w=3.56e-07 $l=2.5e-08 $layer=POLY_cond $X=3.445 $Y=1.202
+ $X2=3.47 $Y2=1.202
r61 25 27 59.573 $w=3.56e-07 $l=4.4e-07 $layer=POLY_cond $X=3.005 $Y=1.202
+ $X2=3.445 $Y2=1.202
r62 25 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.005
+ $Y=1.16 $X2=3.005 $Y2=1.16
r63 23 25 4.73876 $w=3.56e-07 $l=3.5e-08 $layer=POLY_cond $X=2.97 $Y=1.202
+ $X2=3.005 $Y2=1.202
r64 17 37 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=2.98 $Y=1.305
+ $X2=2.985 $Y2=1.305
r65 17 34 10.0316 $w=6.18e-07 $l=5.2e-07 $layer=LI1_cond $X=2.98 $Y=1.305
+ $X2=2.46 $Y2=1.305
r66 15 34 0.192916 $w=6.18e-07 $l=1e-08 $layer=LI1_cond $X=2.45 $Y=1.305
+ $X2=2.46 $Y2=1.305
r67 15 30 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=2.45 $Y=1.305
+ $X2=2.445 $Y2=1.305
r68 12 28 23.0368 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.47 $Y=0.995
+ $X2=3.47 $Y2=1.202
r69 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.47 $Y=0.995
+ $X2=3.47 $Y2=0.56
r70 9 27 18.7059 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.445 $Y=1.41
+ $X2=3.445 $Y2=1.202
r71 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.445 $Y=1.41
+ $X2=3.445 $Y2=1.985
r72 6 23 23.0368 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.97 $Y=0.995
+ $X2=2.97 $Y2=1.202
r73 6 8 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.97 $Y=0.995 $X2=2.97
+ $Y2=0.56
r74 4 23 10.4875 $w=3.56e-07 $l=9.3675e-08 $layer=POLY_cond $X=2.895 $Y=1.16
+ $X2=2.97 $Y2=1.202
r75 4 5 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.895 $Y=1.16
+ $X2=2.475 $Y2=1.16
r76 1 5 30.0773 $w=3.3e-07 $l=2.95804e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.475 $Y2=1.16
r77 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%B1 1 3 4 6 7 9 11 12 14 15 16 17 18 24 28
+ 32
c54 28 0 1.44908e-19 $X=4.715 $Y=1.175
r55 28 32 19.4091 $w=1.98e-07 $l=3.5e-07 $layer=LI1_cond $X=4.715 $Y=1.175
+ $X2=4.365 $Y2=1.175
r56 24 26 29.0521 $w=3.65e-07 $l=2.2e-07 $layer=POLY_cond $X=4.555 $Y=1.202
+ $X2=4.775 $Y2=1.202
r57 23 24 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=4.53 $Y=1.202
+ $X2=4.555 $Y2=1.202
r58 17 28 3.6174 $w=2e-07 $l=1.12e-07 $layer=LI1_cond $X=4.827 $Y=1.175
+ $X2=4.715 $Y2=1.175
r59 17 18 9.55671 $w=3.93e-07 $l=2.55e-07 $layer=LI1_cond $X=4.827 $Y=1.275
+ $X2=4.827 $Y2=1.53
r60 17 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.775
+ $Y=1.16 $X2=4.775 $Y2=1.16
r61 16 32 3.32727 $w=1.98e-07 $l=6e-08 $layer=LI1_cond $X=4.305 $Y=1.175
+ $X2=4.365 $Y2=1.175
r62 12 24 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.555 $Y=1.41
+ $X2=4.555 $Y2=1.202
r63 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.555 $Y=1.41
+ $X2=4.555 $Y2=1.985
r64 9 23 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.53 $Y=0.995
+ $X2=4.53 $Y2=1.202
r65 9 11 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.53 $Y=0.995
+ $X2=4.53 $Y2=0.56
r66 8 15 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=4.105 $Y=1.16
+ $X2=4.005 $Y2=1.202
r67 7 23 10.4484 $w=3.65e-07 $l=9.3675e-08 $layer=POLY_cond $X=4.455 $Y=1.16
+ $X2=4.53 $Y2=1.202
r68 7 8 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=4.455 $Y=1.16
+ $X2=4.105 $Y2=1.16
r69 4 15 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=4.005 $Y=1.41
+ $X2=4.005 $Y2=1.202
r70 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.005 $Y=1.41
+ $X2=4.005 $Y2=1.985
r71 1 15 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=3.98 $Y=0.995
+ $X2=4.005 $Y2=1.202
r72 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.98 $Y=0.995 $X2=3.98
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%A_27_297# 1 2 3 4 5 18 22 26 28 29 30 31
+ 34 37 39 41
r67 32 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.79 $Y=2.295
+ $X2=4.79 $Y2=1.96
r68 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.705 $Y=2.38
+ $X2=4.79 $Y2=2.295
r69 30 31 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=4.705 $Y=2.38
+ $X2=3.855 $Y2=2.38
r70 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.77 $Y=2.295
+ $X2=3.855 $Y2=2.38
r71 28 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=1.955
+ $X2=3.77 $Y2=1.87
r72 28 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.77 $Y=1.955
+ $X2=3.77 $Y2=2.295
r73 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=1.87
+ $X2=2.14 $Y2=1.87
r74 26 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=1.87
+ $X2=3.77 $Y2=1.87
r75 26 27 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=3.685 $Y=1.87
+ $X2=2.225 $Y2=1.87
r76 23 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=1.87 $X2=1.2
+ $Y2=1.87
r77 22 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.87
+ $X2=2.14 $Y2=1.87
r78 22 23 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=1.87
+ $X2=1.285 $Y2=1.87
r79 19 37 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.87
+ $X2=0.26 $Y2=1.87
r80 18 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=1.87 $X2=1.2
+ $Y2=1.87
r81 18 19 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=1.87
+ $X2=0.345 $Y2=1.87
r82 5 34 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.645
+ $Y=1.485 $X2=4.79 $Y2=1.96
r83 4 43 300 $w=1.7e-07 $l=5.70526e-07 $layer=licon1_PDIFF $count=2 $X=3.535
+ $Y=1.485 $X2=3.77 $Y2=1.95
r84 3 41 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.95
r85 2 39 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.95
r86 1 37 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%VPWR 1 2 3 12 16 18 20 25 40 41 44 47 52
+ 55
r71 54 55 11.5558 $w=6.78e-07 $l=2.15e-07 $layer=LI1_cond $X=3.065 $Y=2.465
+ $X2=3.28 $Y2=2.465
r72 50 54 1.3192 $w=6.78e-07 $l=7.5e-08 $layer=LI1_cond $X=2.99 $Y=2.465
+ $X2=3.065 $Y2=2.465
r73 50 52 15.3376 $w=6.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.99 $Y=2.465
+ $X2=2.56 $Y2=2.465
r74 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r75 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r76 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r78 38 41 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r79 38 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r80 37 40 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r81 37 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.28 $Y2=2.72
r82 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 34 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r84 34 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r85 33 52 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.53 $Y=2.72 $X2=2.56
+ $Y2=2.72
r86 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r87 31 47 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=1.645 $Y2=2.72
r88 31 33 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=2.53 $Y2=2.72
r89 29 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r90 29 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r91 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r92 26 44 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r93 26 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 25 47 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.645 $Y2=2.72
r95 25 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r96 20 44 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r97 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r98 18 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r99 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r100 14 47 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2.72
r101 14 16 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2.21
r102 10 44 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r103 10 12 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.21
r104 3 54 300 $w=1.7e-07 $l=9.80115e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=3.065 $Y2=2.21
r105 2 16 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.21
r106 1 12 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%Y 1 2 3 4 13 19 21 23 27 30 34 35 36 45
r75 42 45 0.182927 $w=3.13e-07 $l=5e-09 $layer=LI1_cond $X=3.487 $Y=0.845
+ $X2=3.487 $Y2=0.85
r76 35 36 7.75597 $w=4.83e-07 $l=2.55e-07 $layer=LI1_cond $X=3.487 $Y=1.19
+ $X2=3.487 $Y2=1.445
r77 34 42 2.19354 $w=3.15e-07 $l=1.23288e-07 $layer=LI1_cond $X=3.552 $Y=0.75
+ $X2=3.487 $Y2=0.845
r78 34 35 10.9756 $w=3.13e-07 $l=3e-07 $layer=LI1_cond $X=3.487 $Y=0.89
+ $X2=3.487 $Y2=1.19
r79 34 45 1.46342 $w=3.13e-07 $l=4e-08 $layer=LI1_cond $X=3.487 $Y=0.89
+ $X2=3.487 $Y2=0.85
r80 30 32 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.765 $Y=0.38
+ $X2=4.765 $Y2=0.75
r81 25 27 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.32 $Y=1.615
+ $X2=4.32 $Y2=1.63
r82 24 34 4.00438 $w=1.9e-07 $l=2.23e-07 $layer=LI1_cond $X=3.775 $Y=0.75
+ $X2=3.552 $Y2=0.75
r83 23 32 4.80115 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.575 $Y=0.75
+ $X2=4.765 $Y2=0.75
r84 23 24 46.6986 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=4.575 $Y=0.75
+ $X2=3.775 $Y2=0.75
r85 22 36 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=3.645 $Y=1.53
+ $X2=3.487 $Y2=1.53
r86 21 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.155 $Y=1.53
+ $X2=4.32 $Y2=1.615
r87 21 22 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.155 $Y=1.53
+ $X2=3.645 $Y2=1.53
r88 17 34 2.19354 $w=1.7e-07 $l=1.79315e-07 $layer=LI1_cond $X=3.69 $Y=0.655
+ $X2=3.552 $Y2=0.75
r89 17 19 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.69 $Y=0.655
+ $X2=3.69 $Y2=0.42
r90 13 34 4.00438 $w=1.7e-07 $l=2.26945e-07 $layer=LI1_cond $X=3.33 $Y=0.74
+ $X2=3.552 $Y2=0.75
r91 13 15 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.33 $Y=0.74
+ $X2=2.71 $Y2=0.74
r92 4 27 300 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=2 $X=4.095
+ $Y=1.485 $X2=4.32 $Y2=1.63
r93 3 30 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=4.605
+ $Y=0.235 $X2=4.79 $Y2=0.38
r94 2 34 182 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_NDIFF $count=1 $X=3.545
+ $Y=0.235 $X2=3.69 $Y2=0.76
r95 2 19 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.545
+ $Y=0.235 $X2=3.69 $Y2=0.42
r96 1 15 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.235 $X2=2.71 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%A_27_47# 1 2 3 16
r22 14 16 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.2 $Y=0.74 $X2=2.14
+ $Y2=0.74
r23 11 14 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.26 $Y=0.74 $X2=1.2
+ $Y2=0.74
r24 3 16 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.74
r25 2 14 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.74
r26 1 11 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%VGND 1 2 7 8 14 16 29 30 34
r54 34 37 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.705
+ $Y2=0.38
r55 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r56 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r57 27 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r58 26 27 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r59 24 27 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.91
+ $Y2=0
r60 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r61 23 26 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.91
+ $Y2=0
r62 23 24 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r63 21 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r64 21 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r65 16 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r66 16 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r67 14 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r68 14 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r69 10 29 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.83
+ $Y2=0
r70 8 26 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.025 $Y=0 $X2=3.91
+ $Y2=0
r71 7 12 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=4.215
+ $Y2=0.38
r72 7 10 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=4.405
+ $Y2=0
r73 7 8 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=4.025
+ $Y2=0
r74 2 12 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=4.055
+ $Y=0.235 $X2=4.24 $Y2=0.38
r75 1 37 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31OI_2%A_297_47# 1 2 11
r20 8 11 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=1.67 $Y=0.38
+ $X2=3.21 $Y2=0.38
r21 2 11 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=3.045
+ $Y=0.235 $X2=3.21 $Y2=0.38
r22 1 8 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.38
.ends

