# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.300000 1.075000 8.760000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.380000 0.995000 7.600000 1.445000 ;
        RECT 7.380000 1.445000 8.010000 1.665000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.255000 0.995000 2.940000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.517500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.330000 0.660000 0.930000 0.925000 ;
        RECT 0.330000 0.925000 0.695000 1.440000 ;
        RECT 0.330000 1.440000 0.905000 2.045000 ;
        RECT 0.655000 2.045000 0.905000 2.465000 ;
        RECT 0.680000 0.350000 0.930000 0.660000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.105000  0.085000 0.435000 0.465000 ;
      RECT 0.105000  2.215000 0.435000 2.635000 ;
      RECT 1.095000  0.995000 1.295000 1.325000 ;
      RECT 1.105000  0.085000 1.355000 0.525000 ;
      RECT 1.125000  0.695000 1.745000 0.865000 ;
      RECT 1.125000  0.865000 1.295000 0.995000 ;
      RECT 1.125000  1.325000 1.295000 1.875000 ;
      RECT 1.125000  1.875000 1.865000 2.045000 ;
      RECT 1.125000  2.215000 1.460000 2.635000 ;
      RECT 1.525000  0.255000 3.190000 0.425000 ;
      RECT 1.525000  0.425000 1.745000 0.695000 ;
      RECT 1.530000  1.535000 3.280000 1.705000 ;
      RECT 1.645000  2.045000 1.865000 2.235000 ;
      RECT 1.645000  2.235000 3.340000 2.405000 ;
      RECT 1.915000  0.595000 2.085000 1.535000 ;
      RECT 2.265000  1.895000 3.670000 2.065000 ;
      RECT 2.365000  0.655000 3.575000 0.825000 ;
      RECT 2.785000  0.425000 3.190000 0.455000 ;
      RECT 3.110000  0.995000 3.435000 1.325000 ;
      RECT 3.110000  1.325000 3.280000 1.535000 ;
      RECT 3.360000  0.255000 4.255000 0.425000 ;
      RECT 3.360000  0.425000 3.575000 0.655000 ;
      RECT 3.500000  1.525000 4.030000 1.695000 ;
      RECT 3.500000  1.695000 3.670000 1.895000 ;
      RECT 3.605000  2.235000 4.010000 2.405000 ;
      RECT 3.745000  0.595000 3.915000 1.375000 ;
      RECT 3.745000  1.375000 4.030000 1.525000 ;
      RECT 3.840000  1.895000 5.115000 2.065000 ;
      RECT 3.840000  2.065000 4.010000 2.235000 ;
      RECT 4.085000  0.425000 4.255000 1.035000 ;
      RECT 4.085000  1.035000 4.370000 1.205000 ;
      RECT 4.180000  2.235000 4.510000 2.635000 ;
      RECT 4.200000  1.205000 4.370000 1.895000 ;
      RECT 4.425000  0.085000 4.595000 0.865000 ;
      RECT 4.600000  1.445000 5.115000 1.715000 ;
      RECT 4.825000  0.415000 5.115000 1.445000 ;
      RECT 4.945000  2.065000 5.115000 2.275000 ;
      RECT 4.945000  2.275000 8.240000 2.445000 ;
      RECT 5.290000  0.265000 5.705000 0.485000 ;
      RECT 5.290000  0.485000 5.510000 0.595000 ;
      RECT 5.290000  0.595000 5.460000 2.105000 ;
      RECT 5.630000  0.720000 6.095000 0.825000 ;
      RECT 5.630000  0.825000 5.900000 0.890000 ;
      RECT 5.630000  0.890000 5.800000 2.275000 ;
      RECT 5.680000  0.655000 6.095000 0.720000 ;
      RECT 5.925000  0.320000 6.095000 0.655000 ;
      RECT 6.040000  1.445000 6.870000 1.615000 ;
      RECT 6.040000  1.615000 6.455000 2.045000 ;
      RECT 6.055000  0.995000 6.480000 1.270000 ;
      RECT 6.265000  0.630000 6.480000 0.995000 ;
      RECT 6.700000  0.255000 7.895000 0.425000 ;
      RECT 6.700000  0.425000 6.870000 1.445000 ;
      RECT 7.040000  0.595000 7.210000 1.935000 ;
      RECT 7.040000  1.935000 9.550000 2.105000 ;
      RECT 7.380000  0.425000 7.895000 0.465000 ;
      RECT 7.770000  0.730000 7.975000 0.945000 ;
      RECT 7.770000  0.945000 8.090000 1.275000 ;
      RECT 8.230000  1.495000 9.100000 1.705000 ;
      RECT 8.270000  0.295000 8.560000 0.735000 ;
      RECT 8.270000  0.735000 9.100000 0.750000 ;
      RECT 8.310000  0.750000 9.100000 0.905000 ;
      RECT 8.650000  2.275000 9.035000 2.635000 ;
      RECT 8.780000  0.085000 8.950000 0.565000 ;
      RECT 8.930000  0.905000 9.100000 0.995000 ;
      RECT 8.930000  0.995000 9.210000 1.325000 ;
      RECT 8.930000  1.325000 9.100000 1.495000 ;
      RECT 9.015000  1.875000 9.550000 1.935000 ;
      RECT 9.250000  0.255000 9.550000 0.585000 ;
      RECT 9.255000  2.105000 9.550000 2.465000 ;
      RECT 9.380000  0.585000 9.550000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.860000  1.445000 4.030000 1.615000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 4.830000  0.765000 5.000000 0.935000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.340000  0.425000 5.510000 0.595000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.310000  0.765000 6.480000 0.935000 ;
      RECT 6.310000  1.445000 6.480000 1.615000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.790000  0.765000 7.960000 0.935000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.300000  0.425000 8.470000 0.595000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 3.800000 1.415000 4.090000 1.460000 ;
      RECT 3.800000 1.460000 6.540000 1.600000 ;
      RECT 3.800000 1.600000 4.090000 1.645000 ;
      RECT 4.770000 0.735000 5.060000 0.780000 ;
      RECT 4.770000 0.780000 8.020000 0.920000 ;
      RECT 4.770000 0.920000 5.060000 0.965000 ;
      RECT 5.280000 0.395000 5.570000 0.440000 ;
      RECT 5.280000 0.440000 8.530000 0.580000 ;
      RECT 5.280000 0.580000 5.570000 0.625000 ;
      RECT 6.250000 0.735000 6.540000 0.780000 ;
      RECT 6.250000 0.920000 6.540000 0.965000 ;
      RECT 6.250000 1.415000 6.540000 1.460000 ;
      RECT 6.250000 1.600000 6.540000 1.645000 ;
      RECT 7.730000 0.735000 8.020000 0.780000 ;
      RECT 7.730000 0.920000 8.020000 0.965000 ;
      RECT 8.240000 0.395000 8.530000 0.440000 ;
      RECT 8.240000 0.580000 8.530000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor3_2
