# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o211a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o211a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.825000 1.035000 5.155000 1.495000 ;
        RECT 4.825000 1.495000 6.815000 1.685000 ;
        RECT 6.300000 1.035000 6.815000 1.495000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.340000 1.035000 6.115000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 0.995000 3.085000 1.445000 ;
        RECT 2.790000 1.445000 4.600000 1.685000 ;
        RECT 4.270000 1.035000 4.600000 1.445000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255000 1.035000 4.090000 1.275000 ;
    END
  END C1
  PIN VGND
    ANTENNADIFFAREA  1.069250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.795000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  1.016000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 1.755000 0.805000 ;
        RECT 0.085000 0.805000 0.365000 1.435000 ;
        RECT 0.085000 1.435000 2.230000 1.700000 ;
        RECT 0.645000 0.255000 0.815000 0.615000 ;
        RECT 0.645000 0.615000 1.755000 0.635000 ;
        RECT 1.080000 1.700000 1.260000 2.465000 ;
        RECT 1.585000 0.255000 1.755000 0.615000 ;
        RECT 2.040000 1.700000 2.230000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.480000  1.870000 0.860000 2.635000 ;
      RECT 0.535000  1.065000 2.620000 1.265000 ;
      RECT 1.035000  0.085000 1.365000 0.445000 ;
      RECT 1.440000  1.870000 1.820000 2.635000 ;
      RECT 1.925000  0.085000 2.340000 0.465000 ;
      RECT 2.400000  0.635000 3.820000 0.815000 ;
      RECT 2.400000  0.815000 2.620000 1.065000 ;
      RECT 2.400000  1.265000 2.620000 1.855000 ;
      RECT 2.400000  1.855000 5.845000 2.025000 ;
      RECT 2.400000  2.200000 2.780000 2.635000 ;
      RECT 2.580000  0.255000 4.805000 0.465000 ;
      RECT 3.000000  2.025000 3.360000 2.465000 ;
      RECT 3.535000  2.195000 3.915000 2.635000 ;
      RECT 4.085000  2.025000 4.415000 2.465000 ;
      RECT 4.475000  0.465000 4.805000 0.695000 ;
      RECT 4.475000  0.695000 6.805000 0.865000 ;
      RECT 4.595000  2.195000 4.860000 2.635000 ;
      RECT 4.980000  0.085000 5.295000 0.525000 ;
      RECT 5.465000  0.255000 5.845000 0.695000 ;
      RECT 5.465000  2.025000 5.845000 2.465000 ;
      RECT 6.065000  0.085000 6.255000 0.525000 ;
      RECT 6.425000  0.255000 6.805000 0.695000 ;
      RECT 6.425000  1.915000 6.805000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211a_4
