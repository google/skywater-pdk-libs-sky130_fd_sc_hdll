* File: sky130_fd_sc_hdll__or4b_4.pxi.spice
* Created: Wed Sep  2 08:49:49 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR4B_4%D_N N_D_N_c_94_n N_D_N_c_95_n N_D_N_M1003_g
+ N_D_N_M1013_g D_N D_N D_N N_D_N_c_91_n N_D_N_c_92_n N_D_N_c_93_n
+ PM_SKY130_FD_SC_HDLL__OR4B_4%D_N
x_PM_SKY130_FD_SC_HDLL__OR4B_4%A_117_413# N_A_117_413#_M1013_d
+ N_A_117_413#_M1003_d N_A_117_413#_c_121_n N_A_117_413#_M1017_g
+ N_A_117_413#_c_116_n N_A_117_413#_M1014_g N_A_117_413#_c_117_n
+ N_A_117_413#_c_118_n N_A_117_413#_c_119_n N_A_117_413#_c_124_n
+ N_A_117_413#_c_120_n PM_SKY130_FD_SC_HDLL__OR4B_4%A_117_413#
x_PM_SKY130_FD_SC_HDLL__OR4B_4%C N_C_c_165_n N_C_M1008_g N_C_c_166_n N_C_M1012_g
+ C C N_C_c_167_n PM_SKY130_FD_SC_HDLL__OR4B_4%C
x_PM_SKY130_FD_SC_HDLL__OR4B_4%B N_B_c_198_n N_B_M1006_g N_B_c_199_n N_B_M1007_g
+ B B N_B_c_200_n PM_SKY130_FD_SC_HDLL__OR4B_4%B
x_PM_SKY130_FD_SC_HDLL__OR4B_4%A N_A_c_229_n N_A_M1005_g N_A_c_230_n N_A_M1001_g
+ A N_A_c_231_n A PM_SKY130_FD_SC_HDLL__OR4B_4%A
x_PM_SKY130_FD_SC_HDLL__OR4B_4%A_225_297# N_A_225_297#_M1014_d
+ N_A_225_297#_M1007_d N_A_225_297#_M1017_s N_A_225_297#_c_267_n
+ N_A_225_297#_M1002_g N_A_225_297#_c_275_n N_A_225_297#_M1000_g
+ N_A_225_297#_c_268_n N_A_225_297#_M1010_g N_A_225_297#_c_276_n
+ N_A_225_297#_M1004_g N_A_225_297#_c_269_n N_A_225_297#_M1015_g
+ N_A_225_297#_c_277_n N_A_225_297#_M1009_g N_A_225_297#_c_278_n
+ N_A_225_297#_M1011_g N_A_225_297#_c_270_n N_A_225_297#_M1016_g
+ N_A_225_297#_c_279_n N_A_225_297#_c_271_n N_A_225_297#_c_291_n
+ N_A_225_297#_c_300_n N_A_225_297#_c_292_n N_A_225_297#_c_391_p
+ N_A_225_297#_c_312_n N_A_225_297#_c_272_n N_A_225_297#_c_273_n
+ N_A_225_297#_c_341_p N_A_225_297#_c_307_n N_A_225_297#_c_274_n
+ PM_SKY130_FD_SC_HDLL__OR4B_4%A_225_297#
x_PM_SKY130_FD_SC_HDLL__OR4B_4%VPWR N_VPWR_M1003_s N_VPWR_M1001_d N_VPWR_M1004_d
+ N_VPWR_M1011_d N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n N_VPWR_c_412_n
+ N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n
+ N_VPWR_c_418_n VPWR N_VPWR_c_419_n N_VPWR_c_408_n
+ PM_SKY130_FD_SC_HDLL__OR4B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__OR4B_4%X N_X_M1002_d N_X_M1015_d N_X_M1000_s N_X_M1009_s
+ N_X_c_486_n N_X_c_530_n N_X_c_495_n N_X_c_487_n N_X_c_480_n N_X_c_481_n
+ N_X_c_513_n N_X_c_534_n N_X_c_488_n N_X_c_482_n N_X_c_483_n N_X_c_489_n X
+ N_X_c_485_n PM_SKY130_FD_SC_HDLL__OR4B_4%X
x_PM_SKY130_FD_SC_HDLL__OR4B_4%VGND N_VGND_M1013_s N_VGND_M1014_s N_VGND_M1012_d
+ N_VGND_M1005_d N_VGND_M1010_s N_VGND_M1016_s N_VGND_c_559_n N_VGND_c_560_n
+ N_VGND_c_561_n N_VGND_c_562_n N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n
+ N_VGND_c_566_n N_VGND_c_567_n N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n
+ N_VGND_c_571_n N_VGND_c_572_n N_VGND_c_573_n VGND N_VGND_c_574_n
+ N_VGND_c_575_n N_VGND_c_576_n PM_SKY130_FD_SC_HDLL__OR4B_4%VGND
cc_1 VNB N_D_N_c_91_n 0.0364574f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_2 VNB N_D_N_c_92_n 0.0178988f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_3 VNB N_D_N_c_93_n 0.0216313f $X=-0.19 $Y=-0.24 $X2=0.42 $Y2=0.995
cc_4 VNB N_A_117_413#_c_116_n 0.0210474f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_5 VNB N_A_117_413#_c_117_n 0.0285858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_117_413#_c_118_n 0.013179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_117_413#_c_119_n 0.00623381f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_8 VNB N_A_117_413#_c_120_n 0.0128281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C_c_165_n 0.0240388f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_10 VNB N_C_c_166_n 0.0176935f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_11 VNB N_C_c_167_n 0.00325865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_198_n 0.0236499f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_13 VNB N_B_c_199_n 0.01695f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_14 VNB N_B_c_200_n 0.00358189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_c_229_n 0.0177853f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_16 VNB N_A_c_230_n 0.0240735f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_17 VNB N_A_c_231_n 0.00326942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_225_297#_c_267_n 0.0171624f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_19 VNB N_A_225_297#_c_268_n 0.0167557f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_20 VNB N_A_225_297#_c_269_n 0.0171987f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.19
cc_21 VNB N_A_225_297#_c_270_n 0.0200831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_225_297#_c_271_n 0.00303358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_225_297#_c_272_n 0.0016277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_225_297#_c_273_n 0.00376665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_225_297#_c_274_n 0.0762306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_408_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_480_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_481_n 0.0017592f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.53
cc_29 VNB N_X_c_482_n 0.00123315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_483_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB X 0.0203361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_485_n 0.00836446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_559_n 0.0099134f $X=-0.19 $Y=-0.24 $X2=0.42 $Y2=1.325
cc_34 VNB N_VGND_c_560_n 0.035093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_561_n 0.0222418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_562_n 0.0122395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_563_n 0.00226425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_564_n 0.00260546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_565_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_566_n 0.0116103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_567_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_568_n 0.0195679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_569_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_570_n 0.0173964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_571_n 0.00609289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_572_n 0.0178379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_573_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_574_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_575_n 0.00478242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_576_n 0.296804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VPB N_D_N_c_94_n 0.0403638f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_52 VPB N_D_N_c_95_n 0.0325653f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_53 VPB N_D_N_c_91_n 0.00774063f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_54 VPB N_D_N_c_92_n 0.029026f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_55 VPB N_A_117_413#_c_121_n 0.0202626f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.675
cc_56 VPB N_A_117_413#_c_117_n 0.0106932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_117_413#_c_118_n 0.00700981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_117_413#_c_124_n 0.0177562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_117_413#_c_120_n 0.00867269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_C_c_165_n 0.0272173f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_61 VPB N_C_c_167_n 0.00221474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_B_c_198_n 0.0248843f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_63 VPB N_B_c_200_n 0.00213307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_c_230_n 0.0258087f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_65 VPB A 0.00423925f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.675
cc_66 VPB N_A_c_231_n 0.0026021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_225_297#_c_275_n 0.0171649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_225_297#_c_276_n 0.0159743f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.325
cc_69 VPB N_A_225_297#_c_277_n 0.0159556f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.87
cc_70 VPB N_A_225_297#_c_278_n 0.0191486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_225_297#_c_279_n 0.00719937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_225_297#_c_271_n 0.00315676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_225_297#_c_274_n 0.0467455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_409_n 0.0102718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_410_n 0.0197397f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.16
cc_76 VPB N_VPWR_c_411_n 0.00519418f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.325
cc_77 VPB N_VPWR_c_412_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_413_n 0.012247f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.87
cc_79 VPB N_VPWR_c_414_n 0.00518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_415_n 0.0795937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_416_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_417_n 0.0213107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_418_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_419_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_408_n 0.0560021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_X_c_486_n 0.00190706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_X_c_487_n 0.00206401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_X_c_488_n 0.0110582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_X_c_489_n 0.00161374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB X 0.00758585f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 N_D_N_c_91_n N_A_117_413#_c_117_n 0.0076468f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_92 N_D_N_c_93_n N_A_117_413#_c_119_n 0.00656725f $X=0.42 $Y=0.995 $X2=0 $Y2=0
cc_93 N_D_N_c_94_n N_A_117_413#_c_124_n 0.0164501f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_94 N_D_N_c_95_n N_A_117_413#_c_124_n 0.00608791f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_95 N_D_N_c_92_n N_A_117_413#_c_124_n 0.0422858f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_96 N_D_N_c_91_n N_A_117_413#_c_120_n 0.00410583f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_97 N_D_N_c_92_n N_A_117_413#_c_120_n 0.02434f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_98 N_D_N_c_95_n N_VPWR_c_410_n 0.00465874f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_99 N_D_N_c_92_n N_VPWR_c_410_n 0.0212332f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_100 N_D_N_c_95_n N_VPWR_c_415_n 0.00743866f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_101 N_D_N_c_95_n N_VPWR_c_408_n 0.0141405f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_102 N_D_N_c_92_n N_VPWR_c_408_n 0.00400376f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_103 N_D_N_c_91_n N_VGND_c_560_n 9.41854e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_104 N_D_N_c_92_n N_VGND_c_560_n 0.021392f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_105 N_D_N_c_93_n N_VGND_c_560_n 0.00624463f $X=0.42 $Y=0.995 $X2=0 $Y2=0
cc_106 N_D_N_c_93_n N_VGND_c_561_n 0.00510437f $X=0.42 $Y=0.995 $X2=0 $Y2=0
cc_107 N_D_N_c_93_n N_VGND_c_562_n 0.00284681f $X=0.42 $Y=0.995 $X2=0 $Y2=0
cc_108 N_D_N_c_93_n N_VGND_c_576_n 0.00512902f $X=0.42 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_117_413#_c_121_n N_C_c_165_n 0.0336954f $X=1.485 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_110 N_A_117_413#_c_118_n N_C_c_165_n 0.0180946f $X=1.485 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_117_413#_c_116_n N_C_c_166_n 0.0203587f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_117_413#_c_121_n N_C_c_167_n 0.00613269f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_117_413#_c_118_n N_C_c_167_n 5.28091e-19 $X=1.485 $Y=1.202 $X2=0
+ $Y2=0
cc_114 N_A_117_413#_c_121_n N_A_225_297#_c_279_n 0.0127789f $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_115 N_A_117_413#_c_124_n N_A_225_297#_c_279_n 0.0425016f $X=0.73 $Y=2.275
+ $X2=0 $Y2=0
cc_116 N_A_117_413#_c_121_n N_A_225_297#_c_271_n 0.0228366f $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_117 N_A_117_413#_c_116_n N_A_225_297#_c_271_n 0.0064014f $X=1.51 $Y=0.995
+ $X2=0 $Y2=0
cc_118 N_A_117_413#_c_117_n N_A_225_297#_c_271_n 0.00719285f $X=1.385 $Y=1.16
+ $X2=0 $Y2=0
cc_119 N_A_117_413#_c_118_n N_A_225_297#_c_271_n 0.0134001f $X=1.485 $Y=1.202
+ $X2=0 $Y2=0
cc_120 N_A_117_413#_c_119_n N_A_225_297#_c_271_n 0.00429539f $X=0.73 $Y=0.74
+ $X2=0 $Y2=0
cc_121 N_A_117_413#_c_124_n N_A_225_297#_c_271_n 0.0173144f $X=0.73 $Y=2.275
+ $X2=0 $Y2=0
cc_122 N_A_117_413#_c_120_n N_A_225_297#_c_271_n 0.0290772f $X=1.18 $Y=1.16
+ $X2=0 $Y2=0
cc_123 N_A_117_413#_c_116_n N_A_225_297#_c_291_n 0.00446123f $X=1.51 $Y=0.995
+ $X2=0 $Y2=0
cc_124 N_A_117_413#_c_116_n N_A_225_297#_c_292_n 0.00923831f $X=1.51 $Y=0.995
+ $X2=0 $Y2=0
cc_125 N_A_117_413#_c_119_n N_A_225_297#_c_292_n 0.00445089f $X=0.73 $Y=0.74
+ $X2=0 $Y2=0
cc_126 N_A_117_413#_c_121_n N_VPWR_c_415_n 0.00674013f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_127 N_A_117_413#_c_124_n N_VPWR_c_415_n 0.0124228f $X=0.73 $Y=2.275 $X2=0
+ $Y2=0
cc_128 N_A_117_413#_M1003_d N_VPWR_c_408_n 0.00480007f $X=0.585 $Y=2.065 $X2=0
+ $Y2=0
cc_129 N_A_117_413#_c_121_n N_VPWR_c_408_n 0.0135759f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_130 N_A_117_413#_c_124_n N_VPWR_c_408_n 0.00720598f $X=0.73 $Y=2.275 $X2=0
+ $Y2=0
cc_131 N_A_117_413#_c_119_n N_VGND_c_560_n 0.0107285f $X=0.73 $Y=0.74 $X2=0
+ $Y2=0
cc_132 N_A_117_413#_c_119_n N_VGND_c_561_n 0.00616648f $X=0.73 $Y=0.74 $X2=0
+ $Y2=0
cc_133 N_A_117_413#_c_116_n N_VGND_c_562_n 0.00725468f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_A_117_413#_c_117_n N_VGND_c_562_n 0.00593141f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_117_413#_c_119_n N_VGND_c_562_n 0.00879006f $X=0.73 $Y=0.74 $X2=0
+ $Y2=0
cc_136 N_A_117_413#_c_120_n N_VGND_c_562_n 0.00758226f $X=1.18 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_117_413#_c_116_n N_VGND_c_563_n 0.0013206f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_138 N_A_117_413#_c_116_n N_VGND_c_568_n 0.00501458f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_139 N_A_117_413#_c_116_n N_VGND_c_576_n 0.00982726f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_140 N_A_117_413#_c_119_n N_VGND_c_576_n 0.00646895f $X=0.73 $Y=0.74 $X2=0
+ $Y2=0
cc_141 N_C_c_165_n N_B_c_198_n 0.0781262f $X=2.065 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_142 N_C_c_167_n N_B_c_198_n 0.00296382f $X=1.98 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_143 N_C_c_166_n N_B_c_199_n 0.0215326f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_144 N_C_c_165_n N_B_c_200_n 0.00396354f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_145 N_C_c_167_n N_B_c_200_n 0.0688036f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_146 N_C_c_165_n N_A_225_297#_c_279_n 9.12912e-19 $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_147 N_C_c_167_n N_A_225_297#_c_279_n 0.0216532f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_148 N_C_c_165_n N_A_225_297#_c_271_n 0.00354158f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_149 N_C_c_166_n N_A_225_297#_c_271_n 0.00340748f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_150 N_C_c_167_n N_A_225_297#_c_271_n 0.0588966f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_151 N_C_c_166_n N_A_225_297#_c_291_n 0.00540738f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_152 N_C_c_165_n N_A_225_297#_c_300_n 7.10472e-19 $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_153 N_C_c_166_n N_A_225_297#_c_300_n 0.0120102f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_154 N_C_c_167_n N_A_225_297#_c_300_n 0.0195869f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_155 N_C_c_165_n N_A_225_297#_c_292_n 0.00189854f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_156 N_C_c_165_n N_VPWR_c_415_n 0.00450951f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_157 N_C_c_167_n N_VPWR_c_415_n 0.0106463f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_158 N_C_c_165_n N_VPWR_c_408_n 0.00647188f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_159 N_C_c_167_n N_VPWR_c_408_n 0.00970516f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_160 N_C_c_167_n A_315_297# 0.0114441f $X=1.98 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_161 N_C_c_166_n N_VGND_c_563_n 0.0117441f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_162 N_C_c_166_n N_VGND_c_568_n 0.00199015f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_163 N_C_c_166_n N_VGND_c_576_n 0.00304119f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B_c_199_n N_A_c_229_n 0.0249402f $X=2.56 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_165 N_B_c_198_n N_A_c_230_n 0.0757342f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B_c_200_n N_A_c_230_n 0.0113106f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_167 N_B_c_198_n A 2.18932e-19 $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_168 N_B_c_200_n A 0.00854992f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_169 N_B_c_198_n N_A_c_231_n 0.00138994f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B_c_200_n N_A_c_231_n 0.0371899f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_171 N_B_c_198_n N_A_225_297#_c_300_n 6.39977e-19 $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B_c_199_n N_A_225_297#_c_300_n 0.01167f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B_c_200_n N_A_225_297#_c_300_n 0.0200207f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B_c_200_n N_A_225_297#_c_307_n 0.00136476f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_175 N_B_c_200_n N_VPWR_c_411_n 0.021614f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_176 N_B_c_198_n N_VPWR_c_415_n 0.00450951f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_177 N_B_c_200_n N_VPWR_c_415_n 0.0118327f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_178 N_B_c_198_n N_VPWR_c_408_n 0.00622433f $X=2.535 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B_c_200_n N_VPWR_c_408_n 0.0111733f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B_c_200_n A_431_297# 0.00821046f $X=2.54 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_181 N_B_c_200_n A_525_297# 0.0113974f $X=2.54 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_182 N_B_c_199_n N_VGND_c_563_n 0.00176556f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B_c_199_n N_VGND_c_570_n 0.00428022f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B_c_199_n N_VGND_c_576_n 0.00585784f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_c_229_n N_A_225_297#_c_267_n 0.0169356f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_c_230_n N_A_225_297#_c_275_n 0.0300561f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_187 A N_A_225_297#_c_275_n 0.00138904f $X=3.155 $Y=1.445 $X2=0 $Y2=0
cc_188 N_A_c_231_n N_A_225_297#_c_275_n 7.11862e-19 $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_c_229_n N_A_225_297#_c_312_n 0.0121804f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_230_n N_A_225_297#_c_312_n 0.00208416f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_191 A N_A_225_297#_c_312_n 0.00494055f $X=3.155 $Y=1.445 $X2=0 $Y2=0
cc_192 N_A_c_231_n N_A_225_297#_c_312_n 0.019282f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_c_229_n N_A_225_297#_c_272_n 0.00323346f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_230_n N_A_225_297#_c_272_n 5.19892e-19 $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_c_231_n N_A_225_297#_c_272_n 0.005931f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_c_230_n N_A_225_297#_c_273_n 0.00127183f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_197 A N_A_225_297#_c_273_n 0.00707041f $X=3.155 $Y=1.445 $X2=0 $Y2=0
cc_198 N_A_c_231_n N_A_225_297#_c_273_n 0.0142427f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_c_230_n N_A_225_297#_c_274_n 0.0187825f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_c_231_n N_A_225_297#_c_274_n 0.00252151f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_201 A N_VPWR_M1001_d 0.00517956f $X=3.155 $Y=1.445 $X2=0 $Y2=0
cc_202 N_A_c_230_n N_VPWR_c_411_n 0.0131142f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_203 A N_VPWR_c_411_n 0.0193325f $X=3.155 $Y=1.445 $X2=0 $Y2=0
cc_204 N_A_c_230_n N_VPWR_c_415_n 0.00702461f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_c_230_n N_VPWR_c_408_n 0.0130026f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_206 A N_X_c_486_n 0.00201115f $X=3.155 $Y=1.445 $X2=0 $Y2=0
cc_207 N_A_c_229_n N_VGND_c_564_n 0.00473127f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_c_229_n N_VGND_c_570_n 0.00428022f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_c_229_n N_VGND_c_576_n 0.00626581f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_225_297#_c_275_n N_VPWR_c_411_n 0.0101706f $X=3.585 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_225_297#_c_276_n N_VPWR_c_412_n 0.00300743f $X=4.055 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_225_297#_c_277_n N_VPWR_c_412_n 0.00300743f $X=4.525 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_225_297#_c_278_n N_VPWR_c_414_n 0.00479105f $X=4.995 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_225_297#_c_279_n N_VPWR_c_415_n 0.0192697f $X=1.25 $Y=2.34 $X2=0
+ $Y2=0
cc_215 N_A_225_297#_c_275_n N_VPWR_c_417_n 0.00702461f $X=3.585 $Y=1.41 $X2=0
+ $Y2=0
cc_216 N_A_225_297#_c_276_n N_VPWR_c_417_n 0.00702461f $X=4.055 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A_225_297#_c_277_n N_VPWR_c_419_n 0.00702461f $X=4.525 $Y=1.41 $X2=0
+ $Y2=0
cc_218 N_A_225_297#_c_278_n N_VPWR_c_419_n 0.00702461f $X=4.995 $Y=1.41 $X2=0
+ $Y2=0
cc_219 N_A_225_297#_M1017_s N_VPWR_c_408_n 0.00218082f $X=1.125 $Y=1.485 $X2=0
+ $Y2=0
cc_220 N_A_225_297#_c_275_n N_VPWR_c_408_n 0.0128986f $X=3.585 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_225_297#_c_276_n N_VPWR_c_408_n 0.0124092f $X=4.055 $Y=1.41 $X2=0
+ $Y2=0
cc_222 N_A_225_297#_c_277_n N_VPWR_c_408_n 0.0124092f $X=4.525 $Y=1.41 $X2=0
+ $Y2=0
cc_223 N_A_225_297#_c_278_n N_VPWR_c_408_n 0.0133474f $X=4.995 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_225_297#_c_279_n N_VPWR_c_408_n 0.0123945f $X=1.25 $Y=2.34 $X2=0
+ $Y2=0
cc_225 N_A_225_297#_c_271_n A_315_297# 0.00634131f $X=1.615 $Y=1.575 $X2=-0.19
+ $Y2=-0.24
cc_226 N_A_225_297#_c_275_n N_X_c_486_n 3.19638e-19 $X=3.585 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A_225_297#_c_341_p N_X_c_486_n 0.0172229f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_225_297#_c_274_n N_X_c_486_n 0.00674235f $X=4.995 $Y=1.202 $X2=0
+ $Y2=0
cc_229 N_A_225_297#_c_267_n N_X_c_495_n 0.00489827f $X=3.56 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_225_297#_c_268_n N_X_c_495_n 0.00766092f $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_225_297#_c_269_n N_X_c_495_n 5.47877e-19 $X=4.5 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_225_297#_c_312_n N_X_c_495_n 0.00459795f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_225_297#_c_276_n N_X_c_487_n 0.0158555f $X=4.055 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A_225_297#_c_277_n N_X_c_487_n 0.0159162f $X=4.525 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_225_297#_c_341_p N_X_c_487_n 0.0406907f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_225_297#_c_274_n N_X_c_487_n 0.00881912f $X=4.995 $Y=1.202 $X2=0
+ $Y2=0
cc_237 N_A_225_297#_c_268_n N_X_c_480_n 0.00901745f $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A_225_297#_c_269_n N_X_c_480_n 0.00895898f $X=4.5 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_225_297#_c_341_p N_X_c_480_n 0.0392656f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_225_297#_c_274_n N_X_c_480_n 0.00345541f $X=4.995 $Y=1.202 $X2=0
+ $Y2=0
cc_241 N_A_225_297#_c_267_n N_X_c_481_n 0.00157721f $X=3.56 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_225_297#_c_268_n N_X_c_481_n 0.00270583f $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_225_297#_c_312_n N_X_c_481_n 0.00715387f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_225_297#_c_272_n N_X_c_481_n 0.00518689f $X=3.43 $Y=1.075 $X2=0 $Y2=0
cc_245 N_A_225_297#_c_341_p N_X_c_481_n 0.0199589f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A_225_297#_c_274_n N_X_c_481_n 0.0033272f $X=4.995 $Y=1.202 $X2=0 $Y2=0
cc_247 N_A_225_297#_c_268_n N_X_c_513_n 5.24597e-19 $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_225_297#_c_269_n N_X_c_513_n 0.00651696f $X=4.5 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_225_297#_c_278_n N_X_c_488_n 0.0186158f $X=4.995 $Y=1.41 $X2=0 $Y2=0
cc_250 N_A_225_297#_c_341_p N_X_c_488_n 0.00405064f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A_225_297#_c_274_n N_X_c_488_n 9.44246e-19 $X=4.995 $Y=1.202 $X2=0
+ $Y2=0
cc_252 N_A_225_297#_c_270_n N_X_c_482_n 0.0138528f $X=5.02 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_225_297#_c_341_p N_X_c_482_n 0.00208021f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_225_297#_c_269_n N_X_c_483_n 0.00119564f $X=4.5 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A_225_297#_c_341_p N_X_c_483_n 0.0304076f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A_225_297#_c_274_n N_X_c_483_n 0.00486271f $X=4.995 $Y=1.202 $X2=0
+ $Y2=0
cc_257 N_A_225_297#_c_341_p N_X_c_489_n 0.0172229f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_225_297#_c_274_n N_X_c_489_n 0.0065364f $X=4.995 $Y=1.202 $X2=0 $Y2=0
cc_259 N_A_225_297#_c_278_n X 0.00174663f $X=4.995 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A_225_297#_c_270_n X 0.0197067f $X=5.02 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_225_297#_c_341_p X 0.0113286f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A_225_297#_c_300_n N_VGND_M1012_d 0.00842454f $X=2.685 $Y=0.74 $X2=0
+ $Y2=0
cc_263 N_A_225_297#_c_312_n N_VGND_M1005_d 0.00762812f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_264 N_A_225_297#_c_272_n N_VGND_M1005_d 7.52091e-19 $X=3.43 $Y=1.075 $X2=0
+ $Y2=0
cc_265 N_A_225_297#_c_291_n N_VGND_c_562_n 0.011573f $X=1.8 $Y=0.49 $X2=0 $Y2=0
cc_266 N_A_225_297#_c_291_n N_VGND_c_563_n 0.0118543f $X=1.8 $Y=0.49 $X2=0 $Y2=0
cc_267 N_A_225_297#_c_300_n N_VGND_c_563_n 0.0214497f $X=2.685 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_225_297#_c_267_n N_VGND_c_564_n 0.00816884f $X=3.56 $Y=0.995 $X2=0
+ $Y2=0
cc_269 N_A_225_297#_c_268_n N_VGND_c_564_n 0.00115121f $X=4.03 $Y=0.995 $X2=0
+ $Y2=0
cc_270 N_A_225_297#_c_312_n N_VGND_c_564_n 0.0252021f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_271 N_A_225_297#_c_268_n N_VGND_c_565_n 0.00379224f $X=4.03 $Y=0.995 $X2=0
+ $Y2=0
cc_272 N_A_225_297#_c_269_n N_VGND_c_565_n 0.00276126f $X=4.5 $Y=0.995 $X2=0
+ $Y2=0
cc_273 N_A_225_297#_c_270_n N_VGND_c_567_n 0.00438629f $X=5.02 $Y=0.995 $X2=0
+ $Y2=0
cc_274 N_A_225_297#_c_291_n N_VGND_c_568_n 0.00852533f $X=1.8 $Y=0.49 $X2=0
+ $Y2=0
cc_275 N_A_225_297#_c_292_n N_VGND_c_568_n 0.00586573f $X=1.885 $Y=0.74 $X2=0
+ $Y2=0
cc_276 N_A_225_297#_c_300_n N_VGND_c_570_n 0.0029785f $X=2.685 $Y=0.74 $X2=0
+ $Y2=0
cc_277 N_A_225_297#_c_391_p N_VGND_c_570_n 0.00846569f $X=2.77 $Y=0.49 $X2=0
+ $Y2=0
cc_278 N_A_225_297#_c_312_n N_VGND_c_570_n 0.0035399f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_279 N_A_225_297#_c_267_n N_VGND_c_572_n 0.00496106f $X=3.56 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_225_297#_c_268_n N_VGND_c_572_n 0.00423334f $X=4.03 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_225_297#_c_269_n N_VGND_c_574_n 0.00423334f $X=4.5 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A_225_297#_c_270_n N_VGND_c_574_n 0.00437852f $X=5.02 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_225_297#_M1014_d N_VGND_c_576_n 0.00454252f $X=1.585 $Y=0.235 $X2=0
+ $Y2=0
cc_284 N_A_225_297#_M1007_d N_VGND_c_576_n 0.00256656f $X=2.635 $Y=0.235 $X2=0
+ $Y2=0
cc_285 N_A_225_297#_c_267_n N_VGND_c_576_n 0.0083553f $X=3.56 $Y=0.995 $X2=0
+ $Y2=0
cc_286 N_A_225_297#_c_268_n N_VGND_c_576_n 0.00613677f $X=4.03 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_225_297#_c_269_n N_VGND_c_576_n 0.00608558f $X=4.5 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_A_225_297#_c_270_n N_VGND_c_576_n 0.00711083f $X=5.02 $Y=0.995 $X2=0
+ $Y2=0
cc_289 N_A_225_297#_c_291_n N_VGND_c_576_n 0.00618681f $X=1.8 $Y=0.49 $X2=0
+ $Y2=0
cc_290 N_A_225_297#_c_300_n N_VGND_c_576_n 0.00691826f $X=2.685 $Y=0.74 $X2=0
+ $Y2=0
cc_291 N_A_225_297#_c_292_n N_VGND_c_576_n 0.0107733f $X=1.885 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_225_297#_c_391_p N_VGND_c_576_n 0.00625722f $X=2.77 $Y=0.49 $X2=0
+ $Y2=0
cc_293 N_A_225_297#_c_312_n N_VGND_c_576_n 0.00878037f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_408_n A_315_297# 0.0143816f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_295 N_VPWR_c_408_n A_431_297# 0.0090262f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_296 N_VPWR_c_408_n A_525_297# 0.00967957f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_297 N_VPWR_c_408_n N_X_M1000_s 0.00370124f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_298 N_VPWR_c_408_n N_X_M1009_s 0.00370124f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_299 N_VPWR_c_417_n N_X_c_530_n 0.0149311f $X=4.165 $Y=2.72 $X2=0 $Y2=0
cc_300 N_VPWR_c_408_n N_X_c_530_n 0.00955092f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_301 N_VPWR_M1004_d N_X_c_487_n 0.00187091f $X=4.145 $Y=1.485 $X2=0 $Y2=0
cc_302 N_VPWR_c_412_n N_X_c_487_n 0.0143191f $X=4.29 $Y=1.96 $X2=0 $Y2=0
cc_303 N_VPWR_c_419_n N_X_c_534_n 0.0149311f $X=5.105 $Y=2.72 $X2=0 $Y2=0
cc_304 N_VPWR_c_408_n N_X_c_534_n 0.00955092f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_305 N_VPWR_M1011_d N_X_c_488_n 0.00301844f $X=5.085 $Y=1.485 $X2=0 $Y2=0
cc_306 N_VPWR_c_414_n N_X_c_488_n 0.0187873f $X=5.23 $Y=1.96 $X2=0 $Y2=0
cc_307 N_X_c_480_n N_VGND_M1010_s 0.00251047f $X=4.545 $Y=0.815 $X2=0 $Y2=0
cc_308 N_X_c_482_n N_VGND_M1016_s 2.28588e-19 $X=5.175 $Y=0.815 $X2=0 $Y2=0
cc_309 N_X_c_485_n N_VGND_M1016_s 0.00344973f $X=5.295 $Y=0.905 $X2=0 $Y2=0
cc_310 N_X_c_495_n N_VGND_c_564_n 0.0140037f $X=3.82 $Y=0.485 $X2=0 $Y2=0
cc_311 N_X_c_495_n N_VGND_c_565_n 0.0177813f $X=3.82 $Y=0.485 $X2=0 $Y2=0
cc_312 N_X_c_480_n N_VGND_c_565_n 0.0127273f $X=4.545 $Y=0.815 $X2=0 $Y2=0
cc_313 N_X_c_485_n N_VGND_c_566_n 0.00165369f $X=5.295 $Y=0.905 $X2=0 $Y2=0
cc_314 N_X_c_482_n N_VGND_c_567_n 0.00177288f $X=5.175 $Y=0.815 $X2=0 $Y2=0
cc_315 N_X_c_485_n N_VGND_c_567_n 0.0120207f $X=5.295 $Y=0.905 $X2=0 $Y2=0
cc_316 N_X_c_495_n N_VGND_c_572_n 0.0153475f $X=3.82 $Y=0.485 $X2=0 $Y2=0
cc_317 N_X_c_480_n N_VGND_c_572_n 0.00266636f $X=4.545 $Y=0.815 $X2=0 $Y2=0
cc_318 N_X_c_480_n N_VGND_c_574_n 0.00198695f $X=4.545 $Y=0.815 $X2=0 $Y2=0
cc_319 N_X_c_513_n N_VGND_c_574_n 0.0231806f $X=4.76 $Y=0.39 $X2=0 $Y2=0
cc_320 N_X_c_482_n N_VGND_c_574_n 0.00254521f $X=5.175 $Y=0.815 $X2=0 $Y2=0
cc_321 N_X_M1002_d N_VGND_c_576_n 0.00607585f $X=3.635 $Y=0.235 $X2=0 $Y2=0
cc_322 N_X_M1015_d N_VGND_c_576_n 0.00304143f $X=4.575 $Y=0.235 $X2=0 $Y2=0
cc_323 N_X_c_495_n N_VGND_c_576_n 0.00940698f $X=3.82 $Y=0.485 $X2=0 $Y2=0
cc_324 N_X_c_480_n N_VGND_c_576_n 0.00972452f $X=4.545 $Y=0.815 $X2=0 $Y2=0
cc_325 N_X_c_513_n N_VGND_c_576_n 0.0143352f $X=4.76 $Y=0.39 $X2=0 $Y2=0
cc_326 N_X_c_482_n N_VGND_c_576_n 0.00509281f $X=5.175 $Y=0.815 $X2=0 $Y2=0
cc_327 N_X_c_485_n N_VGND_c_576_n 0.00345847f $X=5.295 $Y=0.905 $X2=0 $Y2=0
