# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.070000 0.940000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.070000 0.330000 1.615000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.240000 1.075000 4.950000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.315000 1.075000 6.295000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.368000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.185000 0.655000 2.630000 1.445000 ;
        RECT 2.185000 1.445000 5.875000 1.665000 ;
        RECT 2.185000 1.665000 2.485000 2.465000 ;
        RECT 3.125000 1.665000 3.505000 2.465000 ;
        RECT 3.495000 1.075000 4.045000 1.445000 ;
        RECT 4.555000 1.665000 4.935000 2.465000 ;
        RECT 5.495000 1.665000 5.875000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.440000 0.085000 ;
        RECT 0.515000  0.085000 0.815000 0.545000 ;
        RECT 5.625000  0.085000 5.795000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.440000 2.805000 ;
        RECT 0.540000 2.195000 0.815000 2.635000 ;
        RECT 1.845000 1.495000 2.015000 2.635000 ;
        RECT 2.655000 1.835000 2.955000 2.635000 ;
        RECT 3.725000 1.835000 4.385000 2.635000 ;
        RECT 5.155000 1.835000 5.325000 2.635000 ;
        RECT 6.095000 1.445000 6.345000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 0.345000 0.730000 ;
      RECT 0.085000 0.730000 1.330000 0.900000 ;
      RECT 0.085000 1.785000 1.330000 1.980000 ;
      RECT 0.085000 1.980000 0.370000 2.440000 ;
      RECT 0.985000 0.255000 1.675000 0.560000 ;
      RECT 0.985000 2.150000 1.675000 2.465000 ;
      RECT 1.160000 0.900000 1.330000 1.785000 ;
      RECT 1.500000 0.560000 1.675000 2.150000 ;
      RECT 1.845000 0.255000 3.975000 0.485000 ;
      RECT 1.845000 0.485000 2.015000 0.585000 ;
      RECT 2.945000 1.075000 3.325000 1.275000 ;
      RECT 3.125000 0.655000 4.935000 0.905000 ;
      RECT 4.165000 0.255000 5.405000 0.485000 ;
      RECT 5.155000 0.485000 5.405000 0.735000 ;
      RECT 5.155000 0.735000 6.345000 0.905000 ;
      RECT 5.965000 0.255000 6.345000 0.735000 ;
    LAYER mcon ;
      RECT 1.160000 1.105000 1.330000 1.275000 ;
      RECT 3.155000 1.105000 3.325000 1.275000 ;
    LAYER met1 ;
      RECT 1.100000 1.075000 3.385000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4bb_2
