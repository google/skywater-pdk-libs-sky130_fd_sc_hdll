* File: sky130_fd_sc_hdll__nor2_2.pex.spice
* Created: Thu Aug 27 19:15:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR2_2%A 1 3 4 6 7 9 10 12 13 14 22
c36 14 0 1.09908e-19 $X=0.6 $Y=1.11
c37 7 0 1.24829e-19 $X=0.985 $Y=1.41
r38 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.01 $Y2=1.202
r39 20 22 43.1263 $w=3.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.645 $Y=1.202
+ $X2=0.985 $Y2=1.202
r40 18 20 16.4895 $w=3.8e-07 $l=1.3e-07 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.645 $Y2=1.202
r41 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r42 14 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r43 13 14 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.645 $Y2=1.175
r44 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.202
r45 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r46 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r47 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r48 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r49 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r50 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_2%B 1 3 4 6 7 9 10 12 13 14 22
c48 22 0 1.09908e-19 $X=1.925 $Y=1.202
r49 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r50 20 22 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=1.69 $Y=1.202
+ $X2=1.925 $Y2=1.202
r51 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.69 $Y2=1.202
r52 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r53 14 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.16 $X2=1.69 $Y2=1.16
r54 13 14 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.605 $Y2=1.175
r55 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r56 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r57 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r58 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r59 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r60 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r61 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995 $X2=1.43
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_2%A_27_297# 1 2 3 10 12 14 16 17 18 22
r39 20 22 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=2.225 $Y=2.295
+ $X2=2.225 $Y2=2
r40 19 29 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=2.38
+ $X2=1.22 $Y2=2.38
r41 18 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.075 $Y=2.38
+ $X2=2.225 $Y2=2.295
r42 18 19 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.075 $Y=2.38
+ $X2=1.305 $Y2=2.38
r43 17 29 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.295
+ $X2=1.22 $Y2=2.38
r44 16 27 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.56
r45 16 17 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=2.295
r46 15 25 3.96222 $w=2.1e-07 $l=1.38e-07 $layer=LI1_cond $X=0.365 $Y=1.56
+ $X2=0.227 $Y2=1.56
r47 14 27 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=1.56
+ $X2=1.22 $Y2=1.56
r48 14 15 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=1.56
+ $X2=0.365 $Y2=1.56
r49 10 25 3.01473 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=0.227 $Y=1.665
+ $X2=0.227 $Y2=1.56
r50 10 12 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=0.227 $Y=1.665
+ $X2=0.227 $Y2=2.3
r51 3 22 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2
r52 2 29 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r53 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r54 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r55 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_2%VPWR 1 6 8 10 20 21 24
r31 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r32 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r33 18 21 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r34 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r35 17 20 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r37 15 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=0.725 $Y2=2.72
r38 15 17 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r39 10 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.725 $Y2=2.72
r40 10 12 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r41 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r43 4 24 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=2.72
r44 4 6 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=2
r45 1 6 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_2%Y 1 2 3 12 14 15 18 20 22 25 26 27 30
c61 27 0 1.24829e-19 $X=1.665 $Y=1.665
r62 27 30 6.21713 $w=3.78e-07 $l=2.05e-07 $layer=LI1_cond $X=1.665 $Y=1.665
+ $X2=1.665 $Y2=1.87
r63 27 29 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.665 $Y=1.665
+ $X2=1.665 $Y2=1.555
r64 24 25 28.9451 $w=2.13e-07 $l=5.4e-07 $layer=LI1_cond $X=2.202 $Y=0.905
+ $X2=2.202 $Y2=1.445
r65 23 29 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=1.555
+ $X2=1.665 $Y2=1.555
r66 22 25 6.81766 $w=2.2e-07 $l=1.54499e-07 $layer=LI1_cond $X=2.095 $Y=1.555
+ $X2=2.202 $Y2=1.445
r67 22 23 12.5721 $w=2.18e-07 $l=2.4e-07 $layer=LI1_cond $X=2.095 $Y=1.555
+ $X2=1.855 $Y2=1.555
r68 21 26 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=1.855 $Y=0.82
+ $X2=1.665 $Y2=0.815
r69 20 24 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=2.095 $Y=0.82
+ $X2=2.202 $Y2=0.905
r70 20 21 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.095 $Y=0.82
+ $X2=1.855 $Y2=0.82
r71 16 26 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.815
r72 16 18 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.39
r73 14 26 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=1.665 $Y2=0.815
r74 14 15 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=0.915 $Y2=0.815
r75 10 15 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.815
r76 10 12 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r77 3 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.62
r78 2 18 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r79 1 12 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_2%VGND 1 2 3 10 12 14 18 22 24 25 26 27 35 40
r39 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r40 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r41 32 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r42 32 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r43 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r44 29 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r45 29 31 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=2.07
+ $Y2=0
r46 27 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r47 27 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r48 25 31 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.07
+ $Y2=0
r49 25 26 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.31
+ $Y2=0
r50 24 34 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.53
+ $Y2=0
r51 24 26 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.31
+ $Y2=0
r52 20 26 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=0.085
+ $X2=2.31 $Y2=0
r53 20 22 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=2.31 $Y=0.085
+ $X2=2.31 $Y2=0.39
r54 16 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r55 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r56 15 37 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r57 14 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r58 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.365
+ $Y2=0
r59 10 37 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r60 10 12 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r61 3 22 182 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.275 $Y2=0.39
r62 2 18 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
r63 1 12 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

