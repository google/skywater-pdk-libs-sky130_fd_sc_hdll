* File: sky130_fd_sc_hdll__o2bb2ai_4.pxi.spice
* Created: Thu Aug 27 19:22:18 2020
* 
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A2_N N_A2_N_c_156_n N_A2_N_M1003_g
+ N_A2_N_c_162_n N_A2_N_M1002_g N_A2_N_c_157_n N_A2_N_M1021_g N_A2_N_c_163_n
+ N_A2_N_M1010_g N_A2_N_c_158_n N_A2_N_M1022_g N_A2_N_c_164_n N_A2_N_M1018_g
+ N_A2_N_c_165_n N_A2_N_M1029_g N_A2_N_c_159_n N_A2_N_M1037_g A2_N
+ N_A2_N_c_160_n N_A2_N_c_161_n A2_N PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A2_N
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A1_N N_A1_N_c_221_n N_A1_N_M1015_g
+ N_A1_N_c_227_n N_A1_N_M1001_g N_A1_N_c_222_n N_A1_N_M1017_g N_A1_N_c_228_n
+ N_A1_N_M1023_g N_A1_N_c_223_n N_A1_N_M1031_g N_A1_N_c_229_n N_A1_N_M1035_g
+ N_A1_N_c_230_n N_A1_N_M1039_g N_A1_N_c_224_n N_A1_N_M1038_g A1_N
+ N_A1_N_c_225_n N_A1_N_c_226_n A1_N PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A1_N
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_113_47# N_A_113_47#_M1003_s
+ N_A_113_47#_M1022_s N_A_113_47#_M1002_d N_A_113_47#_M1018_d
+ N_A_113_47#_M1001_d N_A_113_47#_M1035_d N_A_113_47#_c_313_n
+ N_A_113_47#_M1004_g N_A_113_47#_c_302_n N_A_113_47#_M1006_g
+ N_A_113_47#_c_314_n N_A_113_47#_M1007_g N_A_113_47#_c_303_n
+ N_A_113_47#_M1008_g N_A_113_47#_c_315_n N_A_113_47#_M1019_g
+ N_A_113_47#_c_304_n N_A_113_47#_M1028_g N_A_113_47#_c_316_n
+ N_A_113_47#_M1036_g N_A_113_47#_c_305_n N_A_113_47#_M1033_g
+ N_A_113_47#_c_306_n N_A_113_47#_c_307_n N_A_113_47#_c_308_n
+ N_A_113_47#_c_318_n N_A_113_47#_c_319_n N_A_113_47#_c_379_p
+ N_A_113_47#_c_320_n N_A_113_47#_c_381_p N_A_113_47#_c_321_n
+ N_A_113_47#_c_383_p N_A_113_47#_c_322_n N_A_113_47#_c_395_p
+ N_A_113_47#_c_323_n N_A_113_47#_c_309_n N_A_113_47#_c_310_n
+ N_A_113_47#_c_311_n N_A_113_47#_c_325_n N_A_113_47#_c_326_n
+ N_A_113_47#_c_327_n N_A_113_47#_c_328_n N_A_113_47#_c_312_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_113_47#
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%B2 N_B2_c_464_n N_B2_M1000_g N_B2_c_470_n
+ N_B2_M1011_g N_B2_c_465_n N_B2_M1013_g N_B2_c_471_n N_B2_M1024_g N_B2_c_466_n
+ N_B2_M1016_g N_B2_c_472_n N_B2_M1030_g N_B2_c_473_n N_B2_M1032_g N_B2_c_467_n
+ N_B2_M1034_g B2 N_B2_c_468_n N_B2_c_469_n B2
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_4%B2
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%B1 N_B1_c_549_n N_B1_M1009_g N_B1_c_555_n
+ N_B1_M1005_g N_B1_c_550_n N_B1_M1012_g N_B1_c_556_n N_B1_M1014_g N_B1_c_551_n
+ N_B1_M1026_g N_B1_c_557_n N_B1_M1020_g N_B1_c_558_n N_B1_M1025_g N_B1_c_552_n
+ N_B1_M1027_g B1 N_B1_c_553_n N_B1_c_554_n B1
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_4%B1
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%VPWR N_VPWR_M1002_s N_VPWR_M1010_s
+ N_VPWR_M1029_s N_VPWR_M1023_s N_VPWR_M1039_s N_VPWR_M1007_d N_VPWR_M1036_d
+ N_VPWR_M1005_d N_VPWR_M1020_d N_VPWR_c_625_n N_VPWR_c_626_n N_VPWR_c_627_n
+ N_VPWR_c_628_n N_VPWR_c_629_n N_VPWR_c_630_n N_VPWR_c_631_n N_VPWR_c_632_n
+ N_VPWR_c_633_n N_VPWR_c_634_n N_VPWR_c_635_n N_VPWR_c_636_n N_VPWR_c_637_n
+ N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_640_n N_VPWR_c_641_n N_VPWR_c_642_n
+ N_VPWR_c_643_n N_VPWR_c_644_n N_VPWR_c_645_n VPWR N_VPWR_c_646_n
+ N_VPWR_c_647_n N_VPWR_c_624_n N_VPWR_c_649_n N_VPWR_c_650_n N_VPWR_c_651_n
+ N_VPWR_c_652_n VPWR PM_SKY130_FD_SC_HDLL__O2BB2AI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%Y N_Y_M1006_d N_Y_M1028_d N_Y_M1004_s
+ N_Y_M1019_s N_Y_M1011_d N_Y_M1030_d N_Y_c_774_n N_Y_c_776_n N_Y_c_829_n
+ N_Y_c_777_n N_Y_c_833_n N_Y_c_778_n N_Y_c_779_n N_Y_c_780_n N_Y_c_781_n
+ N_Y_c_782_n N_Y_c_783_n Y PM_SKY130_FD_SC_HDLL__O2BB2AI_4%Y
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_1361_297# N_A_1361_297#_M1011_s
+ N_A_1361_297#_M1024_s N_A_1361_297#_M1032_s N_A_1361_297#_M1014_s
+ N_A_1361_297#_M1025_s N_A_1361_297#_c_863_n N_A_1361_297#_c_871_n
+ N_A_1361_297#_c_864_n N_A_1361_297#_c_921_n N_A_1361_297#_c_873_n
+ N_A_1361_297#_c_865_n N_A_1361_297#_c_901_n N_A_1361_297#_c_866_n
+ N_A_1361_297#_c_905_n N_A_1361_297#_c_867_n N_A_1361_297#_c_868_n
+ N_A_1361_297#_c_869_n N_A_1361_297#_c_911_n N_A_1361_297#_c_870_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_1361_297#
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_27_47# N_A_27_47#_M1003_d N_A_27_47#_M1021_d
+ N_A_27_47#_M1037_d N_A_27_47#_M1017_s N_A_27_47#_M1038_s N_A_27_47#_c_927_n
+ N_A_27_47#_c_938_n N_A_27_47#_c_928_n N_A_27_47#_c_929_n N_A_27_47#_c_946_n
+ N_A_27_47#_c_930_n N_A_27_47#_c_931_n N_A_27_47#_c_932_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%VGND N_VGND_M1015_d N_VGND_M1031_d
+ N_VGND_M1000_d N_VGND_M1016_d N_VGND_M1009_d N_VGND_M1026_d N_VGND_c_1004_n
+ N_VGND_c_1005_n N_VGND_c_1006_n N_VGND_c_1007_n N_VGND_c_1008_n
+ N_VGND_c_1009_n N_VGND_c_1010_n N_VGND_c_1011_n N_VGND_c_1012_n
+ N_VGND_c_1013_n N_VGND_c_1014_n N_VGND_c_1015_n N_VGND_c_1016_n
+ N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n N_VGND_c_1020_n
+ N_VGND_c_1021_n VGND N_VGND_c_1022_n N_VGND_c_1023_n VGND
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_4%VGND
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_887_47# N_A_887_47#_M1006_s
+ N_A_887_47#_M1008_s N_A_887_47#_M1033_s N_A_887_47#_M1013_s
+ N_A_887_47#_M1034_s N_A_887_47#_M1012_s N_A_887_47#_M1027_s
+ N_A_887_47#_c_1164_n N_A_887_47#_c_1165_n N_A_887_47#_c_1230_n
+ N_A_887_47#_c_1170_n N_A_887_47#_c_1155_n N_A_887_47#_c_1156_n
+ N_A_887_47#_c_1181_n N_A_887_47#_c_1157_n N_A_887_47#_c_1189_n
+ N_A_887_47#_c_1158_n N_A_887_47#_c_1203_n N_A_887_47#_c_1159_n
+ N_A_887_47#_c_1160_n N_A_887_47#_c_1161_n N_A_887_47#_c_1162_n
+ N_A_887_47#_c_1163_n PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_887_47#
cc_1 VNB N_A2_N_c_156_n 0.0197108f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A2_N_c_157_n 0.0167462f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_3 VNB N_A2_N_c_158_n 0.017207f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_4 VNB N_A2_N_c_159_n 0.0171597f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_5 VNB N_A2_N_c_160_n 0.00156728f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=1.16
cc_6 VNB N_A2_N_c_161_n 0.0766663f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_7 VNB N_A1_N_c_221_n 0.0164797f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_A1_N_c_222_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_9 VNB N_A1_N_c_223_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_10 VNB N_A1_N_c_224_n 0.0223965f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_11 VNB N_A1_N_c_225_n 0.00378123f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=1.16
cc_12 VNB N_A1_N_c_226_n 0.0795575f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_13 VNB N_A_113_47#_c_302_n 0.0220755f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_14 VNB N_A_113_47#_c_303_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_15 VNB N_A_113_47#_c_304_n 0.0171839f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=1.202
cc_16 VNB N_A_113_47#_c_305_n 0.0201615f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.202
cc_17 VNB N_A_113_47#_c_306_n 0.0190508f $X=-0.19 $Y=-0.24 $X2=1.14 $Y2=1.19
cc_18 VNB N_A_113_47#_c_307_n 0.0116419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_113_47#_c_308_n 0.00988729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_113_47#_c_309_n 5.22495e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_113_47#_c_310_n 0.00772394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_113_47#_c_311_n 0.0159479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_113_47#_c_312_n 0.0855028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_B2_c_464_n 0.0198703f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_25 VNB N_B2_c_465_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_26 VNB N_B2_c_466_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_27 VNB N_B2_c_467_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_28 VNB N_B2_c_468_n 0.0036326f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=1.16
cc_29 VNB N_B2_c_469_n 0.0773639f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_30 VNB N_B1_c_549_n 0.0164927f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_31 VNB N_B1_c_550_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_32 VNB N_B1_c_551_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_33 VNB N_B1_c_552_n 0.0223965f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_34 VNB N_B1_c_553_n 0.0241581f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=1.16
cc_35 VNB N_B1_c_554_n 0.0801709f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_36 VNB N_VPWR_c_624_n 0.459507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_774_n 0.0104258f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_38 VNB Y 0.0116109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_27_47#_c_927_n 0.00973351f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_40 VNB N_A_27_47#_c_928_n 0.00357343f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_41 VNB N_A_27_47#_c_929_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_42 VNB N_A_27_47#_c_930_n 0.00916719f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_43 VNB N_A_27_47#_c_931_n 0.00482775f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=1.202
cc_44 VNB N_A_27_47#_c_932_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.202
cc_45 VNB N_VGND_c_1004_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.985
cc_46 VNB N_VGND_c_1005_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.105
cc_47 VNB N_VGND_c_1006_n 0.00463499f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.202
cc_48 VNB N_VGND_c_1007_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_49 VNB N_VGND_c_1008_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=1.16
cc_50 VNB N_VGND_c_1009_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.18
cc_51 VNB N_VGND_c_1010_n 0.060673f $X=-0.19 $Y=-0.24 $X2=1.14 $Y2=1.19
cc_52 VNB N_VGND_c_1011_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1012_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=1.18
cc_54 VNB N_VGND_c_1013_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1014_n 0.085512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1015_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1016_n 0.019187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1017_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1018_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1019_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1020_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1021_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1022_n 0.0211936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1023_n 0.51896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_887_47#_c_1155_n 0.00247032f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=1.202
cc_66 VNB N_A_887_47#_c_1156_n 0.00155757f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.202
cc_67 VNB N_A_887_47#_c_1157_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.202
cc_68 VNB N_A_887_47#_c_1158_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.24 $Y2=1.18
cc_69 VNB N_A_887_47#_c_1159_n 0.0132268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_887_47#_c_1160_n 0.0187437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_887_47#_c_1161_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_887_47#_c_1162_n 0.00384439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_887_47#_c_1163_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VPB N_A2_N_c_162_n 0.019185f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_75 VPB N_A2_N_c_163_n 0.0159561f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_76 VPB N_A2_N_c_164_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_77 VPB N_A2_N_c_165_n 0.0161064f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_78 VPB N_A2_N_c_161_n 0.0456213f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_79 VPB N_A1_N_c_227_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_80 VPB N_A1_N_c_228_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_81 VPB N_A1_N_c_229_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_82 VPB N_A1_N_c_230_n 0.0192379f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_83 VPB N_A1_N_c_226_n 0.045749f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_84 VPB N_A_113_47#_c_313_n 0.0194469f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_85 VPB N_A_113_47#_c_314_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.105
cc_86 VPB N_A_113_47#_c_315_n 0.0159563f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_87 VPB N_A_113_47#_c_316_n 0.0192098f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=1.16
cc_88 VPB N_A_113_47#_c_306_n 0.00741836f $X=-0.19 $Y=1.305 $X2=1.14 $Y2=1.19
cc_89 VPB N_A_113_47#_c_318_n 0.00231882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_113_47#_c_319_n 0.00935576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_113_47#_c_320_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_113_47#_c_321_n 0.00539591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_113_47#_c_322_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_113_47#_c_323_n 0.00437675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_113_47#_c_309_n 0.0041058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_113_47#_c_325_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_113_47#_c_326_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_113_47#_c_327_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_113_47#_c_328_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_113_47#_c_312_n 0.0481798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_B2_c_470_n 0.019253f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_102 VPB N_B2_c_471_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_103 VPB N_B2_c_472_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_104 VPB N_B2_c_473_n 0.0164231f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_105 VPB N_B2_c_469_n 0.046689f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_106 VPB N_B1_c_555_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_107 VPB N_B1_c_556_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_108 VPB N_B1_c_557_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_109 VPB N_B1_c_558_n 0.0203443f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_110 VPB N_B1_c_554_n 0.048391f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_111 VPB N_VPWR_c_625_n 0.011928f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_112 VPB N_VPWR_c_626_n 0.00518f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_113 VPB N_VPWR_c_627_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.202
cc_114 VPB N_VPWR_c_628_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=1.202
cc_115 VPB N_VPWR_c_629_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=1.16
cc_116 VPB N_VPWR_c_630_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_631_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.14 $Y2=1.19
cc_118 VPB N_VPWR_c_632_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_633_n 0.00789678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_634_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_635_n 0.00518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_636_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_637_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_638_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_639_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_640_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_641_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_642_n 0.0624384f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_643_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_644_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_645_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_646_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_647_n 0.021362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_624_n 0.0594653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_649_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_650_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_651_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_652_n 0.0142078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_Y_c_776_n 0.00184257f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.105
cc_140 VPB N_Y_c_777_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.202
cc_141 VPB N_Y_c_778_n 0.00263282f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.202
cc_142 VPB N_Y_c_779_n 0.00743367f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=1.16
cc_143 VPB N_Y_c_780_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.18
cc_144 VPB N_Y_c_781_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_Y_c_782_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_Y_c_783_n 0.00174485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB Y 0.0168489f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_1361_297#_c_863_n 0.00486153f $X=-0.19 $Y=1.305 $X2=1.455
+ $Y2=1.985
cc_149 VPB N_A_1361_297#_c_864_n 0.00179668f $X=-0.19 $Y=1.305 $X2=1.925
+ $Y2=1.985
cc_150 VPB N_A_1361_297#_c_865_n 0.00359595f $X=-0.19 $Y=1.305 $X2=0.515
+ $Y2=1.202
cc_151 VPB N_A_1361_297#_c_866_n 0.00196267f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_152 VPB N_A_1361_297#_c_867_n 0.00196267f $X=-0.19 $Y=1.305 $X2=1.76
+ $Y2=1.202
cc_153 VPB N_A_1361_297#_c_868_n 0.010205f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=1.16
cc_154 VPB N_A_1361_297#_c_869_n 0.032524f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=1.202
cc_155 VPB N_A_1361_297#_c_870_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 N_A2_N_c_159_n N_A1_N_c_221_n 0.0175316f $X=1.95 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_157 N_A2_N_c_165_n N_A1_N_c_227_n 0.0216822f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A2_N_c_160_n N_A1_N_c_225_n 0.0121231f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_N_c_161_n N_A1_N_c_225_n 2.62535e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_160 N_A2_N_c_160_n N_A1_N_c_226_n 2.62535e-19 $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A2_N_c_161_n N_A1_N_c_226_n 0.0175316f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_162 N_A2_N_c_156_n N_A_113_47#_c_306_n 0.0167836f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A2_N_c_162_n N_A_113_47#_c_306_n 0.00153799f $X=0.515 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A2_N_c_160_n N_A_113_47#_c_306_n 0.0166223f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A2_N_c_156_n N_A_113_47#_c_308_n 0.0134143f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A2_N_c_157_n N_A_113_47#_c_308_n 0.0114491f $X=0.96 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A2_N_c_158_n N_A_113_47#_c_308_n 0.0114446f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_168 N_A2_N_c_159_n N_A_113_47#_c_308_n 2.03781e-19 $X=1.95 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A2_N_c_160_n N_A_113_47#_c_308_n 0.105727f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A2_N_c_161_n N_A_113_47#_c_308_n 0.0117089f $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_171 N_A2_N_c_162_n N_A_113_47#_c_318_n 0.0170402f $X=0.515 $Y=1.41 $X2=0
+ $Y2=0
cc_172 N_A2_N_c_160_n N_A_113_47#_c_318_n 0.0138171f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A2_N_c_161_n N_A_113_47#_c_318_n 9.33689e-19 $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_174 N_A2_N_c_163_n N_A_113_47#_c_320_n 0.0156273f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_175 N_A2_N_c_164_n N_A_113_47#_c_320_n 0.0156273f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A2_N_c_160_n N_A_113_47#_c_320_n 0.0486996f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A2_N_c_161_n N_A_113_47#_c_320_n 0.00864922f $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_178 N_A2_N_c_165_n N_A_113_47#_c_321_n 0.0155843f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_179 N_A2_N_c_160_n N_A_113_47#_c_321_n 0.0145434f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A2_N_c_161_n N_A_113_47#_c_321_n 8.84531e-19 $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_181 N_A2_N_c_160_n N_A_113_47#_c_325_n 0.0204509f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A2_N_c_161_n N_A_113_47#_c_325_n 0.00656533f $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_183 N_A2_N_c_160_n N_A_113_47#_c_326_n 0.0204509f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A2_N_c_161_n N_A_113_47#_c_326_n 0.00635938f $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_185 N_A2_N_c_162_n N_VPWR_c_626_n 0.00479105f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A2_N_c_162_n N_VPWR_c_627_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A2_N_c_163_n N_VPWR_c_627_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A2_N_c_163_n N_VPWR_c_628_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A2_N_c_164_n N_VPWR_c_628_n 0.00300743f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A2_N_c_164_n N_VPWR_c_629_n 0.00702461f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A2_N_c_165_n N_VPWR_c_629_n 0.00702461f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A2_N_c_165_n N_VPWR_c_630_n 0.00300743f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A2_N_c_162_n N_VPWR_c_624_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A2_N_c_163_n N_VPWR_c_624_n 0.0124092f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A2_N_c_164_n N_VPWR_c_624_n 0.0124092f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A2_N_c_165_n N_VPWR_c_624_n 0.0124344f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A2_N_c_156_n N_A_27_47#_c_927_n 0.00931157f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A2_N_c_157_n N_A_27_47#_c_927_n 0.00931157f $X=0.96 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A2_N_c_158_n N_A_27_47#_c_927_n 0.00964761f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A2_N_c_159_n N_A_27_47#_c_927_n 0.0117007f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A2_N_c_160_n N_A_27_47#_c_927_n 0.0039487f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A2_N_c_156_n N_VGND_c_1010_n 0.00357877f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A2_N_c_157_n N_VGND_c_1010_n 0.00357877f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A2_N_c_158_n N_VGND_c_1010_n 0.00357877f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A2_N_c_159_n N_VGND_c_1010_n 0.00357877f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A2_N_c_156_n N_VGND_c_1023_n 0.0063299f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A2_N_c_157_n N_VGND_c_1023_n 0.00548399f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A2_N_c_158_n N_VGND_c_1023_n 0.00560377f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A2_N_c_159_n N_VGND_c_1023_n 0.005504f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A1_N_c_227_n N_A_113_47#_c_321_n 0.0155843f $X=2.395 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A1_N_c_225_n N_A_113_47#_c_321_n 0.0145434f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A1_N_c_226_n N_A_113_47#_c_321_n 8.84531e-19 $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_213 N_A1_N_c_228_n N_A_113_47#_c_322_n 0.0156273f $X=2.865 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A1_N_c_229_n N_A_113_47#_c_322_n 0.0156273f $X=3.335 $Y=1.41 $X2=0
+ $Y2=0
cc_215 N_A1_N_c_225_n N_A_113_47#_c_322_n 0.0486996f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A1_N_c_226_n N_A_113_47#_c_322_n 0.00864922f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_217 N_A1_N_c_230_n N_A_113_47#_c_323_n 0.0172094f $X=3.805 $Y=1.41 $X2=0
+ $Y2=0
cc_218 N_A1_N_c_225_n N_A_113_47#_c_323_n 0.0145434f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A1_N_c_226_n N_A_113_47#_c_323_n 8.84531e-19 $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_220 N_A1_N_c_230_n N_A_113_47#_c_309_n 0.00141146f $X=3.805 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A1_N_c_226_n N_A_113_47#_c_309_n 0.00431362f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_222 N_A1_N_c_225_n N_A_113_47#_c_310_n 0.0143012f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A1_N_c_226_n N_A_113_47#_c_310_n 0.00156252f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_224 N_A1_N_c_225_n N_A_113_47#_c_327_n 0.0204509f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A1_N_c_226_n N_A_113_47#_c_327_n 0.00656533f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_226 N_A1_N_c_225_n N_A_113_47#_c_328_n 0.0204509f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A1_N_c_226_n N_A_113_47#_c_328_n 0.00635938f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_228 N_A1_N_c_227_n N_VPWR_c_630_n 0.00300743f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A1_N_c_227_n N_VPWR_c_631_n 0.00702461f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A1_N_c_228_n N_VPWR_c_631_n 0.00702461f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A1_N_c_228_n N_VPWR_c_632_n 0.00300743f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A1_N_c_229_n N_VPWR_c_632_n 0.00300743f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A1_N_c_230_n N_VPWR_c_633_n 0.00513552f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A1_N_c_229_n N_VPWR_c_646_n 0.00702461f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A1_N_c_230_n N_VPWR_c_646_n 0.00702461f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A1_N_c_227_n N_VPWR_c_624_n 0.0124344f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A1_N_c_228_n N_VPWR_c_624_n 0.0124092f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_238 N_A1_N_c_229_n N_VPWR_c_624_n 0.0124092f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A1_N_c_230_n N_VPWR_c_624_n 0.0136915f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A1_N_c_221_n N_A_27_47#_c_938_n 0.00282739f $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A1_N_c_221_n N_A_27_47#_c_928_n 0.00513032f $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A1_N_c_222_n N_A_27_47#_c_928_n 4.74935e-19 $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A1_N_c_225_n N_A_27_47#_c_928_n 0.00231036f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A1_N_c_221_n N_A_27_47#_c_929_n 0.00901745f $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A1_N_c_222_n N_A_27_47#_c_929_n 0.00895898f $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A1_N_c_225_n N_A_27_47#_c_929_n 0.0398926f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A1_N_c_226_n N_A_27_47#_c_929_n 0.00345541f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_248 N_A1_N_c_221_n N_A_27_47#_c_946_n 5.24597e-19 $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_A1_N_c_222_n N_A_27_47#_c_946_n 0.00651696f $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_A1_N_c_223_n N_A_27_47#_c_946_n 0.00693563f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A1_N_c_224_n N_A_27_47#_c_946_n 5.34196e-19 $X=3.83 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A1_N_c_223_n N_A_27_47#_c_930_n 0.00929182f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A1_N_c_224_n N_A_27_47#_c_930_n 0.00936658f $X=3.83 $Y=0.995 $X2=0
+ $Y2=0
cc_254 N_A1_N_c_225_n N_A_27_47#_c_930_n 0.0462421f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A1_N_c_226_n N_A_27_47#_c_930_n 0.00468948f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_256 N_A1_N_c_223_n N_A_27_47#_c_931_n 5.69266e-19 $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_A1_N_c_224_n N_A_27_47#_c_931_n 0.00857123f $X=3.83 $Y=0.995 $X2=0
+ $Y2=0
cc_258 N_A1_N_c_222_n N_A_27_47#_c_932_n 0.00116636f $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A1_N_c_223_n N_A_27_47#_c_932_n 0.00116636f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_A1_N_c_225_n N_A_27_47#_c_932_n 0.0307014f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A1_N_c_226_n N_A_27_47#_c_932_n 0.00358305f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_262 N_A1_N_c_221_n N_VGND_c_1004_n 0.00378935f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A1_N_c_222_n N_VGND_c_1004_n 0.00276126f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A1_N_c_223_n N_VGND_c_1005_n 0.00385467f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A1_N_c_224_n N_VGND_c_1005_n 0.00365402f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A1_N_c_221_n N_VGND_c_1010_n 0.00421816f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A1_N_c_222_n N_VGND_c_1012_n 0.00423334f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A1_N_c_223_n N_VGND_c_1012_n 0.00423334f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A1_N_c_224_n N_VGND_c_1014_n 0.00396605f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A1_N_c_221_n N_VGND_c_1023_n 0.00600232f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A1_N_c_222_n N_VGND_c_1023_n 0.00597024f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A1_N_c_223_n N_VGND_c_1023_n 0.00620835f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A1_N_c_224_n N_VGND_c_1023_n 0.00712929f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_113_47#_c_318_n N_VPWR_M1002_s 0.00119058f $X=0.625 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_275 N_A_113_47#_c_319_n N_VPWR_M1002_s 0.00289527f $X=0.255 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_276 N_A_113_47#_c_320_n N_VPWR_M1010_s 0.00187091f $X=1.565 $Y=1.54 $X2=0
+ $Y2=0
cc_277 N_A_113_47#_c_321_n N_VPWR_M1029_s 0.00187091f $X=2.505 $Y=1.54 $X2=0
+ $Y2=0
cc_278 N_A_113_47#_c_322_n N_VPWR_M1023_s 0.00187091f $X=3.445 $Y=1.54 $X2=0
+ $Y2=0
cc_279 N_A_113_47#_c_323_n N_VPWR_M1039_s 0.00796532f $X=4.145 $Y=1.54 $X2=0
+ $Y2=0
cc_280 N_A_113_47#_c_318_n N_VPWR_c_626_n 0.00915704f $X=0.625 $Y=1.54 $X2=0
+ $Y2=0
cc_281 N_A_113_47#_c_319_n N_VPWR_c_626_n 0.00892602f $X=0.255 $Y=1.54 $X2=0
+ $Y2=0
cc_282 N_A_113_47#_c_379_p N_VPWR_c_627_n 0.0149311f $X=0.75 $Y=2.3 $X2=0 $Y2=0
cc_283 N_A_113_47#_c_320_n N_VPWR_c_628_n 0.0143191f $X=1.565 $Y=1.54 $X2=0
+ $Y2=0
cc_284 N_A_113_47#_c_381_p N_VPWR_c_629_n 0.0149311f $X=1.69 $Y=2.3 $X2=0 $Y2=0
cc_285 N_A_113_47#_c_321_n N_VPWR_c_630_n 0.0143191f $X=2.505 $Y=1.54 $X2=0
+ $Y2=0
cc_286 N_A_113_47#_c_383_p N_VPWR_c_631_n 0.0149311f $X=2.63 $Y=2.3 $X2=0 $Y2=0
cc_287 N_A_113_47#_c_322_n N_VPWR_c_632_n 0.0143191f $X=3.445 $Y=1.54 $X2=0
+ $Y2=0
cc_288 N_A_113_47#_c_313_n N_VPWR_c_633_n 0.00513552f $X=4.765 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_113_47#_c_323_n N_VPWR_c_633_n 0.0307558f $X=4.145 $Y=1.54 $X2=0
+ $Y2=0
cc_290 N_A_113_47#_c_311_n N_VPWR_c_633_n 0.0121586f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A_113_47#_c_314_n N_VPWR_c_634_n 0.00300743f $X=5.235 $Y=1.41 $X2=0
+ $Y2=0
cc_292 N_A_113_47#_c_315_n N_VPWR_c_634_n 0.00300743f $X=5.705 $Y=1.41 $X2=0
+ $Y2=0
cc_293 N_A_113_47#_c_316_n N_VPWR_c_635_n 0.00479105f $X=6.175 $Y=1.41 $X2=0
+ $Y2=0
cc_294 N_A_113_47#_c_313_n N_VPWR_c_638_n 0.00702461f $X=4.765 $Y=1.41 $X2=0
+ $Y2=0
cc_295 N_A_113_47#_c_314_n N_VPWR_c_638_n 0.00702461f $X=5.235 $Y=1.41 $X2=0
+ $Y2=0
cc_296 N_A_113_47#_c_315_n N_VPWR_c_640_n 0.00702461f $X=5.705 $Y=1.41 $X2=0
+ $Y2=0
cc_297 N_A_113_47#_c_316_n N_VPWR_c_640_n 0.00702461f $X=6.175 $Y=1.41 $X2=0
+ $Y2=0
cc_298 N_A_113_47#_c_395_p N_VPWR_c_646_n 0.0149311f $X=3.57 $Y=2.3 $X2=0 $Y2=0
cc_299 N_A_113_47#_M1002_d N_VPWR_c_624_n 0.00370124f $X=0.605 $Y=1.485 $X2=0
+ $Y2=0
cc_300 N_A_113_47#_M1018_d N_VPWR_c_624_n 0.00370124f $X=1.545 $Y=1.485 $X2=0
+ $Y2=0
cc_301 N_A_113_47#_M1001_d N_VPWR_c_624_n 0.00370124f $X=2.485 $Y=1.485 $X2=0
+ $Y2=0
cc_302 N_A_113_47#_M1035_d N_VPWR_c_624_n 0.00370124f $X=3.425 $Y=1.485 $X2=0
+ $Y2=0
cc_303 N_A_113_47#_c_313_n N_VPWR_c_624_n 0.0136915f $X=4.765 $Y=1.41 $X2=0
+ $Y2=0
cc_304 N_A_113_47#_c_314_n N_VPWR_c_624_n 0.0124092f $X=5.235 $Y=1.41 $X2=0
+ $Y2=0
cc_305 N_A_113_47#_c_315_n N_VPWR_c_624_n 0.0124092f $X=5.705 $Y=1.41 $X2=0
+ $Y2=0
cc_306 N_A_113_47#_c_316_n N_VPWR_c_624_n 0.0136915f $X=6.175 $Y=1.41 $X2=0
+ $Y2=0
cc_307 N_A_113_47#_c_379_p N_VPWR_c_624_n 0.00955092f $X=0.75 $Y=2.3 $X2=0 $Y2=0
cc_308 N_A_113_47#_c_381_p N_VPWR_c_624_n 0.00955092f $X=1.69 $Y=2.3 $X2=0 $Y2=0
cc_309 N_A_113_47#_c_383_p N_VPWR_c_624_n 0.00955092f $X=2.63 $Y=2.3 $X2=0 $Y2=0
cc_310 N_A_113_47#_c_395_p N_VPWR_c_624_n 0.00955092f $X=3.57 $Y=2.3 $X2=0 $Y2=0
cc_311 N_A_113_47#_c_302_n N_Y_c_774_n 3.30826e-19 $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_113_47#_c_303_n N_Y_c_774_n 0.0114127f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A_113_47#_c_304_n N_Y_c_774_n 0.0114769f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A_113_47#_c_305_n N_Y_c_774_n 0.0138468f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A_113_47#_c_311_n N_Y_c_774_n 0.106439f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A_113_47#_c_312_n N_Y_c_774_n 0.0117089f $X=6.175 $Y=1.202 $X2=0 $Y2=0
cc_317 N_A_113_47#_c_313_n N_Y_c_776_n 4.79893e-19 $X=4.765 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_113_47#_c_323_n N_Y_c_776_n 0.00376966f $X=4.145 $Y=1.54 $X2=0 $Y2=0
cc_319 N_A_113_47#_c_311_n N_Y_c_776_n 0.0204509f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_113_47#_c_312_n N_Y_c_776_n 0.00656533f $X=6.175 $Y=1.202 $X2=0 $Y2=0
cc_321 N_A_113_47#_c_314_n N_Y_c_777_n 0.0155666f $X=5.235 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A_113_47#_c_315_n N_Y_c_777_n 0.0156273f $X=5.705 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A_113_47#_c_311_n N_Y_c_777_n 0.0486996f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A_113_47#_c_312_n N_Y_c_777_n 0.00864922f $X=6.175 $Y=1.202 $X2=0 $Y2=0
cc_325 N_A_113_47#_c_316_n N_Y_c_778_n 0.0176272f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A_113_47#_c_311_n N_Y_c_778_n 0.0167226f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A_113_47#_c_312_n N_Y_c_778_n 0.001713f $X=6.175 $Y=1.202 $X2=0 $Y2=0
cc_328 N_A_113_47#_c_311_n N_Y_c_781_n 0.0204509f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_113_47#_c_312_n N_Y_c_781_n 0.00635938f $X=6.175 $Y=1.202 $X2=0 $Y2=0
cc_330 N_A_113_47#_c_316_n Y 0.00159364f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_331 N_A_113_47#_c_305_n Y 0.0068951f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_113_47#_c_311_n Y 0.0174544f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A_113_47#_c_312_n Y 0.00648765f $X=6.175 $Y=1.202 $X2=0 $Y2=0
cc_334 N_A_113_47#_c_307_n N_A_27_47#_M1003_d 0.00261124f $X=0.255 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_335 N_A_113_47#_c_308_n N_A_27_47#_M1003_d 0.00106131f $X=1.69 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_336 N_A_113_47#_c_308_n N_A_27_47#_M1021_d 0.00214342f $X=1.69 $Y=0.73 $X2=0
+ $Y2=0
cc_337 N_A_113_47#_M1003_s N_A_27_47#_c_927_n 0.00400389f $X=0.565 $Y=0.235
+ $X2=0 $Y2=0
cc_338 N_A_113_47#_M1022_s N_A_27_47#_c_927_n 0.00507817f $X=1.505 $Y=0.235
+ $X2=0 $Y2=0
cc_339 N_A_113_47#_c_307_n N_A_27_47#_c_927_n 0.0122591f $X=0.255 $Y=0.775 $X2=0
+ $Y2=0
cc_340 N_A_113_47#_c_308_n N_A_27_47#_c_927_n 0.0863013f $X=1.69 $Y=0.73 $X2=0
+ $Y2=0
cc_341 N_A_113_47#_c_308_n N_A_27_47#_c_928_n 0.00140356f $X=1.69 $Y=0.73 $X2=0
+ $Y2=0
cc_342 N_A_113_47#_c_321_n N_A_27_47#_c_928_n 0.00817864f $X=2.505 $Y=1.54 $X2=0
+ $Y2=0
cc_343 N_A_113_47#_c_302_n N_A_27_47#_c_930_n 0.00152401f $X=4.77 $Y=0.995 $X2=0
+ $Y2=0
cc_344 N_A_113_47#_c_323_n N_A_27_47#_c_930_n 0.00890545f $X=4.145 $Y=1.54 $X2=0
+ $Y2=0
cc_345 N_A_113_47#_c_310_n N_A_27_47#_c_930_n 0.00551491f $X=4.315 $Y=1.18 $X2=0
+ $Y2=0
cc_346 N_A_113_47#_c_302_n N_A_27_47#_c_931_n 7.67377e-19 $X=4.77 $Y=0.995 $X2=0
+ $Y2=0
cc_347 N_A_113_47#_c_307_n N_VGND_c_1010_n 2.98364e-19 $X=0.255 $Y=0.775 $X2=0
+ $Y2=0
cc_348 N_A_113_47#_c_302_n N_VGND_c_1014_n 0.00357877f $X=4.77 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A_113_47#_c_303_n N_VGND_c_1014_n 0.00357877f $X=5.24 $Y=0.995 $X2=0
+ $Y2=0
cc_350 N_A_113_47#_c_304_n N_VGND_c_1014_n 0.00357877f $X=5.71 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_113_47#_c_305_n N_VGND_c_1014_n 0.00357877f $X=6.23 $Y=0.995 $X2=0
+ $Y2=0
cc_352 N_A_113_47#_M1003_s N_VGND_c_1023_n 0.00256987f $X=0.565 $Y=0.235 $X2=0
+ $Y2=0
cc_353 N_A_113_47#_M1022_s N_VGND_c_1023_n 0.00297142f $X=1.505 $Y=0.235 $X2=0
+ $Y2=0
cc_354 N_A_113_47#_c_302_n N_VGND_c_1023_n 0.00677297f $X=4.77 $Y=0.995 $X2=0
+ $Y2=0
cc_355 N_A_113_47#_c_303_n N_VGND_c_1023_n 0.00548399f $X=5.24 $Y=0.995 $X2=0
+ $Y2=0
cc_356 N_A_113_47#_c_304_n N_VGND_c_1023_n 0.00560377f $X=5.71 $Y=0.995 $X2=0
+ $Y2=0
cc_357 N_A_113_47#_c_305_n N_VGND_c_1023_n 0.00680287f $X=6.23 $Y=0.995 $X2=0
+ $Y2=0
cc_358 N_A_113_47#_c_307_n N_VGND_c_1023_n 8.363e-19 $X=0.255 $Y=0.775 $X2=0
+ $Y2=0
cc_359 N_A_113_47#_c_311_n N_A_887_47#_c_1164_n 0.0116182f $X=6.03 $Y=1.16 $X2=0
+ $Y2=0
cc_360 N_A_113_47#_c_302_n N_A_887_47#_c_1165_n 0.0138413f $X=4.77 $Y=0.995
+ $X2=0 $Y2=0
cc_361 N_A_113_47#_c_303_n N_A_887_47#_c_1165_n 0.00923997f $X=5.24 $Y=0.995
+ $X2=0 $Y2=0
cc_362 N_A_113_47#_c_304_n N_A_887_47#_c_1165_n 0.00964761f $X=5.71 $Y=0.995
+ $X2=0 $Y2=0
cc_363 N_A_113_47#_c_305_n N_A_887_47#_c_1165_n 0.00964761f $X=6.23 $Y=0.995
+ $X2=0 $Y2=0
cc_364 N_A_113_47#_c_311_n N_A_887_47#_c_1165_n 0.00464238f $X=6.03 $Y=1.16
+ $X2=0 $Y2=0
cc_365 N_A_113_47#_c_305_n N_A_887_47#_c_1170_n 0.00260271f $X=6.23 $Y=0.995
+ $X2=0 $Y2=0
cc_366 N_A_113_47#_c_305_n N_A_887_47#_c_1156_n 5.08187e-19 $X=6.23 $Y=0.995
+ $X2=0 $Y2=0
cc_367 N_B2_c_467_n N_B1_c_549_n 0.0175833f $X=8.6 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_368 N_B2_c_473_n N_B1_c_555_n 0.00971598f $X=8.575 $Y=1.41 $X2=0 $Y2=0
cc_369 N_B2_c_468_n N_B1_c_553_n 0.0185441f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_370 N_B2_c_469_n N_B1_c_553_n 8.21108e-19 $X=8.575 $Y=1.202 $X2=0 $Y2=0
cc_371 N_B2_c_468_n N_B1_c_554_n 2.16854e-19 $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_372 N_B2_c_469_n N_B1_c_554_n 0.0175833f $X=8.575 $Y=1.202 $X2=0 $Y2=0
cc_373 N_B2_c_470_n N_VPWR_c_635_n 0.00213375f $X=7.165 $Y=1.41 $X2=0 $Y2=0
cc_374 N_B2_c_470_n N_VPWR_c_642_n 0.00429453f $X=7.165 $Y=1.41 $X2=0 $Y2=0
cc_375 N_B2_c_471_n N_VPWR_c_642_n 0.00429453f $X=7.635 $Y=1.41 $X2=0 $Y2=0
cc_376 N_B2_c_472_n N_VPWR_c_642_n 0.00429453f $X=8.105 $Y=1.41 $X2=0 $Y2=0
cc_377 N_B2_c_473_n N_VPWR_c_642_n 0.00429453f $X=8.575 $Y=1.41 $X2=0 $Y2=0
cc_378 N_B2_c_470_n N_VPWR_c_624_n 0.00734734f $X=7.165 $Y=1.41 $X2=0 $Y2=0
cc_379 N_B2_c_471_n N_VPWR_c_624_n 0.00606499f $X=7.635 $Y=1.41 $X2=0 $Y2=0
cc_380 N_B2_c_472_n N_VPWR_c_624_n 0.00606499f $X=8.105 $Y=1.41 $X2=0 $Y2=0
cc_381 N_B2_c_473_n N_VPWR_c_624_n 0.00609021f $X=8.575 $Y=1.41 $X2=0 $Y2=0
cc_382 N_B2_c_464_n N_Y_c_774_n 0.00166811f $X=7.14 $Y=0.995 $X2=0 $Y2=0
cc_383 N_B2_c_470_n N_Y_c_779_n 0.0148794f $X=7.165 $Y=1.41 $X2=0 $Y2=0
cc_384 N_B2_c_468_n N_Y_c_779_n 0.0145434f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_385 N_B2_c_469_n N_Y_c_779_n 8.84531e-19 $X=8.575 $Y=1.202 $X2=0 $Y2=0
cc_386 N_B2_c_471_n N_Y_c_780_n 0.0128795f $X=7.635 $Y=1.41 $X2=0 $Y2=0
cc_387 N_B2_c_472_n N_Y_c_780_n 0.0128188f $X=8.105 $Y=1.41 $X2=0 $Y2=0
cc_388 N_B2_c_468_n N_Y_c_780_n 0.0486996f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_389 N_B2_c_469_n N_Y_c_780_n 0.00864922f $X=8.575 $Y=1.202 $X2=0 $Y2=0
cc_390 N_B2_c_468_n N_Y_c_782_n 0.0204252f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_391 N_B2_c_469_n N_Y_c_782_n 0.00655199f $X=8.575 $Y=1.202 $X2=0 $Y2=0
cc_392 N_B2_c_473_n N_Y_c_783_n 2.98195e-19 $X=8.575 $Y=1.41 $X2=0 $Y2=0
cc_393 N_B2_c_468_n N_Y_c_783_n 0.0204252f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_394 N_B2_c_469_n N_Y_c_783_n 0.00634604f $X=8.575 $Y=1.202 $X2=0 $Y2=0
cc_395 N_B2_c_464_n Y 0.00626083f $X=7.14 $Y=0.995 $X2=0 $Y2=0
cc_396 N_B2_c_470_n Y 0.00149476f $X=7.165 $Y=1.41 $X2=0 $Y2=0
cc_397 N_B2_c_468_n Y 0.0126857f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_398 N_B2_c_469_n Y 0.00602197f $X=8.575 $Y=1.202 $X2=0 $Y2=0
cc_399 N_B2_c_470_n N_A_1361_297#_c_871_n 0.01161f $X=7.165 $Y=1.41 $X2=0 $Y2=0
cc_400 N_B2_c_471_n N_A_1361_297#_c_871_n 0.01161f $X=7.635 $Y=1.41 $X2=0 $Y2=0
cc_401 N_B2_c_472_n N_A_1361_297#_c_873_n 0.01161f $X=8.105 $Y=1.41 $X2=0 $Y2=0
cc_402 N_B2_c_473_n N_A_1361_297#_c_873_n 0.0143578f $X=8.575 $Y=1.41 $X2=0
+ $Y2=0
cc_403 N_B2_c_473_n N_A_1361_297#_c_865_n 2.98195e-19 $X=8.575 $Y=1.41 $X2=0
+ $Y2=0
cc_404 N_B2_c_464_n N_VGND_c_1006_n 0.00358858f $X=7.14 $Y=0.995 $X2=0 $Y2=0
cc_405 N_B2_c_465_n N_VGND_c_1006_n 0.00276126f $X=7.61 $Y=0.995 $X2=0 $Y2=0
cc_406 N_B2_c_466_n N_VGND_c_1007_n 0.00385467f $X=8.08 $Y=0.995 $X2=0 $Y2=0
cc_407 N_B2_c_467_n N_VGND_c_1007_n 0.00365402f $X=8.6 $Y=0.995 $X2=0 $Y2=0
cc_408 N_B2_c_464_n N_VGND_c_1014_n 0.00395719f $X=7.14 $Y=0.995 $X2=0 $Y2=0
cc_409 N_B2_c_465_n N_VGND_c_1016_n 0.00424416f $X=7.61 $Y=0.995 $X2=0 $Y2=0
cc_410 N_B2_c_466_n N_VGND_c_1016_n 0.00423334f $X=8.08 $Y=0.995 $X2=0 $Y2=0
cc_411 N_B2_c_467_n N_VGND_c_1018_n 0.00396605f $X=8.6 $Y=0.995 $X2=0 $Y2=0
cc_412 N_B2_c_464_n N_VGND_c_1023_n 0.00703448f $X=7.14 $Y=0.995 $X2=0 $Y2=0
cc_413 N_B2_c_465_n N_VGND_c_1023_n 0.00599001f $X=7.61 $Y=0.995 $X2=0 $Y2=0
cc_414 N_B2_c_466_n N_VGND_c_1023_n 0.00620835f $X=8.08 $Y=0.995 $X2=0 $Y2=0
cc_415 N_B2_c_467_n N_VGND_c_1023_n 0.00583042f $X=8.6 $Y=0.995 $X2=0 $Y2=0
cc_416 N_B2_c_464_n N_A_887_47#_c_1165_n 0.00373464f $X=7.14 $Y=0.995 $X2=0
+ $Y2=0
cc_417 N_B2_c_464_n N_A_887_47#_c_1170_n 0.00724188f $X=7.14 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_B2_c_465_n N_A_887_47#_c_1170_n 5.42894e-19 $X=7.61 $Y=0.995 $X2=0
+ $Y2=0
cc_419 N_B2_c_464_n N_A_887_47#_c_1155_n 0.0060427f $X=7.14 $Y=0.995 $X2=0 $Y2=0
cc_420 N_B2_c_465_n N_A_887_47#_c_1155_n 0.00874287f $X=7.61 $Y=0.995 $X2=0
+ $Y2=0
cc_421 N_B2_c_468_n N_A_887_47#_c_1155_n 0.0362711f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_422 N_B2_c_469_n N_A_887_47#_c_1155_n 0.00345061f $X=8.575 $Y=1.202 $X2=0
+ $Y2=0
cc_423 N_B2_c_464_n N_A_887_47#_c_1156_n 0.00515933f $X=7.14 $Y=0.995 $X2=0
+ $Y2=0
cc_424 N_B2_c_468_n N_A_887_47#_c_1156_n 0.00616095f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_425 N_B2_c_464_n N_A_887_47#_c_1181_n 5.15068e-19 $X=7.14 $Y=0.995 $X2=0
+ $Y2=0
cc_426 N_B2_c_465_n N_A_887_47#_c_1181_n 0.0063752f $X=7.61 $Y=0.995 $X2=0 $Y2=0
cc_427 N_B2_c_466_n N_A_887_47#_c_1181_n 0.00693563f $X=8.08 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_B2_c_467_n N_A_887_47#_c_1181_n 5.34196e-19 $X=8.6 $Y=0.995 $X2=0 $Y2=0
cc_429 N_B2_c_466_n N_A_887_47#_c_1157_n 0.00929182f $X=8.08 $Y=0.995 $X2=0
+ $Y2=0
cc_430 N_B2_c_467_n N_A_887_47#_c_1157_n 0.00650032f $X=8.6 $Y=0.995 $X2=0 $Y2=0
cc_431 N_B2_c_468_n N_A_887_47#_c_1157_n 0.0400808f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_432 N_B2_c_469_n N_A_887_47#_c_1157_n 0.00468948f $X=8.575 $Y=1.202 $X2=0
+ $Y2=0
cc_433 N_B2_c_466_n N_A_887_47#_c_1189_n 5.69266e-19 $X=8.08 $Y=0.995 $X2=0
+ $Y2=0
cc_434 N_B2_c_467_n N_A_887_47#_c_1189_n 0.00857123f $X=8.6 $Y=0.995 $X2=0 $Y2=0
cc_435 N_B2_c_465_n N_A_887_47#_c_1161_n 0.00131596f $X=7.61 $Y=0.995 $X2=0
+ $Y2=0
cc_436 N_B2_c_466_n N_A_887_47#_c_1161_n 0.00116636f $X=8.08 $Y=0.995 $X2=0
+ $Y2=0
cc_437 N_B2_c_468_n N_A_887_47#_c_1161_n 0.0307014f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_438 N_B2_c_469_n N_A_887_47#_c_1161_n 0.00358305f $X=8.575 $Y=1.202 $X2=0
+ $Y2=0
cc_439 N_B2_c_467_n N_A_887_47#_c_1162_n 0.00269873f $X=8.6 $Y=0.995 $X2=0 $Y2=0
cc_440 N_B2_c_468_n N_A_887_47#_c_1162_n 0.00616124f $X=8.4 $Y=1.16 $X2=0 $Y2=0
cc_441 N_B1_c_555_n N_VPWR_c_636_n 0.00300743f $X=9.045 $Y=1.41 $X2=0 $Y2=0
cc_442 N_B1_c_556_n N_VPWR_c_636_n 0.00300743f $X=9.515 $Y=1.41 $X2=0 $Y2=0
cc_443 N_B1_c_557_n N_VPWR_c_637_n 0.00300743f $X=9.985 $Y=1.41 $X2=0 $Y2=0
cc_444 N_B1_c_558_n N_VPWR_c_637_n 0.00300743f $X=10.455 $Y=1.41 $X2=0 $Y2=0
cc_445 N_B1_c_555_n N_VPWR_c_642_n 0.00702461f $X=9.045 $Y=1.41 $X2=0 $Y2=0
cc_446 N_B1_c_556_n N_VPWR_c_644_n 0.00702461f $X=9.515 $Y=1.41 $X2=0 $Y2=0
cc_447 N_B1_c_557_n N_VPWR_c_644_n 0.00702461f $X=9.985 $Y=1.41 $X2=0 $Y2=0
cc_448 N_B1_c_558_n N_VPWR_c_647_n 0.00702461f $X=10.455 $Y=1.41 $X2=0 $Y2=0
cc_449 N_B1_c_555_n N_VPWR_c_624_n 0.0124344f $X=9.045 $Y=1.41 $X2=0 $Y2=0
cc_450 N_B1_c_556_n N_VPWR_c_624_n 0.0124092f $X=9.515 $Y=1.41 $X2=0 $Y2=0
cc_451 N_B1_c_557_n N_VPWR_c_624_n 0.0124092f $X=9.985 $Y=1.41 $X2=0 $Y2=0
cc_452 N_B1_c_558_n N_VPWR_c_624_n 0.0133942f $X=10.455 $Y=1.41 $X2=0 $Y2=0
cc_453 N_B1_c_553_n N_A_1361_297#_c_865_n 0.00771248f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_454 N_B1_c_555_n N_A_1361_297#_c_866_n 0.0155666f $X=9.045 $Y=1.41 $X2=0
+ $Y2=0
cc_455 N_B1_c_556_n N_A_1361_297#_c_866_n 0.0156273f $X=9.515 $Y=1.41 $X2=0
+ $Y2=0
cc_456 N_B1_c_553_n N_A_1361_297#_c_866_n 0.0487385f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_457 N_B1_c_554_n N_A_1361_297#_c_866_n 0.00837544f $X=10.455 $Y=1.202 $X2=0
+ $Y2=0
cc_458 N_B1_c_557_n N_A_1361_297#_c_867_n 0.0156273f $X=9.985 $Y=1.41 $X2=0
+ $Y2=0
cc_459 N_B1_c_558_n N_A_1361_297#_c_867_n 0.0158589f $X=10.455 $Y=1.41 $X2=0
+ $Y2=0
cc_460 N_B1_c_553_n N_A_1361_297#_c_867_n 0.0487385f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_461 N_B1_c_554_n N_A_1361_297#_c_867_n 0.00816971f $X=10.455 $Y=1.202 $X2=0
+ $Y2=0
cc_462 N_B1_c_553_n N_A_1361_297#_c_868_n 0.0265652f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_463 N_B1_c_553_n N_A_1361_297#_c_870_n 0.0204509f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_464 N_B1_c_554_n N_A_1361_297#_c_870_n 0.00656533f $X=10.455 $Y=1.202 $X2=0
+ $Y2=0
cc_465 N_B1_c_549_n N_VGND_c_1008_n 0.00379224f $X=9.02 $Y=0.995 $X2=0 $Y2=0
cc_466 N_B1_c_550_n N_VGND_c_1008_n 0.00276126f $X=9.49 $Y=0.995 $X2=0 $Y2=0
cc_467 N_B1_c_551_n N_VGND_c_1009_n 0.00385467f $X=9.96 $Y=0.995 $X2=0 $Y2=0
cc_468 N_B1_c_552_n N_VGND_c_1009_n 0.00365402f $X=10.48 $Y=0.995 $X2=0 $Y2=0
cc_469 N_B1_c_549_n N_VGND_c_1018_n 0.00423334f $X=9.02 $Y=0.995 $X2=0 $Y2=0
cc_470 N_B1_c_550_n N_VGND_c_1020_n 0.00423334f $X=9.49 $Y=0.995 $X2=0 $Y2=0
cc_471 N_B1_c_551_n N_VGND_c_1020_n 0.00423334f $X=9.96 $Y=0.995 $X2=0 $Y2=0
cc_472 N_B1_c_552_n N_VGND_c_1022_n 0.00396605f $X=10.48 $Y=0.995 $X2=0 $Y2=0
cc_473 N_B1_c_549_n N_VGND_c_1023_n 0.00599324f $X=9.02 $Y=0.995 $X2=0 $Y2=0
cc_474 N_B1_c_550_n N_VGND_c_1023_n 0.00597024f $X=9.49 $Y=0.995 $X2=0 $Y2=0
cc_475 N_B1_c_551_n N_VGND_c_1023_n 0.00620835f $X=9.96 $Y=0.995 $X2=0 $Y2=0
cc_476 N_B1_c_552_n N_VGND_c_1023_n 0.00683325f $X=10.48 $Y=0.995 $X2=0 $Y2=0
cc_477 N_B1_c_549_n N_A_887_47#_c_1189_n 0.00686626f $X=9.02 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_B1_c_550_n N_A_887_47#_c_1189_n 5.45498e-19 $X=9.49 $Y=0.995 $X2=0
+ $Y2=0
cc_479 N_B1_c_549_n N_A_887_47#_c_1158_n 0.00901745f $X=9.02 $Y=0.995 $X2=0
+ $Y2=0
cc_480 N_B1_c_550_n N_A_887_47#_c_1158_n 0.00901745f $X=9.49 $Y=0.995 $X2=0
+ $Y2=0
cc_481 N_B1_c_553_n N_A_887_47#_c_1158_n 0.0398926f $X=10.25 $Y=1.16 $X2=0 $Y2=0
cc_482 N_B1_c_554_n N_A_887_47#_c_1158_n 0.00345541f $X=10.455 $Y=1.202 $X2=0
+ $Y2=0
cc_483 N_B1_c_549_n N_A_887_47#_c_1203_n 5.24597e-19 $X=9.02 $Y=0.995 $X2=0
+ $Y2=0
cc_484 N_B1_c_550_n N_A_887_47#_c_1203_n 0.00651696f $X=9.49 $Y=0.995 $X2=0
+ $Y2=0
cc_485 N_B1_c_551_n N_A_887_47#_c_1203_n 0.00693563f $X=9.96 $Y=0.995 $X2=0
+ $Y2=0
cc_486 N_B1_c_552_n N_A_887_47#_c_1203_n 5.34196e-19 $X=10.48 $Y=0.995 $X2=0
+ $Y2=0
cc_487 N_B1_c_551_n N_A_887_47#_c_1159_n 0.00929182f $X=9.96 $Y=0.995 $X2=0
+ $Y2=0
cc_488 N_B1_c_552_n N_A_887_47#_c_1159_n 0.00936658f $X=10.48 $Y=0.995 $X2=0
+ $Y2=0
cc_489 N_B1_c_553_n N_A_887_47#_c_1159_n 0.071856f $X=10.25 $Y=1.16 $X2=0 $Y2=0
cc_490 N_B1_c_554_n N_A_887_47#_c_1159_n 0.00468948f $X=10.455 $Y=1.202 $X2=0
+ $Y2=0
cc_491 N_B1_c_551_n N_A_887_47#_c_1160_n 5.69266e-19 $X=9.96 $Y=0.995 $X2=0
+ $Y2=0
cc_492 N_B1_c_552_n N_A_887_47#_c_1160_n 0.00857123f $X=10.48 $Y=0.995 $X2=0
+ $Y2=0
cc_493 N_B1_c_549_n N_A_887_47#_c_1162_n 0.00112787f $X=9.02 $Y=0.995 $X2=0
+ $Y2=0
cc_494 N_B1_c_553_n N_A_887_47#_c_1162_n 0.0108485f $X=10.25 $Y=1.16 $X2=0 $Y2=0
cc_495 N_B1_c_550_n N_A_887_47#_c_1163_n 0.00116636f $X=9.49 $Y=0.995 $X2=0
+ $Y2=0
cc_496 N_B1_c_551_n N_A_887_47#_c_1163_n 0.00116636f $X=9.96 $Y=0.995 $X2=0
+ $Y2=0
cc_497 N_B1_c_553_n N_A_887_47#_c_1163_n 0.0307014f $X=10.25 $Y=1.16 $X2=0 $Y2=0
cc_498 N_B1_c_554_n N_A_887_47#_c_1163_n 0.00358305f $X=10.455 $Y=1.202 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_624_n N_Y_M1004_s 0.00370124f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_500 N_VPWR_c_624_n N_Y_M1019_s 0.00370124f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_501 N_VPWR_c_624_n N_Y_M1011_d 0.00232895f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_502 N_VPWR_c_624_n N_Y_M1030_d 0.00232895f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_503 N_VPWR_c_638_n N_Y_c_829_n 0.0149311f $X=5.345 $Y=2.72 $X2=0 $Y2=0
cc_504 N_VPWR_c_624_n N_Y_c_829_n 0.00955092f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_505 N_VPWR_M1007_d N_Y_c_777_n 0.00187091f $X=5.325 $Y=1.485 $X2=0 $Y2=0
cc_506 N_VPWR_c_634_n N_Y_c_777_n 0.0143191f $X=5.47 $Y=1.96 $X2=0 $Y2=0
cc_507 N_VPWR_c_640_n N_Y_c_833_n 0.0149311f $X=6.285 $Y=2.72 $X2=0 $Y2=0
cc_508 N_VPWR_c_624_n N_Y_c_833_n 0.00955092f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_509 N_VPWR_M1036_d N_Y_c_778_n 0.00183891f $X=6.265 $Y=1.485 $X2=0 $Y2=0
cc_510 N_VPWR_c_635_n N_Y_c_778_n 0.0124114f $X=6.41 $Y=1.96 $X2=0 $Y2=0
cc_511 N_VPWR_M1036_d Y 0.00111785f $X=6.265 $Y=1.485 $X2=0 $Y2=0
cc_512 N_VPWR_c_635_n Y 0.00531954f $X=6.41 $Y=1.96 $X2=0 $Y2=0
cc_513 N_VPWR_c_624_n N_A_1361_297#_M1011_s 0.00217519f $X=10.81 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_514 N_VPWR_c_624_n N_A_1361_297#_M1024_s 0.00231264f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_624_n N_A_1361_297#_M1032_s 0.00297222f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_624_n N_A_1361_297#_M1014_s 0.00370124f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_624_n N_A_1361_297#_M1025_s 0.00303344f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_635_n N_A_1361_297#_c_863_n 0.0308496f $X=6.41 $Y=1.96 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_642_n N_A_1361_297#_c_871_n 0.0386815f $X=9.155 $Y=2.72 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_624_n N_A_1361_297#_c_871_n 0.0239144f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_635_n N_A_1361_297#_c_864_n 0.0113145f $X=6.41 $Y=1.96 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_642_n N_A_1361_297#_c_864_n 0.0183872f $X=9.155 $Y=2.72 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_624_n N_A_1361_297#_c_864_n 0.0107739f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_642_n N_A_1361_297#_c_873_n 0.0386815f $X=9.155 $Y=2.72 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_624_n N_A_1361_297#_c_873_n 0.0239144f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_642_n N_A_1361_297#_c_901_n 0.015002f $X=9.155 $Y=2.72 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_624_n N_A_1361_297#_c_901_n 0.00962794f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_528 N_VPWR_M1005_d N_A_1361_297#_c_866_n 0.00187091f $X=9.135 $Y=1.485 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_636_n N_A_1361_297#_c_866_n 0.0143191f $X=9.28 $Y=1.96 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_644_n N_A_1361_297#_c_905_n 0.0149311f $X=10.095 $Y=2.72 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_624_n N_A_1361_297#_c_905_n 0.00955092f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_532 N_VPWR_M1020_d N_A_1361_297#_c_867_n 0.00187091f $X=10.075 $Y=1.485 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_637_n N_A_1361_297#_c_867_n 0.0143191f $X=10.22 $Y=1.96 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_647_n N_A_1361_297#_c_869_n 0.0204581f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_624_n N_A_1361_297#_c_869_n 0.0118616f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_642_n N_A_1361_297#_c_911_n 0.0149886f $X=9.155 $Y=2.72 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_624_n N_A_1361_297#_c_911_n 0.00962421f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_538 N_Y_c_779_n N_A_1361_297#_M1011_s 0.00293834f $X=7.275 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_539 N_Y_c_780_n N_A_1361_297#_M1024_s 0.00187091f $X=8.215 $Y=1.54 $X2=0
+ $Y2=0
cc_540 N_Y_c_779_n N_A_1361_297#_c_863_n 0.0172719f $X=7.275 $Y=1.54 $X2=0 $Y2=0
cc_541 Y N_A_1361_297#_c_863_n 0.00262061f $X=6.585 $Y=1.445 $X2=0 $Y2=0
cc_542 N_Y_M1011_d N_A_1361_297#_c_871_n 0.00352392f $X=7.255 $Y=1.485 $X2=0
+ $Y2=0
cc_543 N_Y_c_779_n N_A_1361_297#_c_871_n 0.00385532f $X=7.275 $Y=1.54 $X2=0
+ $Y2=0
cc_544 N_Y_c_780_n N_A_1361_297#_c_871_n 0.00385532f $X=8.215 $Y=1.54 $X2=0
+ $Y2=0
cc_545 N_Y_c_782_n N_A_1361_297#_c_871_n 0.013395f $X=7.4 $Y=1.62 $X2=0 $Y2=0
cc_546 N_Y_c_780_n N_A_1361_297#_c_921_n 0.0143018f $X=8.215 $Y=1.54 $X2=0 $Y2=0
cc_547 N_Y_M1030_d N_A_1361_297#_c_873_n 0.00352392f $X=8.195 $Y=1.485 $X2=0
+ $Y2=0
cc_548 N_Y_c_780_n N_A_1361_297#_c_873_n 0.00385532f $X=8.215 $Y=1.54 $X2=0
+ $Y2=0
cc_549 N_Y_c_783_n N_A_1361_297#_c_873_n 0.013395f $X=8.34 $Y=1.62 $X2=0 $Y2=0
cc_550 N_Y_c_783_n N_A_1361_297#_c_865_n 0.00226124f $X=8.34 $Y=1.62 $X2=0 $Y2=0
cc_551 N_Y_c_774_n N_A_27_47#_c_930_n 0.00156115f $X=6.475 $Y=0.775 $X2=0 $Y2=0
cc_552 N_Y_M1006_d N_VGND_c_1023_n 0.00256987f $X=4.845 $Y=0.235 $X2=0 $Y2=0
cc_553 N_Y_M1028_d N_VGND_c_1023_n 0.00297142f $X=5.785 $Y=0.235 $X2=0 $Y2=0
cc_554 N_Y_c_774_n N_A_887_47#_M1008_s 0.00214342f $X=6.475 $Y=0.775 $X2=0 $Y2=0
cc_555 N_Y_c_774_n N_A_887_47#_M1033_s 0.0111033f $X=6.475 $Y=0.775 $X2=0 $Y2=0
cc_556 N_Y_M1006_d N_A_887_47#_c_1165_n 0.00400389f $X=4.845 $Y=0.235 $X2=0
+ $Y2=0
cc_557 N_Y_M1028_d N_A_887_47#_c_1165_n 0.00507817f $X=5.785 $Y=0.235 $X2=0
+ $Y2=0
cc_558 N_Y_c_774_n N_A_887_47#_c_1165_n 0.112904f $X=6.475 $Y=0.775 $X2=0 $Y2=0
cc_559 N_Y_c_774_n N_A_887_47#_c_1170_n 0.00728572f $X=6.475 $Y=0.775 $X2=0
+ $Y2=0
cc_560 N_Y_c_774_n N_A_887_47#_c_1156_n 0.0153979f $X=6.475 $Y=0.775 $X2=0 $Y2=0
cc_561 N_Y_c_779_n N_A_887_47#_c_1156_n 0.00334581f $X=7.275 $Y=1.54 $X2=0 $Y2=0
cc_562 N_A_1361_297#_c_865_n N_A_887_47#_c_1162_n 0.00658191f $X=8.81 $Y=1.625
+ $X2=0 $Y2=0
cc_563 N_A_27_47#_c_929_n N_VGND_M1015_d 0.00251047f $X=2.885 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_564 N_A_27_47#_c_930_n N_VGND_M1031_d 0.00348805f $X=3.825 $Y=0.815 $X2=0
+ $Y2=0
cc_565 N_A_27_47#_c_938_n N_VGND_c_1004_n 0.0141571f $X=2.2 $Y=0.475 $X2=0 $Y2=0
cc_566 N_A_27_47#_c_928_n N_VGND_c_1004_n 0.00471242f $X=2.2 $Y=0.725 $X2=0
+ $Y2=0
cc_567 N_A_27_47#_c_929_n N_VGND_c_1004_n 0.0127273f $X=2.885 $Y=0.815 $X2=0
+ $Y2=0
cc_568 N_A_27_47#_c_946_n N_VGND_c_1005_n 0.0183628f $X=3.1 $Y=0.39 $X2=0 $Y2=0
cc_569 N_A_27_47#_c_930_n N_VGND_c_1005_n 0.0131987f $X=3.825 $Y=0.815 $X2=0
+ $Y2=0
cc_570 N_A_27_47#_c_931_n N_VGND_c_1005_n 0.0223967f $X=4.04 $Y=0.39 $X2=0 $Y2=0
cc_571 N_A_27_47#_c_927_n N_VGND_c_1010_n 0.113039f $X=2.075 $Y=0.365 $X2=0
+ $Y2=0
cc_572 N_A_27_47#_c_938_n N_VGND_c_1010_n 0.0152108f $X=2.2 $Y=0.475 $X2=0 $Y2=0
cc_573 N_A_27_47#_c_929_n N_VGND_c_1010_n 0.00266636f $X=2.885 $Y=0.815 $X2=0
+ $Y2=0
cc_574 N_A_27_47#_c_929_n N_VGND_c_1012_n 0.00198695f $X=2.885 $Y=0.815 $X2=0
+ $Y2=0
cc_575 N_A_27_47#_c_946_n N_VGND_c_1012_n 0.0223596f $X=3.1 $Y=0.39 $X2=0 $Y2=0
cc_576 N_A_27_47#_c_930_n N_VGND_c_1012_n 0.00266636f $X=3.825 $Y=0.815 $X2=0
+ $Y2=0
cc_577 N_A_27_47#_c_930_n N_VGND_c_1014_n 0.00199443f $X=3.825 $Y=0.815 $X2=0
+ $Y2=0
cc_578 N_A_27_47#_c_931_n N_VGND_c_1014_n 0.024373f $X=4.04 $Y=0.39 $X2=0 $Y2=0
cc_579 N_A_27_47#_M1003_d N_VGND_c_1023_n 0.00225742f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_580 N_A_27_47#_M1021_d N_VGND_c_1023_n 0.00255381f $X=1.035 $Y=0.235 $X2=0
+ $Y2=0
cc_581 N_A_27_47#_M1037_d N_VGND_c_1023_n 0.00215206f $X=2.025 $Y=0.235 $X2=0
+ $Y2=0
cc_582 N_A_27_47#_M1017_s N_VGND_c_1023_n 0.0025535f $X=2.915 $Y=0.235 $X2=0
+ $Y2=0
cc_583 N_A_27_47#_M1038_s N_VGND_c_1023_n 0.00209319f $X=3.905 $Y=0.235 $X2=0
+ $Y2=0
cc_584 N_A_27_47#_c_927_n N_VGND_c_1023_n 0.0709513f $X=2.075 $Y=0.365 $X2=0
+ $Y2=0
cc_585 N_A_27_47#_c_938_n N_VGND_c_1023_n 0.00940698f $X=2.2 $Y=0.475 $X2=0
+ $Y2=0
cc_586 N_A_27_47#_c_929_n N_VGND_c_1023_n 0.00972452f $X=2.885 $Y=0.815 $X2=0
+ $Y2=0
cc_587 N_A_27_47#_c_946_n N_VGND_c_1023_n 0.0141302f $X=3.1 $Y=0.39 $X2=0 $Y2=0
cc_588 N_A_27_47#_c_930_n N_VGND_c_1023_n 0.0100158f $X=3.825 $Y=0.815 $X2=0
+ $Y2=0
cc_589 N_A_27_47#_c_931_n N_VGND_c_1023_n 0.0141066f $X=4.04 $Y=0.39 $X2=0 $Y2=0
cc_590 N_A_27_47#_c_930_n N_A_887_47#_c_1164_n 0.00687335f $X=3.825 $Y=0.815
+ $X2=0 $Y2=0
cc_591 N_A_27_47#_c_931_n N_A_887_47#_c_1164_n 0.0147785f $X=4.04 $Y=0.39 $X2=0
+ $Y2=0
cc_592 N_A_27_47#_c_931_n N_A_887_47#_c_1230_n 0.0143874f $X=4.04 $Y=0.39 $X2=0
+ $Y2=0
cc_593 N_VGND_c_1023_n N_A_887_47#_M1006_s 0.00296916f $X=10.81 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_594 N_VGND_c_1023_n N_A_887_47#_M1008_s 0.00255381f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_c_1023_n N_A_887_47#_M1033_s 0.00615454f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_596 N_VGND_c_1023_n N_A_887_47#_M1013_s 0.0025535f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_597 N_VGND_c_1023_n N_A_887_47#_M1034_s 0.00215201f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_c_1023_n N_A_887_47#_M1012_s 0.0025535f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_599 N_VGND_c_1023_n N_A_887_47#_M1027_s 0.00209319f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_600 N_VGND_c_1006_n N_A_887_47#_c_1165_n 0.0172916f $X=7.4 $Y=0.39 $X2=0
+ $Y2=0
cc_601 N_VGND_c_1014_n N_A_887_47#_c_1165_n 0.145636f $X=7.315 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_c_1023_n N_A_887_47#_c_1165_n 0.0904143f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_603 N_VGND_c_1014_n N_A_887_47#_c_1230_n 0.0126217f $X=7.315 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_1023_n N_A_887_47#_c_1230_n 0.00709554f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_605 N_VGND_c_1006_n N_A_887_47#_c_1170_n 0.00558246f $X=7.4 $Y=0.39 $X2=0
+ $Y2=0
cc_606 N_VGND_M1000_d N_A_887_47#_c_1155_n 0.00255557f $X=7.215 $Y=0.235 $X2=0
+ $Y2=0
cc_607 N_VGND_c_1006_n N_A_887_47#_c_1155_n 0.012101f $X=7.4 $Y=0.39 $X2=0 $Y2=0
cc_608 N_VGND_c_1014_n N_A_887_47#_c_1155_n 0.00194552f $X=7.315 $Y=0 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1016_n N_A_887_47#_c_1155_n 0.00193763f $X=8.255 $Y=0 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1023_n N_A_887_47#_c_1155_n 0.00856326f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1007_n N_A_887_47#_c_1181_n 0.0183628f $X=8.34 $Y=0.39 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1016_n N_A_887_47#_c_1181_n 0.0223596f $X=8.255 $Y=0 $X2=0 $Y2=0
cc_613 N_VGND_c_1023_n N_A_887_47#_c_1181_n 0.0141302f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_M1016_d N_A_887_47#_c_1157_n 0.00348805f $X=8.155 $Y=0.235 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1007_n N_A_887_47#_c_1157_n 0.0131987f $X=8.34 $Y=0.39 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1016_n N_A_887_47#_c_1157_n 0.00266636f $X=8.255 $Y=0 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1018_n N_A_887_47#_c_1157_n 0.00199443f $X=9.195 $Y=0 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1023_n N_A_887_47#_c_1157_n 0.0100158f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_c_1007_n N_A_887_47#_c_1189_n 0.0223967f $X=8.34 $Y=0.39 $X2=0
+ $Y2=0
cc_620 N_VGND_c_1008_n N_A_887_47#_c_1189_n 0.0183628f $X=9.28 $Y=0.39 $X2=0
+ $Y2=0
cc_621 N_VGND_c_1018_n N_A_887_47#_c_1189_n 0.0222529f $X=9.195 $Y=0 $X2=0 $Y2=0
cc_622 N_VGND_c_1023_n N_A_887_47#_c_1189_n 0.0139016f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_623 N_VGND_M1009_d N_A_887_47#_c_1158_n 0.00251047f $X=9.095 $Y=0.235 $X2=0
+ $Y2=0
cc_624 N_VGND_c_1008_n N_A_887_47#_c_1158_n 0.0127273f $X=9.28 $Y=0.39 $X2=0
+ $Y2=0
cc_625 N_VGND_c_1018_n N_A_887_47#_c_1158_n 0.00266636f $X=9.195 $Y=0 $X2=0
+ $Y2=0
cc_626 N_VGND_c_1020_n N_A_887_47#_c_1158_n 0.00198695f $X=10.135 $Y=0 $X2=0
+ $Y2=0
cc_627 N_VGND_c_1023_n N_A_887_47#_c_1158_n 0.00972452f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_628 N_VGND_c_1009_n N_A_887_47#_c_1203_n 0.0183628f $X=10.22 $Y=0.39 $X2=0
+ $Y2=0
cc_629 N_VGND_c_1020_n N_A_887_47#_c_1203_n 0.0223596f $X=10.135 $Y=0 $X2=0
+ $Y2=0
cc_630 N_VGND_c_1023_n N_A_887_47#_c_1203_n 0.0141302f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_631 N_VGND_M1026_d N_A_887_47#_c_1159_n 0.00348805f $X=10.035 $Y=0.235 $X2=0
+ $Y2=0
cc_632 N_VGND_c_1009_n N_A_887_47#_c_1159_n 0.0131987f $X=10.22 $Y=0.39 $X2=0
+ $Y2=0
cc_633 N_VGND_c_1020_n N_A_887_47#_c_1159_n 0.00266636f $X=10.135 $Y=0 $X2=0
+ $Y2=0
cc_634 N_VGND_c_1022_n N_A_887_47#_c_1159_n 0.00199443f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_635 N_VGND_c_1023_n N_A_887_47#_c_1159_n 0.0100158f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_636 N_VGND_c_1009_n N_A_887_47#_c_1160_n 0.0223967f $X=10.22 $Y=0.39 $X2=0
+ $Y2=0
cc_637 N_VGND_c_1022_n N_A_887_47#_c_1160_n 0.024373f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_638 N_VGND_c_1023_n N_A_887_47#_c_1160_n 0.0141066f $X=10.81 $Y=0 $X2=0 $Y2=0
