* File: sky130_fd_sc_hdll__a32oi_1.pxi.spice
* Created: Thu Aug 27 18:56:24 2020
* 
x_PM_SKY130_FD_SC_HDLL__A32OI_1%B2 N_B2_c_52_n N_B2_M1002_g N_B2_c_49_n
+ N_B2_M1005_g B2 N_B2_c_51_n PM_SKY130_FD_SC_HDLL__A32OI_1%B2
x_PM_SKY130_FD_SC_HDLL__A32OI_1%B1 N_B1_c_75_n N_B1_M1001_g N_B1_c_76_n
+ N_B1_M1000_g B1 N_B1_c_77_n PM_SKY130_FD_SC_HDLL__A32OI_1%B1
x_PM_SKY130_FD_SC_HDLL__A32OI_1%A1 N_A1_c_107_n N_A1_M1007_g N_A1_c_108_n
+ N_A1_M1009_g A1 PM_SKY130_FD_SC_HDLL__A32OI_1%A1
x_PM_SKY130_FD_SC_HDLL__A32OI_1%A2 N_A2_c_139_n N_A2_M1004_g N_A2_c_140_n
+ N_A2_M1003_g A2 A2 A2 PM_SKY130_FD_SC_HDLL__A32OI_1%A2
x_PM_SKY130_FD_SC_HDLL__A32OI_1%A3 N_A3_M1006_g N_A3_M1008_g N_A3_c_170_n
+ N_A3_c_171_n N_A3_c_172_n A3 N_A3_c_174_n PM_SKY130_FD_SC_HDLL__A32OI_1%A3
x_PM_SKY130_FD_SC_HDLL__A32OI_1%A_27_297# N_A_27_297#_M1002_s
+ N_A_27_297#_M1000_d N_A_27_297#_M1003_d N_A_27_297#_c_193_n
+ N_A_27_297#_c_194_n N_A_27_297#_c_197_n N_A_27_297#_c_201_n
+ N_A_27_297#_c_203_n N_A_27_297#_c_206_n N_A_27_297#_c_210_n
+ PM_SKY130_FD_SC_HDLL__A32OI_1%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A32OI_1%Y N_Y_M1001_d N_Y_M1002_d N_Y_c_239_n
+ N_Y_c_233_n N_Y_c_234_n Y Y PM_SKY130_FD_SC_HDLL__A32OI_1%Y
x_PM_SKY130_FD_SC_HDLL__A32OI_1%VPWR N_VPWR_M1007_d N_VPWR_M1008_d
+ N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n
+ N_VPWR_c_273_n N_VPWR_c_274_n VPWR N_VPWR_c_267_n
+ PM_SKY130_FD_SC_HDLL__A32OI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A32OI_1%VGND N_VGND_M1005_s N_VGND_M1006_d
+ N_VGND_c_307_n N_VGND_c_308_n N_VGND_c_309_n N_VGND_c_310_n N_VGND_c_311_n
+ N_VGND_c_312_n VGND N_VGND_c_313_n PM_SKY130_FD_SC_HDLL__A32OI_1%VGND
cc_1 VNB N_B2_c_49_n 0.0215673f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB B2 0.0156742f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_B2_c_51_n 0.039201f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_B1_c_75_n 0.0184367f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B1_c_76_n 0.0238712f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_B1_c_77_n 0.00424984f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_7 VNB N_A1_c_107_n 0.025064f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_A1_c_108_n 0.0177301f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB A1 0.00140451f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_10 VNB N_A2_c_139_n 0.0163651f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_A2_c_140_n 0.024438f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_12 VNB A2 0.00115519f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_13 VNB N_A3_c_170_n 0.0138067f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_14 VNB N_A3_c_171_n 0.0189423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A3_c_172_n 0.00202312f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_16 VNB A3 0.0165221f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_17 VNB N_A3_c_174_n 0.0120039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB Y 0.00288657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_267_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_307_n 0.0120242f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_21 VNB N_VGND_c_308_n 0.0145569f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.202
cc_22 VNB N_VGND_c_309_n 0.0280734f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_23 VNB N_VGND_c_310_n 0.0162079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_311_n 0.0589181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_312_n 0.0062884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_313_n 0.180776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VPB N_B2_c_52_n 0.020812f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_28 VPB B2 0.00454807f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_29 VPB N_B2_c_51_n 0.019138f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_30 VPB N_B1_c_76_n 0.0268861f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_31 VPB N_B1_c_77_n 0.00190262f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_32 VPB N_A1_c_107_n 0.027128f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_33 VPB A1 2.71883e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_34 VPB N_A2_c_140_n 0.0256736f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_35 VPB A2 2.71883e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_36 VPB N_A3_c_172_n 0.0323326f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_37 VPB A3 0.00419012f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_38 VPB N_A_27_297#_c_193_n 0.00929745f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_39 VPB N_A_27_297#_c_194_n 0.0165453f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_40 VPB Y 0.00105909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_268_n 0.00456071f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.202
cc_42 VPB N_VPWR_c_269_n 0.0433467f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_43 VPB N_VPWR_c_270_n 0.043319f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_271_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_272_n 0.0108943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_273_n 0.0164023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_274_n 0.00593702f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_267_n 0.0508213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 N_B2_c_49_n N_B1_c_75_n 0.0295873f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_50 N_B2_c_52_n N_B1_c_76_n 0.0343508f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 N_B2_c_51_n N_B1_c_76_n 0.0295873f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_52 N_B2_c_51_n N_B1_c_77_n 3.44518e-19 $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_53 B2 N_A_27_297#_c_194_n 0.00920024f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_54 N_B2_c_51_n N_A_27_297#_c_194_n 0.00155795f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_55 N_B2_c_52_n N_A_27_297#_c_197_n 0.0134476f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_56 N_B2_c_49_n N_Y_c_233_n 0.0125163f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_57 N_B2_c_49_n N_Y_c_234_n 0.00139501f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_58 N_B2_c_52_n Y 0.0281369f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_59 N_B2_c_49_n Y 0.0102688f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_60 B2 Y 0.0238764f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_61 N_B2_c_51_n Y 0.0145635f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_62 N_B2_c_52_n N_VPWR_c_270_n 0.00429453f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_B2_c_52_n N_VPWR_c_267_n 0.00700261f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_64 N_B2_c_49_n N_VGND_c_308_n 0.00495469f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_65 B2 N_VGND_c_308_n 0.00785389f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_66 N_B2_c_51_n N_VGND_c_308_n 0.00357774f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_67 N_B2_c_49_n N_VGND_c_311_n 0.00499818f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_68 N_B2_c_49_n N_VGND_c_313_n 0.00889408f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_69 N_B1_c_76_n N_A1_c_107_n 0.0367193f $X=0.965 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_70 N_B1_c_77_n N_A1_c_107_n 0.00859889f $X=1.03 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_71 N_B1_c_75_n N_A1_c_108_n 0.0132856f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_72 N_B1_c_75_n A1 0.00404323f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_73 N_B1_c_76_n A1 3.50991e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 N_B1_c_77_n A1 0.019417f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_75 N_B1_c_77_n N_A_27_297#_M1000_d 0.00395702f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B1_c_76_n N_A_27_297#_c_197_n 0.0157706f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_77 N_B1_c_77_n N_A_27_297#_c_197_n 0.0052576f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B1_c_76_n N_A_27_297#_c_201_n 0.00182998f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_79 N_B1_c_77_n N_A_27_297#_c_201_n 0.00349239f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B1_c_76_n N_A_27_297#_c_203_n 0.0055061f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_81 N_B1_c_75_n N_Y_c_239_n 0.0122184f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_82 N_B1_c_76_n N_Y_c_239_n 9.59713e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B1_c_77_n N_Y_c_239_n 0.0201443f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B1_c_75_n N_Y_c_234_n 0.00765495f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B1_c_75_n Y 0.00765128f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_86 N_B1_c_76_n Y 0.0126884f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_87 N_B1_c_77_n Y 0.0474677f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_88 N_B1_c_76_n N_VPWR_c_270_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B1_c_76_n N_VPWR_c_267_n 0.00650299f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B1_c_75_n N_VGND_c_311_n 0.00406829f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B1_c_75_n N_VGND_c_313_n 0.00625696f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A1_c_108_n N_A2_c_139_n 0.0290065f $X=1.62 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_93 A1 N_A2_c_139_n 0.00363063f $X=1.5 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_94 N_A1_c_107_n N_A2_c_140_n 0.0677313f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A1_c_108_n A2 0.00305445f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_96 A1 A2 0.0415228f $X=1.5 $Y=0.425 $X2=0 $Y2=0
cc_97 N_A1_c_107_n N_A_27_297#_c_201_n 6.50343e-19 $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A1_c_107_n N_A_27_297#_c_203_n 0.00460856f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A1_c_107_n N_A_27_297#_c_206_n 0.0130084f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_100 A1 N_A_27_297#_c_206_n 0.00679426f $X=1.5 $Y=0.425 $X2=0 $Y2=0
cc_101 A1 N_Y_M1001_d 0.00608208f $X=1.5 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_102 N_A1_c_108_n N_Y_c_239_n 7.03273e-19 $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_103 A1 N_Y_c_239_n 0.0120269f $X=1.5 $Y=0.425 $X2=0 $Y2=0
cc_104 N_A1_c_108_n N_Y_c_234_n 0.00215355f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_105 A1 N_Y_c_234_n 0.0191343f $X=1.5 $Y=0.425 $X2=0 $Y2=0
cc_106 N_A1_c_107_n N_VPWR_c_268_n 0.00300743f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A1_c_107_n N_VPWR_c_270_n 0.00702461f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A1_c_107_n N_VPWR_c_267_n 0.00731696f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A1_c_108_n N_VGND_c_311_n 0.0037719f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_110 A1 N_VGND_c_311_n 0.00820582f $X=1.5 $Y=0.425 $X2=0 $Y2=0
cc_111 N_A1_c_108_n N_VGND_c_313_n 0.00589832f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_112 A1 N_VGND_c_313_n 0.00728499f $X=1.5 $Y=0.425 $X2=0 $Y2=0
cc_113 N_A2_c_140_n N_A3_c_170_n 0.0202968f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_114 A2 N_A3_c_170_n 4.5144e-19 $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_115 N_A2_c_139_n N_A3_c_171_n 0.0316243f $X=2.04 $Y=0.995 $X2=0 $Y2=0
cc_116 A2 N_A3_c_171_n 0.00656315f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_117 N_A2_c_140_n N_A3_c_172_n 0.0243911f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A2_c_140_n A3 0.00198797f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_119 A2 A3 0.0211854f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_120 N_A2_c_140_n N_A_27_297#_c_206_n 0.013235f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_121 A2 N_A_27_297#_c_206_n 0.00625303f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_122 N_A2_c_140_n N_A_27_297#_c_210_n 6.82445e-19 $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A2_c_140_n N_VPWR_c_268_n 0.00159434f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A2_c_140_n N_VPWR_c_269_n 0.00187208f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A2_c_140_n N_VPWR_c_273_n 0.00702461f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A2_c_140_n N_VPWR_c_267_n 0.00700869f $X=2.065 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A2_c_139_n N_VGND_c_309_n 0.00220259f $X=2.04 $Y=0.995 $X2=0 $Y2=0
cc_128 A2 N_VGND_c_309_n 0.0157264f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_129 N_A2_c_139_n N_VGND_c_311_n 0.00416396f $X=2.04 $Y=0.995 $X2=0 $Y2=0
cc_130 A2 N_VGND_c_311_n 0.00567082f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_131 N_A2_c_139_n N_VGND_c_313_n 0.00637074f $X=2.04 $Y=0.995 $X2=0 $Y2=0
cc_132 A2 N_VGND_c_313_n 0.00631895f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_133 A2 A_423_47# 0.00595534f $X=2.015 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_134 N_A3_c_172_n N_VPWR_c_269_n 0.0264811f $X=2.58 $Y=1.41 $X2=0 $Y2=0
cc_135 A3 N_VPWR_c_269_n 0.0223625f $X=2.5 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A3_c_172_n N_VPWR_c_273_n 0.00388479f $X=2.58 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A3_c_172_n N_VPWR_c_267_n 0.00676216f $X=2.58 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A3_c_170_n N_VGND_c_309_n 0.00298992f $X=2.58 $Y=1.095 $X2=0 $Y2=0
cc_139 N_A3_c_171_n N_VGND_c_309_n 0.0156602f $X=2.58 $Y=0.96 $X2=0 $Y2=0
cc_140 A3 N_VGND_c_309_n 0.0181349f $X=2.5 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A3_c_171_n N_VGND_c_311_n 0.00486043f $X=2.58 $Y=0.96 $X2=0 $Y2=0
cc_142 N_A3_c_171_n N_VGND_c_313_n 0.00844905f $X=2.58 $Y=0.96 $X2=0 $Y2=0
cc_143 N_A_27_297#_c_197_n N_Y_M1002_d 0.00355156f $X=1.195 $Y=2.36 $X2=0 $Y2=0
cc_144 N_A_27_297#_c_194_n Y 0.0193539f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_145 N_A_27_297#_c_197_n Y 0.0202507f $X=1.195 $Y=2.36 $X2=0 $Y2=0
cc_146 N_A_27_297#_c_201_n Y 0.00966852f $X=1.32 $Y=1.955 $X2=0 $Y2=0
cc_147 N_A_27_297#_c_203_n Y 0.00677711f $X=1.32 $Y=2.255 $X2=0 $Y2=0
cc_148 N_A_27_297#_c_206_n N_VPWR_M1007_d 0.0085927f $X=2.215 $Y=1.87 $X2=-0.19
+ $Y2=1.305
cc_149 N_A_27_297#_c_206_n N_VPWR_c_268_n 0.0132478f $X=2.215 $Y=1.87 $X2=0
+ $Y2=0
cc_150 N_A_27_297#_c_210_n N_VPWR_c_269_n 0.0553287f $X=2.3 $Y=1.91 $X2=0 $Y2=0
cc_151 N_A_27_297#_c_193_n N_VPWR_c_270_n 0.0182136f $X=0.215 $Y=2.255 $X2=0
+ $Y2=0
cc_152 N_A_27_297#_c_197_n N_VPWR_c_270_n 0.0472019f $X=1.195 $Y=2.36 $X2=0
+ $Y2=0
cc_153 N_A_27_297#_c_203_n N_VPWR_c_270_n 0.0175802f $X=1.32 $Y=2.255 $X2=0
+ $Y2=0
cc_154 N_A_27_297#_c_210_n N_VPWR_c_273_n 0.0118637f $X=2.3 $Y=1.91 $X2=0 $Y2=0
cc_155 N_A_27_297#_M1002_s N_VPWR_c_267_n 0.00217523f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_156 N_A_27_297#_M1000_d N_VPWR_c_267_n 0.00394925f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_157 N_A_27_297#_M1003_d N_VPWR_c_267_n 0.00514355f $X=2.155 $Y=1.485 $X2=0
+ $Y2=0
cc_158 N_A_27_297#_c_193_n N_VPWR_c_267_n 0.00998795f $X=0.215 $Y=2.255 $X2=0
+ $Y2=0
cc_159 N_A_27_297#_c_197_n N_VPWR_c_267_n 0.0300764f $X=1.195 $Y=2.36 $X2=0
+ $Y2=0
cc_160 N_A_27_297#_c_203_n N_VPWR_c_267_n 0.00962794f $X=1.32 $Y=2.255 $X2=0
+ $Y2=0
cc_161 N_A_27_297#_c_206_n N_VPWR_c_267_n 0.0170503f $X=2.215 $Y=1.87 $X2=0
+ $Y2=0
cc_162 N_A_27_297#_c_210_n N_VPWR_c_267_n 0.00647979f $X=2.3 $Y=1.91 $X2=0 $Y2=0
cc_163 N_Y_M1002_d N_VPWR_c_267_n 0.00232895f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_164 N_Y_c_239_n N_VGND_c_311_n 0.00275741f $X=0.965 $Y=0.72 $X2=0 $Y2=0
cc_165 N_Y_c_233_n N_VGND_c_311_n 0.00437317f $X=0.775 $Y=0.72 $X2=0 $Y2=0
cc_166 N_Y_c_234_n N_VGND_c_311_n 0.0147442f $X=1.18 $Y=0.53 $X2=0 $Y2=0
cc_167 N_Y_M1001_d N_VGND_c_313_n 0.0116883f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_168 N_Y_c_239_n N_VGND_c_313_n 0.00487344f $X=0.965 $Y=0.72 $X2=0 $Y2=0
cc_169 N_Y_c_233_n N_VGND_c_313_n 0.00741246f $X=0.775 $Y=0.72 $X2=0 $Y2=0
cc_170 N_Y_c_234_n N_VGND_c_313_n 0.0109258f $X=1.18 $Y=0.53 $X2=0 $Y2=0
cc_171 N_Y_c_239_n A_119_47# 0.00177909f $X=0.965 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_172 N_Y_c_233_n A_119_47# 0.00224858f $X=0.775 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_173 Y A_119_47# 9.24014e-19 $X=0.645 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_174 N_VGND_c_313_n A_119_47# 0.0031505f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_175 N_VGND_c_313_n A_339_47# 0.0115413f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_176 N_VGND_c_313_n A_423_47# 0.0117715f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
