* File: sky130_fd_sc_hdll__xor2_2.spice
* Created: Thu Aug 27 19:29:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__xor2_2.pex.spice"
.subckt sky130_fd_sc_hdll__xor2_2  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_112_47#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.12025 PD=1.85 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_M1015_g N_A_112_47#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1015_d N_B_M1016_g N_A_112_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1017_d N_B_M1017_g N_A_112_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_510_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1003_d N_A_M1007_g N_A_510_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1000 N_X_M1000_d N_B_M1000_g N_A_510_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.138125 AS=0.104 PD=1.075 PS=0.97 NRD=18.456 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1000_d N_B_M1004_g N_A_510_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.138125 AS=0.169 PD=1.075 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_112_47#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_112_47#_M1012_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.285 PD=1.29 PS=2.57 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1001_d N_A_M1013_g N_A_27_297#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1006 N_A_27_297#_M1013_s N_B_M1006_g N_A_112_47#_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1009_d N_B_M1009_g N_A_112_47#_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1018 N_A_510_297#_M1018_d N_A_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1019 N_A_510_297#_M1019_d N_A_M1019_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_510_297#_M1019_d N_B_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.1725 PD=1.29 PS=1.345 NRD=0.9653 NRS=11.8003 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_A_510_297#_M1010_d N_B_M1010_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.1725 PD=2.54 PS=1.345 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1011 N_A_510_297#_M1011_d N_A_112_47#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1014 N_A_510_297#_M1014_d N_A_112_47#_M1014_g N_X_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
*
.include "sky130_fd_sc_hdll__xor2_2.pxi.spice"
*
.ends
*
*
