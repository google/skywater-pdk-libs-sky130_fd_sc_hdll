* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VGND a_1787_159# a_2181_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND a_2266_413# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_455_324# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X3 VPWR a_1611_413# a_1787_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=180000u
X4 Q_N a_851_264# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_955_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X7 VGND SCD a_1373_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_2266_413# a_211_363# a_2360_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X9 a_851_264# a_2266_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR DE a_787_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X11 VPWR a_2266_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_787_369# a_851_264# a_319_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X13 a_2414_47# a_851_264# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_413_47# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_27_47# a_211_363# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_455_324# a_779_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_985_47# a_27_47# a_1611_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X18 a_1738_47# a_1787_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_851_264# a_2266_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X20 VPWR SCD a_1376_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X21 a_985_47# a_211_363# a_1611_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X22 Q a_2266_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_2165_413# a_27_47# a_2266_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X24 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_1611_413# a_1787_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 a_319_47# SCE a_985_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X27 Q_N a_851_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_455_324# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VGND a_851_264# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VPWR a_27_47# a_211_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X31 a_1611_413# a_27_47# a_1712_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X32 a_319_47# D a_413_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_319_47# a_955_21# a_985_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1611_413# a_211_363# a_1738_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X35 a_409_369# a_455_324# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X36 a_955_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X37 a_2181_47# a_211_363# a_2266_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X38 a_779_47# a_851_264# a_319_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1712_413# a_1787_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X40 a_2360_413# a_851_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X41 Q a_2266_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X42 a_2266_413# a_27_47# a_2414_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X43 a_319_47# D a_409_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X44 VPWR a_1787_159# a_2165_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X45 a_1376_369# a_955_21# a_985_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X46 a_1373_119# SCE a_985_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X47 VPWR a_851_264# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
