* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_805_297# B1 a_523_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_79_204# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_1243_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND C1 a_79_204# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND B1 a_79_204# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_79_204# C1 a_805_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VPWR A1 a_523_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_523_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VPWR A2 a_523_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_79_204# A1 a_1243_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A2 a_1051_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_523_297# B1 a_613_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 a_613_297# C1 a_79_204# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_523_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_79_204# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_1051_47# A1 a_79_204# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
