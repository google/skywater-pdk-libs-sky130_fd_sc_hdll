# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a22o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a22o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.350000 1.075000 5.895000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 1.075000 5.130000 1.445000 ;
        RECT 4.750000 1.445000 6.285000 1.615000 ;
        RECT 6.115000 1.075000 6.815000 1.275000 ;
        RECT 6.115000 1.275000 6.285000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 1.075000 4.030000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.620000 1.075000 3.205000 1.445000 ;
        RECT 2.620000 1.445000 4.580000 1.615000 ;
        RECT 4.200000 1.075000 4.580000 1.445000 ;
    END
  END B2
  PIN VGND
    ANTENNADIFFAREA  1.397500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.900000 0.085000 ;
        RECT 0.260000  0.085000 0.430000 0.555000 ;
        RECT 1.200000  0.085000 1.370000 0.555000 ;
        RECT 2.140000  0.085000 2.830000 0.555000 ;
        RECT 4.585000  0.085000 4.755000 0.555000 ;
        RECT 6.500000  0.085000 6.670000 0.895000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.430000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.900000 2.805000 ;
        RECT 0.220000 1.825000 0.470000 2.635000 ;
        RECT 1.160000 1.795000 1.410000 2.635000 ;
        RECT 2.100000 2.125000 2.350000 2.635000 ;
        RECT 5.050000 2.125000 5.300000 2.635000 ;
        RECT 5.990000 2.125000 6.240000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.725000 1.920000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.445000 ;
        RECT 0.085000 1.445000 1.880000 1.615000 ;
        RECT 0.600000 0.265000 0.980000 0.725000 ;
        RECT 0.690000 1.615000 0.940000 2.465000 ;
        RECT 1.540000 0.255000 1.920000 0.725000 ;
        RECT 1.630000 1.615000 1.880000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.540000 1.075000 2.430000 1.275000 ;
      RECT 2.100000 1.275000 2.430000 1.785000 ;
      RECT 2.100000 1.785000 4.280000 1.955000 ;
      RECT 2.140000 0.735000 5.810000 0.905000 ;
      RECT 2.140000 0.905000 2.430000 1.075000 ;
      RECT 2.620000 2.125000 2.870000 2.295000 ;
      RECT 2.620000 2.295000 4.830000 2.465000 ;
      RECT 3.000000 0.255000 4.320000 0.475000 ;
      RECT 3.090000 1.955000 3.340000 2.125000 ;
      RECT 3.420000 0.645000 3.905000 0.735000 ;
      RECT 3.560000 2.125000 3.810000 2.295000 ;
      RECT 4.030000 1.955000 4.280000 2.125000 ;
      RECT 4.500000 1.785000 6.710000 1.955000 ;
      RECT 4.500000 1.955000 4.830000 2.295000 ;
      RECT 4.960000 0.255000 6.280000 0.475000 ;
      RECT 5.385000 0.645000 5.810000 0.735000 ;
      RECT 5.520000 1.955000 5.770000 2.465000 ;
      RECT 6.030000 0.475000 6.280000 0.895000 ;
      RECT 6.505000 1.455000 6.710000 1.785000 ;
      RECT 6.505000 1.955000 6.710000 2.465000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22o_4
