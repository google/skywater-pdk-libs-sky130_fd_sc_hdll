* File: sky130_fd_sc_hdll__buf_8.pex.spice
* Created: Thu Aug 27 19:00:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUF_8%A 1 3 6 8 10 13 15 17 20 22 23 24 38 45 47
c68 24 0 1.25463e-19 $X=1.065 $Y=1.105
r69 45 47 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=1.035 $Y2=1.175
r70 38 39 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.212
+ $X2=1.46 $Y2=1.212
r71 36 38 59.5062 $w=3.24e-07 $l=4e-07 $layer=POLY_cond $X=1.035 $Y=1.212
+ $X2=1.435 $Y2=1.212
r72 36 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.035
+ $Y=1.16 $X2=1.035 $Y2=1.16
r73 34 36 6.69444 $w=3.24e-07 $l=4.5e-08 $layer=POLY_cond $X=0.99 $Y=1.212
+ $X2=1.035 $Y2=1.212
r74 33 34 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.212
+ $X2=0.99 $Y2=1.212
r75 32 33 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.212
+ $X2=0.965 $Y2=1.212
r76 31 32 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.212
+ $X2=0.52 $Y2=1.212
r77 29 31 28.2654 $w=3.24e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.212
+ $X2=0.495 $Y2=1.212
r78 24 47 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=1.15 $Y=1.175
+ $X2=1.035 $Y2=1.175
r79 23 45 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=0.685 $Y=1.175
+ $X2=0.695 $Y2=1.175
r80 22 23 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.685 $Y2=1.175
r81 22 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.305
+ $Y=1.16 $X2=0.305 $Y2=1.16
r82 18 39 20.7868 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.212
r83 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r84 15 38 16.5046 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.212
r85 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r86 11 34 20.7868 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=1.212
r87 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=0.56
r88 8 33 16.5046 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.212
r89 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r90 4 32 20.7868 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=1.212
r91 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=0.56
r92 1 31 16.5046 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.212
r93 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_8%A_27_47# 1 2 3 4 15 17 19 22 24 26 29 31 33
+ 36 38 40 43 45 47 50 52 54 57 59 61 62 64 67 71 77 79 80 81 82 85 91 93 95 98
+ 100 106 109 110 111 128
c229 128 0 1.25463e-19 $X=5.195 $Y=1.217
c230 52 0 1.89091e-19 $X=4.255 $Y=1.41
r231 128 129 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=5.195 $Y=1.217
+ $X2=5.22 $Y2=1.217
r232 127 128 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=4.725 $Y=1.217
+ $X2=5.195 $Y2=1.217
r233 126 127 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.217
+ $X2=4.725 $Y2=1.217
r234 123 124 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.217
+ $X2=4.255 $Y2=1.217
r235 122 123 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=3.785 $Y=1.217
+ $X2=4.23 $Y2=1.217
r236 121 122 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.217
+ $X2=3.785 $Y2=1.217
r237 120 121 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=3.315 $Y=1.217
+ $X2=3.76 $Y2=1.217
r238 119 120 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.217
+ $X2=3.315 $Y2=1.217
r239 118 119 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=3.29 $Y2=1.217
r240 117 118 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.217
+ $X2=2.845 $Y2=1.217
r241 116 117 66.6118 $w=3.22e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.82 $Y2=1.217
r242 115 116 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r243 112 113 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.217
+ $X2=1.905 $Y2=1.217
r244 107 126 62.8696 $w=3.22e-07 $l=4.2e-07 $layer=POLY_cond $X=4.28 $Y=1.217
+ $X2=4.7 $Y2=1.217
r245 107 124 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.217
+ $X2=4.255 $Y2=1.217
r246 106 107 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=4.28
+ $Y=1.16 $X2=4.28 $Y2=1.16
r247 104 115 53.8882 $w=3.22e-07 $l=3.6e-07 $layer=POLY_cond $X=1.99 $Y=1.217
+ $X2=2.35 $Y2=1.217
r248 104 113 12.7236 $w=3.22e-07 $l=8.5e-08 $layer=POLY_cond $X=1.99 $Y=1.217
+ $X2=1.905 $Y2=1.217
r249 103 106 149.401 $w=1.68e-07 $l=2.29e-06 $layer=LI1_cond $X=1.99 $Y=1.16
+ $X2=4.28 $Y2=1.16
r250 103 104 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=1.99
+ $Y=1.16 $X2=1.99 $Y2=1.16
r251 101 111 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=1.745 $Y=1.16
+ $X2=1.657 $Y2=1.16
r252 101 103 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.745 $Y=1.16
+ $X2=1.99 $Y2=1.16
r253 99 111 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.657 $Y=1.245
+ $X2=1.657 $Y2=1.16
r254 99 100 12.6753 $w=1.73e-07 $l=2e-07 $layer=LI1_cond $X=1.657 $Y=1.245
+ $X2=1.657 $Y2=1.445
r255 98 111 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.657 $Y=1.075
+ $X2=1.657 $Y2=1.16
r256 97 98 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=1.657 $Y=0.905
+ $X2=1.657 $Y2=1.075
r257 96 109 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=1.53
+ $X2=1.175 $Y2=1.53
r258 95 100 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.57 $Y=1.53
+ $X2=1.657 $Y2=1.445
r259 95 96 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.57 $Y=1.53
+ $X2=1.365 $Y2=1.53
r260 94 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0.82
+ $X2=1.2 $Y2=0.82
r261 93 97 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.57 $Y=0.82
+ $X2=1.657 $Y2=0.905
r262 93 94 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.57 $Y=0.82
+ $X2=1.285 $Y2=0.82
r263 89 110 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.2 $Y2=0.82
r264 89 91 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.2 $Y2=0.56
r265 85 87 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.175 $Y=1.63
+ $X2=1.175 $Y2=2.31
r266 83 109 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=1.615
+ $X2=1.175 $Y2=1.53
r267 83 85 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.175 $Y=1.615
+ $X2=1.175 $Y2=1.63
r268 81 109 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=1.53
+ $X2=1.175 $Y2=1.53
r269 81 82 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=1.53
+ $X2=0.425 $Y2=1.53
r270 79 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.82
+ $X2=1.2 $Y2=0.82
r271 79 80 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0.82
+ $X2=0.345 $Y2=0.82
r272 75 80 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.345 $Y2=0.82
r273 75 77 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.56
r274 71 73 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r275 69 82 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.425 $Y2=1.53
r276 69 71 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.63
r277 65 129 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.22 $Y=1.025
+ $X2=5.22 $Y2=1.217
r278 65 67 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.22 $Y=1.025
+ $X2=5.22 $Y2=0.56
r279 62 128 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.217
r280 62 64 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r281 59 127 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.217
r282 59 61 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r283 55 126 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=1.217
r284 55 57 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=0.56
r285 52 124 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.217
r286 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r287 48 123 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=1.217
r288 48 50 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=0.56
r289 45 122 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.217
r290 45 47 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r291 41 121 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.76 $Y=1.025
+ $X2=3.76 $Y2=1.217
r292 41 43 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.76 $Y=1.025
+ $X2=3.76 $Y2=0.56
r293 38 120 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r294 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r295 34 119 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r296 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r297 31 118 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r298 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r299 27 117 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=1.217
r300 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=0.56
r301 24 116 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r302 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r303 20 115 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r304 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
r305 17 113 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r306 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r307 13 112 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=1.217
r308 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=0.56
r309 4 87 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.31
r310 4 85 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.63
r311 3 73 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r312 3 71 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r313 2 91 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.56
r314 1 77 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_8%VPWR 1 2 3 4 5 6 21 23 27 31 35 39 41 45 49
+ 51 53 58 63 70 71 73 75 78 81 84 87 90
r103 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r104 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r105 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r106 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r108 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r109 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r110 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.645 $Y=2.72
+ $X2=0.73 $Y2=2.72
r112 71 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r113 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r114 68 90 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=5.405 $Y2=2.72
r115 68 70 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=5.75 $Y2=2.72
r116 67 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r117 67 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r118 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r119 64 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.525 $Y2=2.72
r120 64 66 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.91 $Y2=2.72
r121 63 87 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.275 $Y=2.72
+ $X2=4.465 $Y2=2.72
r122 63 66 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.275 $Y=2.72
+ $X2=3.91 $Y2=2.72
r123 62 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r124 62 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r125 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r126 59 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.585 $Y2=2.72
r127 59 61 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.99 $Y2=2.72
r128 58 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=3.525 $Y2=2.72
r129 58 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=2.99 $Y2=2.72
r130 57 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r131 57 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r132 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r133 54 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=2.72
+ $X2=1.67 $Y2=2.72
r134 54 56 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.755 $Y=2.72
+ $X2=2.07 $Y2=2.72
r135 53 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.585 $Y2=2.72
r136 53 56 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.07 $Y2=2.72
r137 51 76 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r138 49 73 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.235 $Y=2.72
+ $X2=0.645 $Y2=2.72
r139 45 48 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=5.405 $Y=1.66
+ $X2=5.405 $Y2=2.34
r140 43 90 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.405 $Y=2.635
+ $X2=5.405 $Y2=2.72
r141 43 48 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=5.405 $Y=2.635
+ $X2=5.405 $Y2=2.34
r142 42 87 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.655 $Y=2.72
+ $X2=4.465 $Y2=2.72
r143 41 90 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.215 $Y=2.72
+ $X2=5.405 $Y2=2.72
r144 41 42 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.215 $Y=2.72
+ $X2=4.655 $Y2=2.72
r145 37 87 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=2.635
+ $X2=4.465 $Y2=2.72
r146 37 39 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=4.465 $Y=2.635
+ $X2=4.465 $Y2=2
r147 33 84 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=2.635
+ $X2=3.525 $Y2=2.72
r148 33 35 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.525 $Y=2.635
+ $X2=3.525 $Y2=2
r149 29 81 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=2.635
+ $X2=2.585 $Y2=2.72
r150 29 31 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.585 $Y=2.635
+ $X2=2.585 $Y2=2
r151 25 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r152 25 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2
r153 24 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.73 $Y2=2.72
r154 23 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=1.67 $Y2=2.72
r155 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=0.815 $Y2=2.72
r156 19 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r157 19 21 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2
r158 6 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.34
r159 6 45 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.66
r160 5 39 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2
r161 4 35 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2
r162 3 31 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2
r163 2 27 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2
r164 1 21 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_8%X 1 2 3 4 5 6 7 8 27 31 33 34 35 36 39 43 45
+ 47 51 55 57 59 63 65 66 67 68 69 70 71 86
c139 69 0 1.89091e-19 $X=4.825 $Y=0.85
r140 71 86 7.82882 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=4.96 $Y=1.615
+ $X2=4.96 $Y2=1.755
r141 70 71 7.06976 $w=5.23e-07 $l=2.55e-07 $layer=LI1_cond $X=4.867 $Y=1.19
+ $X2=4.867 $Y2=1.445
r142 69 78 3.55013 $w=2.62e-07 $l=8.5e-08 $layer=LI1_cond $X=4.867 $Y=0.82
+ $X2=4.867 $Y2=0.905
r143 69 70 8.76506 $w=3.53e-07 $l=2.7e-07 $layer=LI1_cond $X=4.867 $Y=0.92
+ $X2=4.867 $Y2=1.19
r144 69 78 0.486948 $w=3.53e-07 $l=1.5e-08 $layer=LI1_cond $X=4.867 $Y=0.92
+ $X2=4.867 $Y2=0.905
r145 61 69 3.55013 $w=2.62e-07 $l=1.28662e-07 $layer=LI1_cond $X=4.96 $Y=0.735
+ $X2=4.867 $Y2=0.82
r146 61 63 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.96 $Y=0.735
+ $X2=4.96 $Y2=0.56
r147 60 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=1.53
+ $X2=4.02 $Y2=1.53
r148 59 71 2.9446 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=4.69 $Y=1.53
+ $X2=4.867 $Y2=1.53
r149 59 60 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.69 $Y=1.53
+ $X2=4.105 $Y2=1.53
r150 58 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=0.82
+ $X2=4.02 $Y2=0.82
r151 57 69 2.9446 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=4.69 $Y=0.82
+ $X2=4.867 $Y2=0.82
r152 57 58 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.69 $Y=0.82
+ $X2=4.105 $Y2=0.82
r153 53 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=1.615
+ $X2=4.02 $Y2=1.53
r154 53 55 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.02 $Y=1.615
+ $X2=4.02 $Y2=1.755
r155 49 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.735
+ $X2=4.02 $Y2=0.82
r156 49 51 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.02 $Y=0.735
+ $X2=4.02 $Y2=0.56
r157 48 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=1.53
+ $X2=3.08 $Y2=1.53
r158 47 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=1.53
+ $X2=4.02 $Y2=1.53
r159 47 48 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.935 $Y=1.53
+ $X2=3.165 $Y2=1.53
r160 46 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=0.82
+ $X2=3.08 $Y2=0.82
r161 45 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=0.82
+ $X2=4.02 $Y2=0.82
r162 45 46 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.935 $Y=0.82
+ $X2=3.165 $Y2=0.82
r163 41 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=1.615
+ $X2=3.08 $Y2=1.53
r164 41 43 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.08 $Y=1.615
+ $X2=3.08 $Y2=1.755
r165 37 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.735
+ $X2=3.08 $Y2=0.82
r166 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.08 $Y=0.735
+ $X2=3.08 $Y2=0.56
r167 35 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=1.53
+ $X2=3.08 $Y2=1.53
r168 35 36 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.995 $Y=1.53
+ $X2=2.225 $Y2=1.53
r169 33 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=0.82
+ $X2=3.08 $Y2=0.82
r170 33 34 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.995 $Y=0.82
+ $X2=2.225 $Y2=0.82
r171 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=1.615
+ $X2=2.225 $Y2=1.53
r172 29 31 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.14 $Y=1.615
+ $X2=2.14 $Y2=1.755
r173 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.225 $Y2=0.82
r174 25 27 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.14 $Y2=0.56
r175 8 86 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.755
r176 7 55 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.755
r177 6 43 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.755
r178 5 31 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.755
r179 4 63 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.56
r180 3 51 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.56
r181 2 39 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.56
r182 1 27 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_8%VGND 1 2 3 4 5 6 21 25 29 33 37 39 43 45 47
+ 49 54 56 61 66 71 78 79 82 85 88 91 94 97
r116 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r117 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r118 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r119 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r120 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r121 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r122 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r123 79 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r124 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r125 76 97 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.595 $Y=0 $X2=5.405
+ $Y2=0
r126 76 78 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.595 $Y=0
+ $X2=5.75 $Y2=0
r127 75 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r128 75 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r129 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r130 72 91 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.525
+ $Y2=0
r131 72 74 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.715 $Y=0
+ $X2=3.91 $Y2=0
r132 71 94 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.275 $Y=0 $X2=4.465
+ $Y2=0
r133 71 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.275 $Y=0
+ $X2=3.91 $Y2=0
r134 70 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r135 70 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r136 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r137 67 88 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.585
+ $Y2=0
r138 67 69 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.775 $Y=0
+ $X2=2.99 $Y2=0
r139 66 91 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=0 $X2=3.525
+ $Y2=0
r140 66 69 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.335 $Y=0 $X2=2.99
+ $Y2=0
r141 65 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r142 65 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r143 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r144 62 85 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.645
+ $Y2=0
r145 62 64 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.835 $Y=0
+ $X2=2.07 $Y2=0
r146 61 88 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.585
+ $Y2=0
r147 61 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=0
+ $X2=2.07 $Y2=0
r148 60 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r149 60 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r150 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r151 57 82 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r152 57 59 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r153 56 85 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.645
+ $Y2=0
r154 56 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r155 49 82 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r156 47 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r157 47 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r158 45 49 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.235 $Y=0
+ $X2=0.515 $Y2=0
r159 45 54 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r160 41 97 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.405 $Y=0.085
+ $X2=5.405 $Y2=0
r161 41 43 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=5.405 $Y=0.085
+ $X2=5.405 $Y2=0.38
r162 40 94 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=4.465
+ $Y2=0
r163 39 97 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.405
+ $Y2=0
r164 39 40 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.215 $Y=0
+ $X2=4.655 $Y2=0
r165 35 94 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=0.085
+ $X2=4.465 $Y2=0
r166 35 37 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=4.465 $Y=0.085
+ $X2=4.465 $Y2=0.4
r167 31 91 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0
r168 31 33 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0.4
r169 27 88 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.085
+ $X2=2.585 $Y2=0
r170 27 29 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.585 $Y=0.085
+ $X2=2.585 $Y2=0.4
r171 23 85 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0
r172 23 25 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0.4
r173 19 82 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r174 19 21 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.4
r175 6 43 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.295
+ $Y=0.235 $X2=5.43 $Y2=0.38
r176 5 37 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.4
r177 4 33 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.4
r178 3 29 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.4
r179 2 25 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.4
r180 1 21 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

