* File: sky130_fd_sc_hdll__einvp_2.pex.spice
* Created: Thu Aug 27 19:07:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EINVP_2%TE 3 6 7 9 10 11 12 14 15 17 19 20 21 22
c52 15 0 6.11783e-20 $X=1.39 $Y=1.035
r53 28 29 3.50291 $w=3.44e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.142
+ $X2=0.495 $Y2=1.142
r54 26 28 31.5262 $w=3.44e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.142
+ $X2=0.47 $Y2=1.142
r55 21 22 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.207 $Y=1.16
+ $X2=0.207 $Y2=1.53
r56 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r57 17 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.465 $Y=0.96
+ $X2=1.465 $Y2=0.56
r58 16 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.07 $Y=1.035
+ $X2=0.995 $Y2=1.035
r59 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.39 $Y=1.035
+ $X2=1.465 $Y2=0.96
r60 15 16 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.39 $Y=1.035
+ $X2=1.07 $Y2=1.035
r61 12 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.995 $Y=0.96
+ $X2=0.995 $Y2=1.035
r62 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.995 $Y=0.96
+ $X2=0.995 $Y2=0.56
r63 11 29 29.6109 $w=3.44e-07 $l=1.48825e-07 $layer=POLY_cond $X=0.595 $Y=1.035
+ $X2=0.495 $Y2=1.142
r64 10 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.92 $Y=1.035
+ $X2=0.995 $Y2=1.035
r65 10 11 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.92 $Y=1.035
+ $X2=0.595 $Y2=1.035
r66 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r67 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.67 $X2=0.495
+ $Y2=1.77
r68 5 29 15.449 $w=2e-07 $l=1.83e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.142
r69 5 6 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.67
r70 1 28 22.2144 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=0.47 $Y=0.96
+ $X2=0.47 $Y2=1.142
r71 1 3 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.47 $Y=0.96 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_2%A_27_47# 1 2 7 9 10 11 12 14 16 19 23 26
+ 27 29 30
c73 27 0 1.1096e-19 $X=0.925 $Y=1.16
r74 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.16 $X2=1.92 $Y2=1.16
r75 27 33 6.77082 $w=4.22e-07 $l=2.8562e-07 $layer=LI1_cond $X=0.925 $Y=1.16
+ $X2=0.712 $Y2=0.99
r76 27 29 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=0.925 $Y=1.16
+ $X2=1.92 $Y2=1.16
r77 25 33 0.687693 $w=4.25e-07 $l=3.35e-07 $layer=LI1_cond $X=0.712 $Y=1.325
+ $X2=0.712 $Y2=0.99
r78 25 26 12.4735 $w=4.23e-07 $l=4.6e-07 $layer=LI1_cond $X=0.712 $Y=1.325
+ $X2=0.712 $Y2=1.785
r79 21 26 32.4246 $w=1.68e-07 $l=4.97e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.712 $Y2=1.87
r80 21 23 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=1.955
+ $X2=0.215 $Y2=2.165
r81 17 33 14.3682 $w=4.22e-07 $l=6.43043e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.712 $Y2=0.99
r82 17 19 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r83 15 30 28.8521 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=1.945 $Y=1.32
+ $X2=1.945 $Y2=1.16
r84 15 16 13.0992 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.945 $Y=1.32
+ $X2=1.945 $Y2=1.395
r85 12 16 13.0992 $w=2.5e-07 $l=1.00623e-07 $layer=POLY_cond $X=2.005 $Y=1.47
+ $X2=1.945 $Y2=1.395
r86 12 14 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.005 $Y=1.47
+ $X2=2.005 $Y2=2.015
r87 10 16 12.7694 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.785 $Y=1.395
+ $X2=1.945 $Y2=1.395
r88 10 11 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.785 $Y=1.395
+ $X2=1.625 $Y2=1.395
r89 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.535 $Y=1.47
+ $X2=1.625 $Y2=1.395
r90 7 9 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.535 $Y=1.47
+ $X2=1.535 $Y2=2.015
r91 2 23 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.165
r92 1 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_2%A 1 3 4 6 7 9 10 12 13 14 15 22
r41 22 24 33.7665 $w=3.64e-07 $l=2.55e-07 $layer=POLY_cond $X=3.12 $Y=1.202
+ $X2=3.375 $Y2=1.202
r42 21 22 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=3.095 $Y=1.202
+ $X2=3.12 $Y2=1.202
r43 20 21 62.2363 $w=3.64e-07 $l=4.7e-07 $layer=POLY_cond $X=2.625 $Y=1.202
+ $X2=3.095 $Y2=1.202
r44 19 20 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=2.6 $Y=1.202
+ $X2=2.625 $Y2=1.202
r45 13 15 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.39 $Y=1.16
+ $X2=3.39 $Y2=1.53
r46 13 14 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=3.39 $Y=1.16
+ $X2=3.39 $Y2=0.85
r47 13 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.375
+ $Y=1.16 $X2=3.375 $Y2=1.16
r48 10 22 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.12 $Y=0.995
+ $X2=3.12 $Y2=1.202
r49 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.12 $Y=0.995
+ $X2=3.12 $Y2=0.56
r50 7 21 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.095 $Y=1.41
+ $X2=3.095 $Y2=1.202
r51 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.095 $Y=1.41
+ $X2=3.095 $Y2=1.985
r52 4 20 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.625 $Y=1.41
+ $X2=2.625 $Y2=1.202
r53 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.625 $Y=1.41
+ $X2=2.625 $Y2=1.985
r54 1 19 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.6 $Y=0.995 $X2=2.6
+ $Y2=1.202
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.6 $Y=0.995 $X2=2.6
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_2%VPWR 1 2 9 11 15 17 19 29 30 33 36
r47 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r51 27 30 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 26 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=2.72
+ $X2=1.77 $Y2=2.72
r56 24 26 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.935 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 19 33 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.72 $Y2=2.72
r58 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r59 17 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r60 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r61 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=2.635
+ $X2=1.77 $Y2=2.72
r62 13 15 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.77 $Y=2.635
+ $X2=1.77 $Y2=2.02
r63 12 33 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.72 $Y2=2.72
r64 11 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.77 $Y2=2.72
r65 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=0.925 $Y2=2.72
r66 7 33 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.635 $X2=0.72
+ $Y2=2.72
r67 7 9 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.34
r68 2 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.625
+ $Y=1.545 $X2=1.77 $Y2=2.02
r69 1 9 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.845 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_2%A_235_309# 1 2 3 12 14 15 19 20 21 24
c43 14 0 6.11783e-20 $X=2.185 $Y=1.64
r44 22 24 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=3.387 $Y=2.295
+ $X2=3.387 $Y2=1.96
r45 20 22 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=3.245 $Y=2.38
+ $X2=3.387 $Y2=2.295
r46 20 21 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.245 $Y=2.38
+ $X2=2.355 $Y2=2.38
r47 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.27 $Y=2.295
+ $X2=2.355 $Y2=2.38
r48 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.27 $Y=2.295
+ $X2=2.27 $Y2=1.96
r49 16 19 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.27 $Y=1.725
+ $X2=2.27 $Y2=1.96
r50 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.185 $Y=1.64
+ $X2=2.27 $Y2=1.725
r51 14 15 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=2.185 $Y=1.64
+ $X2=1.385 $Y2=1.64
r52 10 15 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.265 $Y=1.725
+ $X2=1.385 $Y2=1.64
r53 10 12 11.2843 $w=2.38e-07 $l=2.35e-07 $layer=LI1_cond $X=1.265 $Y=1.725
+ $X2=1.265 $Y2=1.96
r54 3 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.185
+ $Y=1.485 $X2=3.33 $Y2=1.96
r55 2 19 300 $w=1.7e-07 $l=4.94823e-07 $layer=licon1_PDIFF $count=2 $X=2.095
+ $Y=1.545 $X2=2.27 $Y2=1.96
r56 1 12 300 $w=1.7e-07 $l=4.73392e-07 $layer=licon1_PDIFF $count=2 $X=1.175
+ $Y=1.545 $X2=1.3 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_2%Z 1 2 7 8 9 10 16
r19 9 10 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.86 $Y=1.53 $X2=2.86
+ $Y2=1.87
r20 8 9 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.86 $Y=1.19 $X2=2.86
+ $Y2=1.53
r21 7 8 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.86 $Y=0.85 $X2=2.86
+ $Y2=1.19
r22 7 16 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=2.86 $Y=0.85 $X2=2.86
+ $Y2=0.76
r23 2 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.715
+ $Y=1.485 $X2=2.86 $Y2=1.61
r24 1 16 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=0.235 $X2=2.86 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_2%VGND 1 2 9 11 13 18 28 29 33 39
r50 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r51 33 36 10.119 $w=4.08e-07 $l=3.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.72
+ $Y2=0.36
r52 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r53 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r54 26 29 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r55 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r56 25 28 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r57 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r58 23 39 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.695
+ $Y2=0
r59 23 25 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.07
+ $Y2=0
r60 22 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r61 22 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r62 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r63 19 33 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.72
+ $Y2=0
r64 19 21 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.15
+ $Y2=0
r65 18 39 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.695
+ $Y2=0
r66 18 21 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.15
+ $Y2=0
r67 13 33 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.72
+ $Y2=0
r68 13 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r69 11 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r70 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r71 7 39 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0
r72 7 9 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0.38
r73 2 9 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.235 $X2=1.695 $Y2=0.38
r74 1 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.76 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_2%A_214_47# 1 2 3 12 14 15 19 20 21
r38 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.245 $Y=0.34
+ $X2=2.475 $Y2=0.34
r39 17 19 4.12815 $w=3.33e-07 $l=1.2e-07 $layer=LI1_cond $X=2.307 $Y=0.655
+ $X2=2.307 $Y2=0.535
r40 16 21 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=2.307 $Y=0.425
+ $X2=2.475 $Y2=0.34
r41 16 19 3.78414 $w=3.33e-07 $l=1.1e-07 $layer=LI1_cond $X=2.307 $Y=0.425
+ $X2=2.307 $Y2=0.535
r42 14 17 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=2.14 $Y=0.74
+ $X2=2.307 $Y2=0.655
r43 14 15 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=2.14 $Y=0.74 $X2=1.34
+ $Y2=0.74
r44 10 15 6.85817 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=1.242 $Y=0.655
+ $X2=1.34 $Y2=0.74
r45 10 12 6.82517 $w=1.93e-07 $l=1.2e-07 $layer=LI1_cond $X=1.242 $Y=0.655
+ $X2=1.242 $Y2=0.535
r46 3 20 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.235 $X2=3.33 $Y2=0.42
r47 2 19 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=2.17
+ $Y=0.235 $X2=2.295 $Y2=0.535
r48 1 12 182 $w=1.7e-07 $l=3.81445e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.255 $Y2=0.535
.ends

