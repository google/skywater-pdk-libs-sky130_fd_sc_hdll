# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__clkinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.664000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.035000 5.565000 1.290000 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA  0.701400 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  2.095000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  2.386400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.695000 6.330000 0.865000 ;
        RECT 0.115000 0.865000 0.285000 1.460000 ;
        RECT 0.115000 1.460000 6.330000 1.630000 ;
        RECT 0.615000 1.630000 0.855000 2.435000 ;
        RECT 1.555000 1.630000 1.795000 2.435000 ;
        RECT 1.685000 0.280000 1.875000 0.695000 ;
        RECT 2.495000 1.630000 2.745000 2.435000 ;
        RECT 2.645000 0.280000 2.835000 0.695000 ;
        RECT 3.430000 1.630000 3.675000 2.435000 ;
        RECT 3.605000 0.280000 3.795000 0.695000 ;
        RECT 4.420000 1.630000 4.725000 2.435000 ;
        RECT 4.665000 0.280000 4.855000 0.695000 ;
        RECT 5.465000 1.630000 5.705000 2.435000 ;
        RECT 6.060000 0.865000 6.330000 1.460000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.135000  1.800000 0.395000 2.635000 ;
      RECT 1.075000  1.800000 1.335000 2.635000 ;
      RECT 1.135000  0.085000 1.465000 0.525000 ;
      RECT 2.015000  1.800000 2.275000 2.635000 ;
      RECT 2.095000  0.085000 2.425000 0.525000 ;
      RECT 2.965000  1.800000 3.210000 2.635000 ;
      RECT 3.055000  0.085000 3.435000 0.525000 ;
      RECT 3.895000  1.800000 4.200000 2.635000 ;
      RECT 4.015000  0.085000 4.445000 0.525000 ;
      RECT 4.945000  1.800000 5.245000 2.635000 ;
      RECT 5.075000  0.085000 5.505000 0.525000 ;
      RECT 5.925000  1.800000 6.180000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_8
END LIBRARY
