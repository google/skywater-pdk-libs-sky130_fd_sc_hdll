* File: sky130_fd_sc_hdll__a21bo_4.pex.spice
* Created: Wed Sep  2 08:16:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21BO_4%B1_N 1 3 4 6 7 14
c31 1 0 1.15164e-19 $X=0.665 $Y=1.41
r32 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=1.16 $X2=0.635 $Y2=1.16
r33 7 14 0.972421 $w=6.13e-07 $l=5e-08 $layer=LI1_cond $X=0.685 $Y=1.317
+ $X2=0.635 $Y2=1.317
r34 4 10 38.578 $w=2.95e-07 $l=1.79374e-07 $layer=POLY_cond $X=0.69 $Y=0.995
+ $X2=0.66 $Y2=1.16
r35 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.69 $Y=0.995 $X2=0.69
+ $Y2=0.56
r36 1 10 48.1208 $w=2.95e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.665 $Y=1.41
+ $X2=0.66 $Y2=1.16
r37 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.665 $Y=1.41
+ $X2=0.665 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_4%A_209_21# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 40 41 42 45 49 51 54 60 72
c141 34 0 1.10898e-19 $X=2.585 $Y=1.16
c142 19 0 6.40318e-20 $X=1.625 $Y=1.41
r143 71 72 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.56 $Y=1.202
+ $X2=2.585 $Y2=1.202
r144 70 71 59.5951 $w=3.68e-07 $l=4.55e-07 $layer=POLY_cond $X=2.105 $Y=1.202
+ $X2=2.56 $Y2=1.202
r145 69 70 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.08 $Y=1.202
+ $X2=2.105 $Y2=1.202
r146 66 67 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.6 $Y=1.202
+ $X2=1.625 $Y2=1.202
r147 65 66 59.5951 $w=3.68e-07 $l=4.55e-07 $layer=POLY_cond $X=1.145 $Y=1.202
+ $X2=1.6 $Y2=1.202
r148 64 65 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.12 $Y=1.202
+ $X2=1.145 $Y2=1.202
r149 60 62 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=5.245 $Y=0.57
+ $X2=5.245 $Y2=0.755
r150 55 72 3.92935 $w=3.68e-07 $l=3e-08 $layer=POLY_cond $X=2.615 $Y=1.202
+ $X2=2.585 $Y2=1.202
r151 54 56 16.7054 $w=2.41e-07 $l=3.3e-07 $layer=LI1_cond $X=2.615 $Y=1.16
+ $X2=2.945 $Y2=1.16
r152 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.615
+ $Y=1.16 $X2=2.615 $Y2=1.16
r153 52 58 3.05 $w=1.7e-07 $l=9.80051e-08 $layer=LI1_cond $X=3.915 $Y=0.755
+ $X2=3.83 $Y2=0.727
r154 51 62 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.105 $Y=0.755
+ $X2=5.245 $Y2=0.755
r155 51 52 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=5.105 $Y=0.755
+ $X2=3.915 $Y2=0.755
r156 47 58 3.05 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.83 $Y=0.84 $X2=3.83
+ $Y2=0.727
r157 47 49 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.83 $Y=0.84
+ $X2=3.83 $Y2=1.62
r158 43 58 3.05 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.83 $Y=0.615 $X2=3.83
+ $Y2=0.727
r159 43 45 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.83 $Y=0.615
+ $X2=3.83 $Y2=0.42
r160 41 58 3.05 $w=1.7e-07 $l=9.75705e-08 $layer=LI1_cond $X=3.745 $Y=0.7
+ $X2=3.83 $Y2=0.727
r161 41 42 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.745 $Y=0.7
+ $X2=3.03 $Y2=0.7
r162 40 56 2.78154 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=0.995
+ $X2=2.945 $Y2=1.16
r163 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.945 $Y=0.785
+ $X2=3.03 $Y2=0.7
r164 39 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.945 $Y=0.785
+ $X2=2.945 $Y2=0.995
r165 37 69 25.5408 $w=3.68e-07 $l=1.95e-07 $layer=POLY_cond $X=1.885 $Y=1.202
+ $X2=2.08 $Y2=1.202
r166 37 67 34.0543 $w=3.68e-07 $l=2.6e-07 $layer=POLY_cond $X=1.885 $Y=1.202
+ $X2=1.625 $Y2=1.202
r167 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.885
+ $Y=1.16 $X2=1.885 $Y2=1.16
r168 34 54 2.01903 $w=3.3e-07 $l=3e-08 $layer=LI1_cond $X=2.585 $Y=1.16
+ $X2=2.615 $Y2=1.16
r169 34 36 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.585 $Y=1.16
+ $X2=1.885 $Y2=1.16
r170 31 72 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.585 $Y=1.41
+ $X2=2.585 $Y2=1.202
r171 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.585 $Y=1.41
+ $X2=2.585 $Y2=1.985
r172 28 71 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.56 $Y=0.995
+ $X2=2.56 $Y2=1.202
r173 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.56 $Y=0.995
+ $X2=2.56 $Y2=0.56
r174 25 70 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.105 $Y2=1.202
r175 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.105 $Y2=1.985
r176 22 69 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.08 $Y=0.995
+ $X2=2.08 $Y2=1.202
r177 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.08 $Y=0.995
+ $X2=2.08 $Y2=0.56
r178 19 67 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.625 $Y=1.41
+ $X2=1.625 $Y2=1.202
r179 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.625 $Y=1.41
+ $X2=1.625 $Y2=1.985
r180 16 66 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.6 $Y=0.995
+ $X2=1.6 $Y2=1.202
r181 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.6 $Y=0.995
+ $X2=1.6 $Y2=0.56
r182 13 65 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.145 $Y=1.41
+ $X2=1.145 $Y2=1.202
r183 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.145 $Y=1.41
+ $X2=1.145 $Y2=1.985
r184 10 64 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.12 $Y=0.995
+ $X2=1.12 $Y2=1.202
r185 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.12 $Y=0.995
+ $X2=1.12 $Y2=0.56
r186 3 49 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.685
+ $Y=1.485 $X2=3.83 $Y2=1.62
r187 2 60 182 $w=1.7e-07 $l=4.17373e-07 $layer=licon1_NDIFF $count=1 $X=5.055
+ $Y=0.235 $X2=5.24 $Y2=0.57
r188 1 58 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.235 $X2=3.83 $Y2=0.76
r189 1 45 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.235 $X2=3.83 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_4%A_36_47# 1 2 7 9 10 12 13 15 16 18 20 21
+ 24 25 27 31 36 46
c104 36 0 1.15164e-19 $X=0.32 $Y=2.02
c105 21 0 1.10898e-19 $X=2.92 $Y=2.02
c106 13 0 1.54054e-19 $X=4.065 $Y=1.41
r107 46 47 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=4.065 $Y=1.202
+ $X2=4.09 $Y2=1.202
r108 45 46 58.1274 $w=3.69e-07 $l=4.45e-07 $layer=POLY_cond $X=3.62 $Y=1.202
+ $X2=4.065 $Y2=1.202
r109 44 45 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=3.595 $Y=1.202
+ $X2=3.62 $Y2=1.202
r110 36 38 8.11401 $w=4.21e-07 $l=2.8e-07 $layer=LI1_cond $X=0.32 $Y=2.02
+ $X2=0.32 $Y2=2.3
r111 35 36 1.73872 $w=4.21e-07 $l=6e-08 $layer=LI1_cond $X=0.32 $Y=1.96 $X2=0.32
+ $Y2=2.02
r112 31 33 16.7678 $w=4.03e-07 $l=4.8e-07 $layer=LI1_cond $X=0.307 $Y=0.36
+ $X2=0.307 $Y2=0.84
r113 28 44 20.2466 $w=3.69e-07 $l=1.55e-07 $layer=POLY_cond $X=3.44 $Y=1.202
+ $X2=3.595 $Y2=1.202
r114 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.16 $X2=3.44 $Y2=1.16
r115 25 39 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.37 $Y=1.44
+ $X2=3.005 $Y2=1.44
r116 25 27 7.24924 $w=3.08e-07 $l=1.95e-07 $layer=LI1_cond $X=3.37 $Y=1.355
+ $X2=3.37 $Y2=1.16
r117 23 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=1.525
+ $X2=3.005 $Y2=1.44
r118 23 24 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.005 $Y=1.525
+ $X2=3.005 $Y2=1.935
r119 22 36 6.09054 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.535 $Y=2.02
+ $X2=0.32 $Y2=2.02
r120 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.92 $Y=2.02
+ $X2=3.005 $Y2=1.935
r121 21 22 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=2.92 $Y=2.02
+ $X2=0.535 $Y2=2.02
r122 20 35 8.32692 $w=4.21e-07 $l=2.1609e-07 $layer=LI1_cond $X=0.202 $Y=1.795
+ $X2=0.32 $Y2=1.96
r123 20 33 54.317 $w=1.93e-07 $l=9.55e-07 $layer=LI1_cond $X=0.202 $Y=1.795
+ $X2=0.202 $Y2=0.84
r124 16 47 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.09 $Y=0.995
+ $X2=4.09 $Y2=1.202
r125 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.09 $Y=0.995
+ $X2=4.09 $Y2=0.56
r126 13 46 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.065 $Y=1.41
+ $X2=4.065 $Y2=1.202
r127 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.065 $Y=1.41
+ $X2=4.065 $Y2=1.985
r128 10 45 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.62 $Y=0.995
+ $X2=3.62 $Y2=1.202
r129 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.62 $Y=0.995
+ $X2=3.62 $Y2=0.56
r130 7 44 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.595 $Y=1.41
+ $X2=3.595 $Y2=1.202
r131 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.595 $Y=1.41
+ $X2=3.595 $Y2=1.985
r132 2 38 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.485 $X2=0.425 $Y2=2.3
r133 2 35 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.485 $X2=0.425 $Y2=1.96
r134 1 31 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.18
+ $Y=0.235 $X2=0.345 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_4%A2 1 3 4 6 7 9 10 12 14 15 16 17 19 28 31
+ 36
c81 31 0 1.1034e-19 $X=5.69 $Y=1.445
c82 14 0 1.54054e-19 $X=4.677 $Y=1.595
r83 31 36 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=1.68
+ $X2=5.745 $Y2=1.595
r84 31 36 3.75797 $w=2.28e-07 $l=7.5e-08 $layer=LI1_cond $X=5.745 $Y=1.52
+ $X2=5.745 $Y2=1.595
r85 30 31 11.5244 $w=2.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.745 $Y=1.29
+ $X2=5.745 $Y2=1.52
r86 25 28 7.26257 $w=2.63e-07 $l=1.67e-07 $layer=LI1_cond $X=4.51 $Y=1.142
+ $X2=4.677 $Y2=1.142
r87 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.51
+ $Y=1.16 $X2=4.51 $Y2=1.16
r88 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.98
+ $Y=1.16 $X2=5.98 $Y2=1.16
r89 17 30 6.81752 $w=2.35e-07 $l=1.65813e-07 $layer=LI1_cond $X=5.86 $Y=1.172
+ $X2=5.745 $Y2=1.29
r90 17 19 3.18761 $w=2.33e-07 $l=6.5e-08 $layer=LI1_cond $X=5.86 $Y=1.172
+ $X2=5.925 $Y2=1.172
r91 15 31 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.63 $Y=1.68
+ $X2=5.745 $Y2=1.68
r92 15 16 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.63 $Y=1.68
+ $X2=4.79 $Y2=1.68
r93 14 16 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=4.677 $Y=1.595
+ $X2=4.79 $Y2=1.68
r94 13 28 1.71951 $w=2.25e-07 $l=1.33e-07 $layer=LI1_cond $X=4.677 $Y=1.275
+ $X2=4.677 $Y2=1.142
r95 13 14 16.3903 $w=2.23e-07 $l=3.2e-07 $layer=LI1_cond $X=4.677 $Y=1.275
+ $X2=4.677 $Y2=1.595
r96 10 22 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=5.945 $Y=1.41
+ $X2=6.005 $Y2=1.16
r97 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.945 $Y=1.41
+ $X2=5.945 $Y2=1.985
r98 7 22 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=5.92 $Y=0.995
+ $X2=6.005 $Y2=1.16
r99 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.92 $Y=0.995 $X2=5.92
+ $Y2=0.56
r100 4 26 38.578 $w=2.95e-07 $l=1.94808e-07 $layer=POLY_cond $X=4.6 $Y=0.995
+ $X2=4.535 $Y2=1.16
r101 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.6 $Y=0.995 $X2=4.6
+ $Y2=0.56
r102 1 26 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=4.535 $Y=1.41
+ $X2=4.535 $Y2=1.16
r103 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.535 $Y=1.41
+ $X2=4.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_4%A1 1 3 4 6 7 9 10 12 13 20
r47 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=1.202
+ $X2=5.5 $Y2=1.202
r48 18 20 33.6132 $w=3.8e-07 $l=2.65e-07 $layer=POLY_cond $X=5.21 $Y=1.202
+ $X2=5.475 $Y2=1.202
r49 16 18 26.0026 $w=3.8e-07 $l=2.05e-07 $layer=POLY_cond $X=5.005 $Y=1.202
+ $X2=5.21 $Y2=1.202
r50 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.98 $Y=1.202
+ $X2=5.005 $Y2=1.202
r51 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.21
+ $Y=1.16 $X2=5.21 $Y2=1.16
r52 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.5 $Y=0.995
+ $X2=5.5 $Y2=1.202
r53 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.5 $Y=0.995 $X2=5.5
+ $Y2=0.56
r54 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.202
r55 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.985
r56 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.005 $Y=1.41
+ $X2=5.005 $Y2=1.202
r57 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.005 $Y=1.41
+ $X2=5.005 $Y2=1.985
r58 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.98 $Y=0.995
+ $X2=4.98 $Y2=1.202
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.98 $Y=0.995 $X2=4.98
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_4%VPWR 1 2 3 4 5 19 22 26 29 32 41 48 55 56
+ 59 62 66 73
r99 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r100 73 76 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.685 $Y=2.36
+ $X2=5.685 $Y2=2.72
r101 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r102 66 69 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.745 $Y=2.36
+ $X2=4.745 $Y2=2.72
r103 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r104 59 62 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.88 $Y=2.36
+ $X2=0.88 $Y2=2.72
r105 56 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r106 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r107 53 76 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.875 $Y=2.72
+ $X2=5.685 $Y2=2.72
r108 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.875 $Y=2.72
+ $X2=6.21 $Y2=2.72
r109 52 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r110 52 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r111 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r112 49 69 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=4.745 $Y2=2.72
r113 49 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=5.29 $Y2=2.72
r114 48 76 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.495 $Y=2.72
+ $X2=5.685 $Y2=2.72
r115 48 51 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.495 $Y=2.72
+ $X2=5.29 $Y2=2.72
r116 47 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r117 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r118 44 47 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r119 43 46 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r120 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r121 41 69 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.555 $Y=2.72
+ $X2=4.745 $Y2=2.72
r122 41 46 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.555 $Y=2.72
+ $X2=4.37 $Y2=2.72
r123 40 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r124 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r125 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r126 37 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r127 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r128 34 62 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.07 $Y=2.72
+ $X2=0.88 $Y2=2.72
r129 34 36 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r130 32 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r131 29 39 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.605 $Y=2.72
+ $X2=2.53 $Y2=2.72
r132 29 43 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.797 $Y=2.72
+ $X2=2.99 $Y2=2.72
r133 26 29 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=2.797 $Y=2.36
+ $X2=2.797 $Y2=2.72
r134 23 39 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.03 $Y=2.72 $X2=2.53
+ $Y2=2.72
r135 22 36 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.65 $Y=2.72 $X2=1.61
+ $Y2=2.72
r136 21 23 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.84 $Y=2.72
+ $X2=2.03 $Y2=2.72
r137 21 22 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.84 $Y=2.72
+ $X2=1.65 $Y2=2.72
r138 19 21 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.84 $Y=2.36
+ $X2=1.84 $Y2=2.72
r139 5 73 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=2.36
r140 4 66 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=1.485 $X2=4.77 $Y2=2.36
r141 3 26 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=1.485 $X2=2.82 $Y2=2.36
r142 2 19 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=1.485 $X2=1.865 $Y2=2.36
r143 1 59 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=1.485 $X2=0.905 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_4%X 1 2 3 4 15 19 21 24 27 30
c47 27 0 6.40318e-20 $X=1.295 $Y=1.595
r48 27 30 1.58663 $w=4.88e-07 $l=6.5e-08 $layer=LI1_cond $X=1.295 $Y=1.595
+ $X2=1.295 $Y2=1.53
r49 24 27 2.35588 $w=4.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=1.68
+ $X2=1.295 $Y2=1.595
r50 24 30 0.244098 $w=4.88e-07 $l=1e-08 $layer=LI1_cond $X=1.295 $Y=1.52
+ $X2=1.295 $Y2=1.53
r51 21 24 17.9412 $w=4.88e-07 $l=7.35e-07 $layer=LI1_cond $X=1.295 $Y=0.785
+ $X2=1.295 $Y2=1.52
r52 21 23 2.35588 $w=4.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.785
+ $X2=1.295 $Y2=0.7
r53 17 24 6.79047 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=1.54 $Y=1.68
+ $X2=1.295 $Y2=1.68
r54 17 19 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.54 $Y=1.68
+ $X2=2.345 $Y2=1.68
r55 13 23 6.79047 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=1.54 $Y=0.7
+ $X2=1.295 $Y2=0.7
r56 13 15 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.54 $Y=0.7
+ $X2=2.345 $Y2=0.7
r57 4 19 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.195
+ $Y=1.485 $X2=2.345 $Y2=1.68
r58 3 24 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.485 $X2=1.385 $Y2=1.68
r59 2 15 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.235 $X2=2.345 $Y2=0.7
r60 1 23 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.235 $X2=1.385 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_4%A_647_297# 1 2 3 4 15 17 18 21 23 29 32
r55 32 33 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=4.295 $Y=2.02
+ $X2=4.295 $Y2=2.295
r56 27 29 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=6.217 $Y=1.935
+ $X2=6.217 $Y2=1.63
r57 24 32 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.385 $Y=2.02 $X2=4.295
+ $Y2=2.02
r58 24 26 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.385 $Y=2.02
+ $X2=5.24 $Y2=2.02
r59 23 27 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=6.09 $Y=2.02
+ $X2=6.217 $Y2=1.935
r60 23 26 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=6.09 $Y=2.02
+ $X2=5.24 $Y2=2.02
r61 19 32 5.23737 $w=1.78e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=1.935
+ $X2=4.295 $Y2=2.02
r62 19 21 20.0253 $w=1.78e-07 $l=3.25e-07 $layer=LI1_cond $X=4.295 $Y=1.935
+ $X2=4.295 $Y2=1.61
r63 17 33 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.205 $Y=2.295
+ $X2=4.295 $Y2=2.295
r64 17 18 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.205 $Y=2.295
+ $X2=3.445 $Y2=2.295
r65 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.36 $Y=2.21
+ $X2=3.445 $Y2=2.295
r66 13 15 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.36 $Y=2.21
+ $X2=3.36 $Y2=1.86
r67 4 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=1.63
r68 3 26 600 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=1 $X=5.095
+ $Y=1.485 $X2=5.24 $Y2=2.02
r69 2 32 600 $w=1.7e-07 $l=6.38396e-07 $layer=licon1_PDIFF $count=1 $X=4.155
+ $Y=1.485 $X2=4.3 $Y2=2.055
r70 2 21 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.155
+ $Y=1.485 $X2=4.3 $Y2=1.61
r71 1 15 300 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=2 $X=3.235
+ $Y=1.485 $X2=3.36 $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_4%VGND 1 2 3 4 5 20 22 24 26 27 33 43 48 58
+ 66 69 71 75
r85 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r86 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r87 68 69 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.34 $Y=0.18
+ $X2=3.505 $Y2=0.18
r88 64 68 7.89863 $w=5.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.99 $Y=0.18
+ $X2=3.34 $Y2=0.18
r89 64 66 11.7354 $w=5.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.99 $Y=0.18
+ $X2=2.735 $Y2=0.18
r90 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r91 58 61 10.6379 $w=3.88e-07 $l=3.6e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.875
+ $Y2=0.36
r92 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r93 55 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r94 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r95 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r96 52 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r97 51 54 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r98 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r99 49 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.505 $Y=0 $X2=4.34
+ $Y2=0
r100 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.505 $Y=0
+ $X2=4.83 $Y2=0
r101 48 74 4.31451 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=6.065 $Y=0
+ $X2=6.252 $Y2=0
r102 48 54 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.065 $Y=0
+ $X2=5.75 $Y2=0
r103 47 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r104 47 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r105 46 69 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.91 $Y=0
+ $X2=3.505 $Y2=0
r106 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r107 43 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.175 $Y=0 $X2=4.34
+ $Y2=0
r108 43 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.175 $Y=0
+ $X2=3.91 $Y2=0
r109 42 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r110 41 66 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.53 $Y=0
+ $X2=2.735 $Y2=0
r111 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r112 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r113 38 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r114 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r115 35 58 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=0.875
+ $Y2=0
r116 35 37 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=1.61
+ $Y2=0
r117 33 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r118 29 41 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.53
+ $Y2=0
r119 27 37 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.61
+ $Y2=0
r120 26 31 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=1.84
+ $Y2=0.36
r121 26 29 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=2.03
+ $Y2=0
r122 26 27 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=1.65
+ $Y2=0
r123 22 74 3.04554 $w=2.8e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.205 $Y=0.085
+ $X2=6.252 $Y2=0
r124 22 24 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=6.205 $Y=0.085
+ $X2=6.205 $Y2=0.38
r125 18 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.085
+ $X2=4.34 $Y2=0
r126 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.34 $Y=0.085
+ $X2=4.34 $Y2=0.36
r127 5 24 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=5.995
+ $Y=0.235 $X2=6.18 $Y2=0.38
r128 4 20 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=4.165
+ $Y=0.235 $X2=4.34 $Y2=0.36
r129 3 68 91 $w=1.7e-07 $l=7.64951e-07 $layer=licon1_NDIFF $count=2 $X=2.635
+ $Y=0.235 $X2=3.34 $Y2=0.36
r130 2 31 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.675
+ $Y=0.235 $X2=1.865 $Y2=0.36
r131 1 61 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.765
+ $Y=0.235 $X2=0.905 $Y2=0.36
.ends

