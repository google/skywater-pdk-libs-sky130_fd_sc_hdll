* File: sky130_fd_sc_hdll__buf_1.pex.spice
* Created: Wed Sep  2 08:24:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUF_1%A 2 3 5 8 10 13
c33 13 0 2.95098e-19 $X=0.46 $Y=1.16
c34 8 0 8.7047e-20 $X=0.52 $Y=0.495
r35 13 16 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.46 $Y=1.16
+ $X2=0.46 $Y2=1.325
r36 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.46 $Y=1.16
+ $X2=0.46 $Y2=0.995
r37 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.46
+ $Y=1.16 $X2=0.46 $Y2=1.16
r38 8 15 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.52 $Y=0.495 $X2=0.52
+ $Y2=0.995
r39 3 5 125.856 $w=1.8e-07 $l=4.7e-07 $layer=POLY_cond $X=0.495 $Y=1.62
+ $X2=0.495 $Y2=2.09
r40 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.52 $X2=0.495
+ $Y2=1.62
r41 2 16 64.6575 $w=2e-07 $l=1.95e-07 $layer=POLY_cond $X=0.495 $Y=1.52
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_1%A_27_47# 1 2 7 9 12 16 20 22 23 24 25 29 31
+ 33
c60 25 0 1.45394e-19 $X=0.345 $Y=1.62
c61 23 0 1.49704e-19 $X=0.345 $Y=0.72
r62 31 34 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.877 $Y=1.225
+ $X2=0.877 $Y2=1.39
r63 31 33 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.877 $Y=1.225
+ $X2=0.877 $Y2=1.06
r64 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.225 $X2=0.95 $Y2=1.225
r65 29 34 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.805 $Y=1.535
+ $X2=0.805 $Y2=1.39
r66 26 33 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.805 $Y=0.805
+ $X2=0.805 $Y2=1.06
r67 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=1.62
+ $X2=0.805 $Y2=1.535
r68 24 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.72 $Y=1.62
+ $X2=0.345 $Y2=1.62
r69 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=0.72
+ $X2=0.805 $Y2=0.805
r70 22 23 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.72 $Y=0.72
+ $X2=0.345 $Y2=0.72
r71 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r72 18 20 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.445
r73 14 25 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.255 $Y=1.705
+ $X2=0.345 $Y2=1.62
r74 14 16 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.255 $Y=1.705
+ $X2=0.255 $Y2=1.96
r75 10 32 39.8325 $w=2.41e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.01 $Y=1.06
+ $X2=0.95 $Y2=1.225
r76 10 12 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.01 $Y=1.06
+ $X2=1.01 $Y2=0.495
r77 7 32 82.1933 $w=2.41e-07 $l=4.12129e-07 $layer=POLY_cond $X=0.985 $Y=1.62
+ $X2=0.95 $Y2=1.225
r78 7 9 125.856 $w=1.8e-07 $l=4.7e-07 $layer=POLY_cond $X=0.985 $Y=1.62
+ $X2=0.985 $Y2=2.09
r79 2 16 300 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.695 $X2=0.26 $Y2=1.96
r80 1 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_1%VPWR 1 6 8 10 12 20 21 24
r22 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r23 21 25 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r24 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r25 18 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.71 $Y2=2.72
r26 18 20 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r27 12 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.71 $Y2=2.72
r28 10 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r29 8 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.525 $Y2=2.72
r30 8 10 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r31 4 24 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.635 $X2=0.71
+ $Y2=2.72
r32 4 6 21.0243 $w=3.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.71 $Y=2.635
+ $X2=0.71 $Y2=1.96
r33 1 6 300 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.695 $X2=0.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_1%X 1 2 9 10 11 12 13 33
c25 33 0 8.7047e-20 $X=1.23 $Y=0.76
r26 12 13 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.23 $Y=1.87
+ $X2=1.23 $Y2=2.21
r27 11 33 7.19178 $w=4.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=0.595
+ $X2=1.23 $Y2=0.76
r28 10 33 49.2929 $w=1.78e-07 $l=8e-07 $layer=LI1_cond $X=1.305 $Y=1.56
+ $X2=1.305 $Y2=0.76
r29 9 12 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.23 $Y=1.725
+ $X2=1.23 $Y2=1.87
r30 9 10 8.12648 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=1.725
+ $X2=1.23 $Y2=1.56
r31 2 12 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.695 $X2=1.22 $Y2=1.895
r32 1 11 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_1%VGND 1 6 8 10 12 17 21 22 25
r23 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r24 22 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r25 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r26 19 25 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.71
+ $Y2=0
r27 19 21 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.61
+ $Y2=0
r28 12 25 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.71
+ $Y2=0
r29 10 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r30 10 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r31 8 12 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.525
+ $Y2=0
r32 8 17 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.23
+ $Y2=0
r33 4 25 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r34 4 6 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.38
r35 1 6 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

