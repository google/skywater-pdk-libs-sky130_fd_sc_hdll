* File: sky130_fd_sc_hdll__ebufn_2.pxi.spice
* Created: Thu Aug 27 19:07:01 2020
* 
x_PM_SKY130_FD_SC_HDLL__EBUFN_2%A N_A_M1010_g N_A_c_75_n N_A_c_76_n N_A_M1000_g
+ A A N_A_c_74_n PM_SKY130_FD_SC_HDLL__EBUFN_2%A
x_PM_SKY130_FD_SC_HDLL__EBUFN_2%TE_B N_TE_B_M1002_g N_TE_B_c_111_n
+ N_TE_B_c_112_n N_TE_B_M1006_g N_TE_B_c_113_n N_TE_B_c_114_n N_TE_B_M1007_g
+ N_TE_B_c_115_n N_TE_B_c_116_n N_TE_B_M1008_g N_TE_B_c_117_n TE_B
+ N_TE_B_c_110_n PM_SKY130_FD_SC_HDLL__EBUFN_2%TE_B
x_PM_SKY130_FD_SC_HDLL__EBUFN_2%A_224_47# N_A_224_47#_M1002_d
+ N_A_224_47#_M1006_d N_A_224_47#_c_177_n N_A_224_47#_M1001_g
+ N_A_224_47#_c_178_n N_A_224_47#_c_179_n N_A_224_47#_M1004_g
+ N_A_224_47#_c_180_n N_A_224_47#_c_187_n N_A_224_47#_c_181_n
+ N_A_224_47#_c_182_n N_A_224_47#_c_183_n N_A_224_47#_c_189_n
+ N_A_224_47#_c_184_n N_A_224_47#_c_185_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_2%A_224_47#
x_PM_SKY130_FD_SC_HDLL__EBUFN_2%A_27_47# N_A_27_47#_M1010_s N_A_27_47#_M1000_s
+ N_A_27_47#_M1005_g N_A_27_47#_c_265_n N_A_27_47#_M1003_g N_A_27_47#_c_266_n
+ N_A_27_47#_M1009_g N_A_27_47#_M1011_g N_A_27_47#_c_260_n N_A_27_47#_c_281_n
+ N_A_27_47#_c_261_n N_A_27_47#_c_262_n N_A_27_47#_c_263_n N_A_27_47#_c_264_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EBUFN_2%VPWR N_VPWR_M1000_d N_VPWR_M1007_s
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n VPWR N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_335_n N_VPWR_c_342_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_2%VPWR
x_PM_SKY130_FD_SC_HDLL__EBUFN_2%A_340_309# N_A_340_309#_M1007_d
+ N_A_340_309#_M1008_d N_A_340_309#_M1009_d N_A_340_309#_c_398_n
+ N_A_340_309#_c_389_n N_A_340_309#_c_390_n N_A_340_309#_c_391_n
+ N_A_340_309#_c_393_n N_A_340_309#_c_396_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_2%A_340_309#
x_PM_SKY130_FD_SC_HDLL__EBUFN_2%Z N_Z_M1005_s N_Z_M1003_s N_Z_c_449_n
+ N_Z_c_437_n Z Z Z Z Z Z Z N_Z_c_440_n Z Z Z N_Z_c_436_n N_Z_c_441_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_2%Z
x_PM_SKY130_FD_SC_HDLL__EBUFN_2%VGND N_VGND_M1010_d N_VGND_M1001_d
+ N_VGND_c_493_n N_VGND_c_494_n VGND N_VGND_c_495_n N_VGND_c_496_n
+ N_VGND_c_497_n N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_2%VGND
x_PM_SKY130_FD_SC_HDLL__EBUFN_2%A_412_47# N_A_412_47#_M1001_s
+ N_A_412_47#_M1004_s N_A_412_47#_M1011_d N_A_412_47#_c_550_n
+ N_A_412_47#_c_556_n N_A_412_47#_c_551_n N_A_412_47#_c_562_n
+ N_A_412_47#_c_563_n N_A_412_47#_c_552_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_2%A_412_47#
cc_1 VNB N_A_M1010_g 0.0331912f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A 0.00515246f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_3 VNB N_A_c_74_n 0.0288146f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_4 VNB N_TE_B_M1002_g 0.0369037f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_5 VNB TE_B 0.00797222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_TE_B_c_110_n 0.0273119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_224_47#_c_177_n 0.017408f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.77
cc_8 VNB N_A_224_47#_c_178_n 0.0385858f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_9 VNB N_A_224_47#_c_179_n 0.00859481f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_10 VNB N_A_224_47#_c_180_n 0.0125944f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_11 VNB N_A_224_47#_c_181_n 0.0130355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_224_47#_c_182_n 0.0013647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_224_47#_c_183_n 0.0228928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_224_47#_c_184_n 0.00280572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_224_47#_c_185_n 0.0153829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_M1005_g 0.0200702f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.165
cc_17 VNB N_A_27_47#_M1011_g 0.0219261f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.85
cc_18 VNB N_A_27_47#_c_260_n 0.0124311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_261_n 0.00175392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_262_n 0.0152409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_263_n 0.0438172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_264_n 0.0424277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_335_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB Z 0.0225392f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=0.995
cc_25 VNB N_Z_c_436_n 0.0109904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_493_n 0.00307453f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.165
cc_27 VNB N_VGND_c_494_n 4.89699e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_495_n 0.0151734f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=0.995
cc_29 VNB N_VGND_c_496_n 0.0385018f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_30 VNB N_VGND_c_497_n 0.0431128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_498_n 0.252128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_499_n 0.00613341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_500_n 0.00502768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_412_47#_c_550_n 0.00499888f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_35 VNB N_A_412_47#_c_551_n 0.00268163f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.16
cc_36 VNB N_A_412_47#_c_552_n 0.00871563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VPB N_A_c_75_n 0.0205511f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_38 VPB N_A_c_76_n 0.0268833f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_39 VPB A 0.00510322f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.765
cc_40 VPB N_A_c_74_n 0.00541359f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_41 VPB N_TE_B_c_111_n 0.0129566f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_42 VPB N_TE_B_c_112_n 0.027196f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_43 VPB N_TE_B_c_113_n 0.0465319f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.765
cc_44 VPB N_TE_B_c_114_n 0.018413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_TE_B_c_115_n 0.0283251f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_46 VPB N_TE_B_c_116_n 0.0191144f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=0.995
cc_47 VPB N_TE_B_c_117_n 0.00735165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_TE_B_c_110_n 0.0110197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_224_47#_c_178_n 0.00914443f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.765
cc_50 VPB N_A_224_47#_c_187_n 0.0107265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_224_47#_c_182_n 7.0588e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_224_47#_c_189_n 0.0130404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_265_n 0.0200905f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_54 VPB N_A_27_47#_c_266_n 0.0191741f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.16
cc_55 VPB N_A_27_47#_c_263_n 0.0159147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_264_n 0.0522423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_336_n 0.00469661f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_58 VPB N_VPWR_c_337_n 0.00556536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_338_n 0.0267715f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_60 VPB N_VPWR_c_339_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_340_n 0.0515168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_335_n 0.0568819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_342_n 0.00663993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_340_309#_c_389_n 0.00131456f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_65 VPB N_A_340_309#_c_390_n 0.00759475f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_66 VPB N_A_340_309#_c_391_n 0.0194249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_Z_c_437_n 0.00195862f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_68 VPB Z 0.00731007f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=0.995
cc_69 VPB Z 0.00953505f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=0.85
cc_70 VPB N_Z_c_440_n 0.00623256f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_Z_c_441_n 0.00143709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 N_A_M1010_g N_TE_B_M1002_g 0.0184879f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_73 A N_TE_B_M1002_g 0.00159023f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_74 N_A_c_74_n N_TE_B_M1002_g 0.0185122f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_c_76_n N_TE_B_c_111_n 0.00653324f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_76 N_A_c_76_n N_TE_B_c_112_n 0.0148662f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_77 N_A_M1010_g TE_B 5.40201e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_78 A TE_B 0.0402744f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_79 N_A_c_74_n TE_B 7.69775e-19 $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_c_75_n N_TE_B_c_110_n 0.00653324f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_81 A N_TE_B_c_110_n 0.00632969f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_82 A N_A_224_47#_c_189_n 0.00993953f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_83 A N_A_27_47#_c_260_n 0.00266482f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_84 N_A_c_74_n N_A_27_47#_c_260_n 0.00266134f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_85 A N_A_27_47#_c_262_n 0.0164018f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_86 N_A_c_74_n N_A_27_47#_c_262_n 0.0116614f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_M1010_g N_A_27_47#_c_264_n 0.0300471f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_c_76_n N_A_27_47#_c_264_n 0.00953388f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_89 A N_A_27_47#_c_264_n 0.0671602f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_90 N_A_c_76_n N_VPWR_c_336_n 0.0271995f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_91 A N_VPWR_c_336_n 0.0201565f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_92 N_A_c_74_n N_VPWR_c_336_n 4.5672e-19 $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_c_76_n N_VPWR_c_339_n 0.00427505f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_94 N_A_c_76_n N_VPWR_c_335_n 0.00835414f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_95 N_A_M1010_g N_VGND_c_493_n 0.0115284f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_96 A N_VGND_c_493_n 0.0196224f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_97 N_A_c_74_n N_VGND_c_493_n 7.77e-19 $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_M1010_g N_VGND_c_495_n 0.0046653f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_M1010_g N_VGND_c_498_n 0.00895857f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_100 A N_VGND_c_498_n 0.00103459f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_101 N_TE_B_c_115_n N_A_224_47#_c_178_n 3.91667e-19 $X=2.44 $Y=1.395 $X2=0
+ $Y2=0
cc_102 N_TE_B_c_115_n N_A_224_47#_c_179_n 0.0136463f $X=2.44 $Y=1.395 $X2=0
+ $Y2=0
cc_103 N_TE_B_M1002_g N_A_224_47#_c_180_n 0.00518275f $X=1.045 $Y=0.445 $X2=0
+ $Y2=0
cc_104 TE_B N_A_224_47#_c_180_n 0.0157345f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_105 N_TE_B_c_110_n N_A_224_47#_c_180_n 6.59347e-19 $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_106 N_TE_B_c_112_n N_A_224_47#_c_187_n 0.010345f $X=1.07 $Y=1.77 $X2=0 $Y2=0
cc_107 N_TE_B_c_114_n N_A_224_47#_c_187_n 0.0059554f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_108 N_TE_B_c_110_n N_A_224_47#_c_187_n 8.70198e-19 $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_109 N_TE_B_M1002_g N_A_224_47#_c_181_n 0.00530078f $X=1.045 $Y=0.445 $X2=0
+ $Y2=0
cc_110 TE_B N_A_224_47#_c_181_n 0.0163628f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_111 N_TE_B_c_110_n N_A_224_47#_c_181_n 2.12603e-19 $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_112 N_TE_B_c_113_n N_A_224_47#_c_182_n 0.0216386f $X=1.97 $Y=1.395 $X2=0
+ $Y2=0
cc_113 N_TE_B_c_110_n N_A_224_47#_c_182_n 0.00161087f $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_114 N_TE_B_c_113_n N_A_224_47#_c_183_n 0.0194291f $X=1.97 $Y=1.395 $X2=0
+ $Y2=0
cc_115 N_TE_B_c_111_n N_A_224_47#_c_189_n 0.0101387f $X=1.07 $Y=1.67 $X2=0 $Y2=0
cc_116 N_TE_B_c_113_n N_A_224_47#_c_189_n 0.016278f $X=1.97 $Y=1.395 $X2=0 $Y2=0
cc_117 N_TE_B_c_114_n N_A_224_47#_c_189_n 0.00613026f $X=2.06 $Y=1.47 $X2=0
+ $Y2=0
cc_118 TE_B N_A_224_47#_c_189_n 0.00561075f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_119 N_TE_B_c_110_n N_A_224_47#_c_189_n 0.00245935f $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_120 N_TE_B_c_113_n N_A_224_47#_c_184_n 4.76658e-19 $X=1.97 $Y=1.395 $X2=0
+ $Y2=0
cc_121 TE_B N_A_224_47#_c_184_n 0.0135202f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_122 N_TE_B_c_110_n N_A_224_47#_c_184_n 0.00459165f $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_123 N_TE_B_c_113_n N_A_27_47#_c_262_n 0.00566409f $X=1.97 $Y=1.395 $X2=0
+ $Y2=0
cc_124 TE_B N_A_27_47#_c_262_n 0.0298487f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_125 N_TE_B_c_110_n N_A_27_47#_c_262_n 0.00229642f $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_126 N_TE_B_c_112_n N_VPWR_c_336_n 0.0140613f $X=1.07 $Y=1.77 $X2=0 $Y2=0
cc_127 TE_B N_VPWR_c_336_n 0.00105855f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_128 N_TE_B_c_114_n N_VPWR_c_337_n 0.010738f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_129 N_TE_B_c_116_n N_VPWR_c_337_n 0.0081454f $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_130 N_TE_B_c_112_n N_VPWR_c_338_n 0.00622633f $X=1.07 $Y=1.77 $X2=0 $Y2=0
cc_131 N_TE_B_c_114_n N_VPWR_c_338_n 0.00309549f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_132 N_TE_B_c_116_n N_VPWR_c_340_n 0.00450253f $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_133 N_TE_B_c_112_n N_VPWR_c_335_n 0.0118107f $X=1.07 $Y=1.77 $X2=0 $Y2=0
cc_134 N_TE_B_c_114_n N_VPWR_c_335_n 0.00495823f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_135 N_TE_B_c_116_n N_VPWR_c_335_n 0.0064627f $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_136 N_TE_B_c_113_n N_A_340_309#_c_389_n 0.00163695f $X=1.97 $Y=1.395 $X2=0
+ $Y2=0
cc_137 N_TE_B_c_114_n N_A_340_309#_c_393_n 0.014254f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_138 N_TE_B_c_115_n N_A_340_309#_c_393_n 4.11517e-19 $X=2.44 $Y=1.395 $X2=0
+ $Y2=0
cc_139 N_TE_B_c_116_n N_A_340_309#_c_393_n 0.015268f $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_140 N_TE_B_c_116_n N_A_340_309#_c_396_n 0.0126492f $X=2.53 $Y=1.47 $X2=0
+ $Y2=0
cc_141 N_TE_B_c_114_n N_Z_c_440_n 0.012f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_142 N_TE_B_c_115_n N_Z_c_440_n 0.00786091f $X=2.44 $Y=1.395 $X2=0 $Y2=0
cc_143 N_TE_B_c_116_n N_Z_c_440_n 0.018198f $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_144 N_TE_B_c_117_n N_Z_c_440_n 0.00206935f $X=2.06 $Y=1.395 $X2=0 $Y2=0
cc_145 N_TE_B_M1002_g N_VGND_c_493_n 0.0066614f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_146 N_TE_B_M1002_g N_VGND_c_496_n 0.00509549f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_147 N_TE_B_M1002_g N_VGND_c_498_n 0.00756462f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_148 TE_B N_VGND_c_498_n 0.00470396f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_149 N_A_224_47#_c_178_n N_A_27_47#_M1005_g 0.0177818f $X=2.84 $Y=1.035 $X2=0
+ $Y2=0
cc_150 N_A_224_47#_c_185_n N_A_27_47#_M1005_g 0.0165303f $X=2.987 $Y=0.96 $X2=0
+ $Y2=0
cc_151 N_A_224_47#_c_183_n N_A_27_47#_c_281_n 6.39895e-19 $X=3 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_224_47#_c_178_n N_A_27_47#_c_261_n 3.49161e-19 $X=2.84 $Y=1.035 $X2=0
+ $Y2=0
cc_153 N_A_224_47#_c_183_n N_A_27_47#_c_261_n 0.0114076f $X=3 $Y=1.16 $X2=0
+ $Y2=0
cc_154 N_A_224_47#_c_180_n N_A_27_47#_c_262_n 0.00958493f $X=1.55 $Y=0.425 $X2=0
+ $Y2=0
cc_155 N_A_224_47#_c_183_n N_A_27_47#_c_262_n 0.0625906f $X=3 $Y=1.16 $X2=0
+ $Y2=0
cc_156 N_A_224_47#_c_189_n N_A_27_47#_c_262_n 0.0127794f $X=1.682 $Y=1.605 $X2=0
+ $Y2=0
cc_157 N_A_224_47#_c_184_n N_A_27_47#_c_262_n 0.024679f $X=1.69 $Y=1.15 $X2=0
+ $Y2=0
cc_158 N_A_224_47#_c_183_n N_A_27_47#_c_263_n 0.00179139f $X=3 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A_224_47#_c_187_n N_VPWR_c_336_n 0.0402328f $X=1.305 $Y=2.22 $X2=0
+ $Y2=0
cc_160 N_A_224_47#_c_187_n N_VPWR_c_338_n 0.0204048f $X=1.305 $Y=2.22 $X2=0
+ $Y2=0
cc_161 N_A_224_47#_M1006_d N_VPWR_c_335_n 0.00430086f $X=1.16 $Y=1.845 $X2=0
+ $Y2=0
cc_162 N_A_224_47#_c_187_n N_VPWR_c_335_n 0.0110999f $X=1.305 $Y=2.22 $X2=0
+ $Y2=0
cc_163 N_A_224_47#_c_189_n N_A_340_309#_M1007_d 0.00378908f $X=1.682 $Y=1.605
+ $X2=-0.19 $Y2=-0.24
cc_164 N_A_224_47#_c_187_n N_A_340_309#_c_398_n 0.0259829f $X=1.305 $Y=2.22
+ $X2=0 $Y2=0
cc_165 N_A_224_47#_c_187_n N_A_340_309#_c_389_n 0.0134641f $X=1.305 $Y=2.22
+ $X2=0 $Y2=0
cc_166 N_A_224_47#_c_183_n N_A_340_309#_c_389_n 0.00244188f $X=3 $Y=1.16 $X2=0
+ $Y2=0
cc_167 N_A_224_47#_c_189_n N_A_340_309#_c_389_n 0.00958694f $X=1.682 $Y=1.605
+ $X2=0 $Y2=0
cc_168 N_A_224_47#_c_184_n N_A_340_309#_c_389_n 4.98355e-19 $X=1.69 $Y=1.15
+ $X2=0 $Y2=0
cc_169 N_A_224_47#_c_183_n N_A_340_309#_c_393_n 0.00130112f $X=3 $Y=1.16 $X2=0
+ $Y2=0
cc_170 N_A_224_47#_c_178_n N_Z_c_440_n 0.00886593f $X=2.84 $Y=1.035 $X2=0 $Y2=0
cc_171 N_A_224_47#_c_183_n N_Z_c_440_n 0.0873067f $X=3 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_224_47#_c_189_n N_Z_c_440_n 0.0275334f $X=1.682 $Y=1.605 $X2=0 $Y2=0
cc_173 N_A_224_47#_c_180_n N_VGND_c_493_n 0.0281689f $X=1.55 $Y=0.425 $X2=0
+ $Y2=0
cc_174 N_A_224_47#_c_177_n N_VGND_c_494_n 0.0115396f $X=2.495 $Y=0.96 $X2=0
+ $Y2=0
cc_175 N_A_224_47#_c_185_n N_VGND_c_494_n 0.0085985f $X=2.987 $Y=0.96 $X2=0
+ $Y2=0
cc_176 N_A_224_47#_c_177_n N_VGND_c_496_n 0.00199015f $X=2.495 $Y=0.96 $X2=0
+ $Y2=0
cc_177 N_A_224_47#_c_180_n N_VGND_c_496_n 0.050181f $X=1.55 $Y=0.425 $X2=0 $Y2=0
cc_178 N_A_224_47#_c_185_n N_VGND_c_497_n 0.00341689f $X=2.987 $Y=0.96 $X2=0
+ $Y2=0
cc_179 N_A_224_47#_M1002_d N_VGND_c_498_n 0.00251142f $X=1.12 $Y=0.235 $X2=0
+ $Y2=0
cc_180 N_A_224_47#_c_177_n N_VGND_c_498_n 0.00403341f $X=2.495 $Y=0.96 $X2=0
+ $Y2=0
cc_181 N_A_224_47#_c_180_n N_VGND_c_498_n 0.028699f $X=1.55 $Y=0.425 $X2=0 $Y2=0
cc_182 N_A_224_47#_c_185_n N_VGND_c_498_n 0.00442061f $X=2.987 $Y=0.96 $X2=0
+ $Y2=0
cc_183 N_A_224_47#_c_177_n N_A_412_47#_c_550_n 0.0116233f $X=2.495 $Y=0.96 $X2=0
+ $Y2=0
cc_184 N_A_224_47#_c_180_n N_A_412_47#_c_550_n 0.0300108f $X=1.55 $Y=0.425 $X2=0
+ $Y2=0
cc_185 N_A_224_47#_c_181_n N_A_412_47#_c_550_n 0.00484117f $X=1.69 $Y=1.025
+ $X2=0 $Y2=0
cc_186 N_A_224_47#_c_177_n N_A_412_47#_c_556_n 0.0140159f $X=2.495 $Y=0.96 $X2=0
+ $Y2=0
cc_187 N_A_224_47#_c_178_n N_A_412_47#_c_556_n 0.00534566f $X=2.84 $Y=1.035
+ $X2=0 $Y2=0
cc_188 N_A_224_47#_c_183_n N_A_412_47#_c_556_n 0.0539283f $X=3 $Y=1.16 $X2=0
+ $Y2=0
cc_189 N_A_224_47#_c_185_n N_A_412_47#_c_556_n 0.0132297f $X=2.987 $Y=0.96 $X2=0
+ $Y2=0
cc_190 N_A_224_47#_c_181_n N_A_412_47#_c_551_n 0.0174869f $X=1.69 $Y=1.025 $X2=0
+ $Y2=0
cc_191 N_A_224_47#_c_183_n N_A_412_47#_c_551_n 0.0248994f $X=3 $Y=1.16 $X2=0
+ $Y2=0
cc_192 N_A_224_47#_c_185_n N_A_412_47#_c_562_n 0.00469463f $X=2.987 $Y=0.96
+ $X2=0 $Y2=0
cc_193 N_A_224_47#_c_185_n N_A_412_47#_c_563_n 0.00191185f $X=2.987 $Y=0.96
+ $X2=0 $Y2=0
cc_194 N_A_27_47#_c_262_n N_VPWR_c_336_n 0.00747039f $X=3.57 $Y=1.145 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_264_n N_VPWR_c_336_n 0.0486687f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_264_n N_VPWR_c_339_n 0.0182101f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_265_n N_VPWR_c_340_n 0.00429453f $X=3.525 $Y=1.41 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_266_n N_VPWR_c_340_n 0.00429453f $X=3.995 $Y=1.41 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_M1000_s N_VPWR_c_335_n 0.00430086f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_265_n N_VPWR_c_335_n 0.00743756f $X=3.525 $Y=1.41 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_266_n N_VPWR_c_335_n 0.00706378f $X=3.995 $Y=1.41 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_264_n N_VPWR_c_335_n 0.00993603f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_265_n N_A_340_309#_c_390_n 0.0148808f $X=3.525 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_266_n N_A_340_309#_c_390_n 0.0102255f $X=3.995 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_265_n N_A_340_309#_c_396_n 0.0126492f $X=3.525 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_M1005_g N_Z_c_449_n 0.00305699f $X=3.5 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A_27_47#_M1011_g N_Z_c_449_n 0.0134839f $X=4.02 $Y=0.56 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_281_n N_Z_c_449_n 0.00260702f $X=3.765 $Y=1.145 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_261_n N_Z_c_449_n 0.0238517f $X=3.765 $Y=1.145 $X2=0 $Y2=0
cc_210 N_A_27_47#_c_263_n N_Z_c_449_n 0.00136944f $X=3.995 $Y=1.217 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_266_n N_Z_c_437_n 0.0108005f $X=3.995 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_263_n N_Z_c_437_n 3.64592e-19 $X=3.995 $Y=1.217 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_266_n Z 0.00126476f $X=3.995 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_27_47#_M1011_g Z 0.0186328f $X=4.02 $Y=0.56 $X2=0 $Y2=0
cc_215 N_A_27_47#_c_281_n Z 0.00151111f $X=3.765 $Y=1.145 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_261_n Z 0.0119436f $X=3.765 $Y=1.145 $X2=0 $Y2=0
cc_217 N_A_27_47#_c_265_n N_Z_c_440_n 0.0204197f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_261_n N_Z_c_440_n 0.00662079f $X=3.765 $Y=1.145 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_262_n N_Z_c_440_n 0.0203903f $X=3.57 $Y=1.145 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_263_n N_Z_c_440_n 5.12501e-19 $X=3.995 $Y=1.217 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_265_n N_Z_c_441_n 0.0124762f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_266_n N_Z_c_441_n 0.0192996f $X=3.995 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_281_n N_Z_c_441_n 0.00256437f $X=3.765 $Y=1.145 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_261_n N_Z_c_441_n 0.0268377f $X=3.765 $Y=1.145 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_263_n N_Z_c_441_n 0.0072138f $X=3.995 $Y=1.217 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_262_n N_VGND_c_493_n 0.00577688f $X=3.57 $Y=1.145 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_M1005_g N_VGND_c_494_n 0.00110864f $X=3.5 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_264_n N_VGND_c_495_n 0.015516f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A_27_47#_M1005_g N_VGND_c_497_n 0.00362032f $X=3.5 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A_27_47#_M1011_g N_VGND_c_497_n 0.00362032f $X=4.02 $Y=0.56 $X2=0 $Y2=0
cc_231 N_A_27_47#_M1010_s N_VGND_c_498_n 0.00388065f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1005_g N_VGND_c_498_n 0.00591554f $X=3.5 $Y=0.56 $X2=0 $Y2=0
cc_233 N_A_27_47#_M1011_g N_VGND_c_498_n 0.00652646f $X=4.02 $Y=0.56 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_264_n N_VGND_c_498_n 0.00981584f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_262_n N_A_412_47#_c_556_n 0.010201f $X=3.57 $Y=1.145 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_262_n N_A_412_47#_c_551_n 0.00217021f $X=3.57 $Y=1.145 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_M1005_g N_A_412_47#_c_552_n 0.0129646f $X=3.5 $Y=0.56 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_M1011_g N_A_412_47#_c_552_n 0.00890228f $X=4.02 $Y=0.56 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_261_n N_A_412_47#_c_552_n 0.00129798f $X=3.765 $Y=1.145
+ $X2=0 $Y2=0
cc_240 N_VPWR_c_335_n N_A_340_309#_M1007_d 0.00235746f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_241 N_VPWR_c_335_n N_A_340_309#_M1008_d 0.00682329f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_335_n N_A_340_309#_M1009_d 0.00233921f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_337_n N_A_340_309#_c_398_n 0.0144065f $X=2.295 $Y=2.36 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_338_n N_A_340_309#_c_398_n 0.0143637f $X=2.08 $Y=2.72 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_335_n N_A_340_309#_c_398_n 0.00795901f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_340_n N_A_340_309#_c_390_n 0.0183322f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_335_n N_A_340_309#_c_390_n 0.0100092f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_248 N_VPWR_M1007_s N_A_340_309#_c_393_n 0.00352612f $X=2.15 $Y=1.545 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_337_n N_A_340_309#_c_393_n 0.0195044f $X=2.295 $Y=2.36 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_338_n N_A_340_309#_c_393_n 0.00250551f $X=2.08 $Y=2.72 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_340_n N_A_340_309#_c_393_n 0.00336306f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_335_n N_A_340_309#_c_393_n 0.0115752f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_337_n N_A_340_309#_c_396_n 0.0129226f $X=2.295 $Y=2.36 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_340_n N_A_340_309#_c_396_n 0.0905296f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_335_n N_A_340_309#_c_396_n 0.0542792f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_335_n N_Z_M1003_s 0.00232895f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_257 N_VPWR_M1007_s N_Z_c_440_n 0.00191236f $X=2.15 $Y=1.545 $X2=0 $Y2=0
cc_258 N_A_340_309#_c_390_n N_Z_M1003_s 0.00352392f $X=4.165 $Y=2.38 $X2=0 $Y2=0
cc_259 N_A_340_309#_M1009_d N_Z_c_437_n 0.00115729f $X=4.085 $Y=1.485 $X2=0
+ $Y2=0
cc_260 N_A_340_309#_c_390_n N_Z_c_437_n 0.00252045f $X=4.165 $Y=2.38 $X2=0 $Y2=0
cc_261 N_A_340_309#_c_391_n N_Z_c_437_n 0.00518396f $X=4.25 $Y=1.96 $X2=0 $Y2=0
cc_262 N_A_340_309#_M1009_d Z 0.002457f $X=4.085 $Y=1.485 $X2=0 $Y2=0
cc_263 N_A_340_309#_c_391_n Z 0.0176452f $X=4.25 $Y=1.96 $X2=0 $Y2=0
cc_264 N_A_340_309#_M1008_d N_Z_c_440_n 0.0145194f $X=2.62 $Y=1.545 $X2=0 $Y2=0
cc_265 N_A_340_309#_c_390_n N_Z_c_440_n 0.00454431f $X=4.165 $Y=2.38 $X2=0 $Y2=0
cc_266 N_A_340_309#_c_393_n N_Z_c_440_n 0.095772f $X=2.68 $Y=2.2 $X2=0 $Y2=0
cc_267 N_A_340_309#_c_390_n N_Z_c_441_n 0.0210394f $X=4.165 $Y=2.38 $X2=0 $Y2=0
cc_268 N_A_340_309#_c_391_n N_Z_c_441_n 0.0255232f $X=4.25 $Y=1.96 $X2=0 $Y2=0
cc_269 N_A_340_309#_c_396_n N_Z_c_441_n 0.0129692f $X=3.375 $Y=2.2 $X2=0 $Y2=0
cc_270 N_Z_c_436_n N_VGND_c_497_n 0.00121826f $X=4.345 $Y=0.855 $X2=0 $Y2=0
cc_271 N_Z_M1005_s N_VGND_c_498_n 0.00298338f $X=3.575 $Y=0.235 $X2=0 $Y2=0
cc_272 N_Z_c_436_n N_VGND_c_498_n 0.00223842f $X=4.345 $Y=0.855 $X2=0 $Y2=0
cc_273 N_Z_c_449_n N_A_412_47#_M1011_d 0.00222098f $X=4.23 $Y=0.745 $X2=0 $Y2=0
cc_274 Z N_A_412_47#_M1011_d 4.69901e-19 $X=4.245 $Y=0.765 $X2=0 $Y2=0
cc_275 N_Z_c_436_n N_A_412_47#_M1011_d 0.00230798f $X=4.345 $Y=0.855 $X2=0 $Y2=0
cc_276 N_Z_c_440_n N_A_412_47#_c_556_n 0.00220399f $X=3.595 $Y=1.605 $X2=0 $Y2=0
cc_277 N_Z_M1005_s N_A_412_47#_c_552_n 0.00512757f $X=3.575 $Y=0.235 $X2=0 $Y2=0
cc_278 N_Z_c_449_n N_A_412_47#_c_552_n 0.0348928f $X=4.23 $Y=0.745 $X2=0 $Y2=0
cc_279 N_Z_c_436_n N_A_412_47#_c_552_n 0.0132977f $X=4.345 $Y=0.855 $X2=0 $Y2=0
cc_280 N_VGND_c_498_n N_A_412_47#_M1001_s 0.00333218f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_281 N_VGND_c_498_n N_A_412_47#_M1004_s 0.00390995f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_498_n N_A_412_47#_M1011_d 0.00210181f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_494_n N_A_412_47#_c_550_n 0.0179998f $X=2.705 $Y=0.36 $X2=0
+ $Y2=0
cc_284 N_VGND_c_496_n N_A_412_47#_c_550_n 0.0222373f $X=2.49 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_498_n N_A_412_47#_c_550_n 0.0122068f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_M1001_d N_A_412_47#_c_556_n 0.00293186f $X=2.57 $Y=0.235 $X2=0
+ $Y2=0
cc_287 N_VGND_c_494_n N_A_412_47#_c_556_n 0.0198656f $X=2.705 $Y=0.36 $X2=0
+ $Y2=0
cc_288 N_VGND_c_496_n N_A_412_47#_c_556_n 0.00234591f $X=2.49 $Y=0 $X2=0 $Y2=0
cc_289 N_VGND_c_497_n N_A_412_47#_c_556_n 0.00313531f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_290 N_VGND_c_498_n N_A_412_47#_c_556_n 0.0116556f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_291 N_VGND_c_494_n N_A_412_47#_c_562_n 0.00124003f $X=2.705 $Y=0.36 $X2=0
+ $Y2=0
cc_292 N_VGND_c_494_n N_A_412_47#_c_563_n 0.0129887f $X=2.705 $Y=0.36 $X2=0
+ $Y2=0
cc_293 N_VGND_c_497_n N_A_412_47#_c_563_n 0.0173458f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_294 N_VGND_c_498_n N_A_412_47#_c_563_n 0.0108223f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_295 N_VGND_c_497_n N_A_412_47#_c_552_n 0.0520305f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_296 N_VGND_c_498_n N_A_412_47#_c_552_n 0.0363595f $X=4.37 $Y=0 $X2=0 $Y2=0
