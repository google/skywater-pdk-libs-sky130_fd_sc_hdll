* File: sky130_fd_sc_hdll__a22o_2.spice
* Created: Thu Aug 27 18:54:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a22o_2.pex.spice"
.subckt sky130_fd_sc_hdll__a22o_2  VNB VPB B2 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1009 A_119_47# N_B2_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65 AD=0.07475
+ AS=0.2015 PD=0.88 PS=1.92 NRD=11.076 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1010 N_A_27_297#_M1010_d N_B1_M1010_g A_119_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.07475 PD=1.92 PS=0.88 NRD=8.304 NRS=11.076 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 A_411_47# N_A1_M1006_g N_A_27_297#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.2015 PD=1.03 PS=1.92 NRD=24.912 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g A_411_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.118625 AS=0.1235 PD=1.015 PS=1.03 NRD=0 NRS=24.912 M=1 R=4.33333
+ SA=75000.8 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1007_d N_A_27_297#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.118625 AS=0.104 PD=1.015 PS=0.97 NRD=16.608 NRS=0 M=1 R=4.33333
+ SA=75001.3 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_27_297#_M1004_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.25675 AS=0.104 PD=2.09 PS=0.97 NRD=23.988 NRS=8.304 M=1 R=4.33333
+ SA=75001.7 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1005 N_A_117_297#_M1005_d N_B2_M1005_g N_A_27_297#_M1005_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1000 N_A_27_297#_M1000_d N_B1_M1000_g N_A_117_297#_M1005_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_A_117_297#_M1008_d N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.27 PD=1.35 PS=2.54 NRD=5.8903 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_117_297#_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1675 AS=0.175 PD=1.335 PS=1.35 NRD=9.8303 NRS=7.8603 M=1 R=5.55556
+ SA=90000.7 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1001 N_X_M1001_d N_A_27_297#_M1001_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.1675 PD=1.29 PS=1.335 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1011 N_X_M1001_d N_A_27_297#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.405 PD=1.29 PS=2.81 NRD=0.9653 NRS=27.5603 M=1 R=5.55556
+ SA=90001.7 SB=90000.3 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__a22o_2.pxi.spice"
*
.ends
*
*
