* File: sky130_fd_sc_hdll__nand3_4.pex.spice
* Created: Thu Aug 27 19:13:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND3_4%C 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 37 51 59 62
c83 32 0 1.98913e-19 $X=1.535 $Y=1.105
r84 51 52 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=1.93 $Y2=1.217
r85 49 51 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=1.67 $Y=1.217
+ $X2=1.905 $Y2=1.217
r86 47 49 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=1.46 $Y=1.217
+ $X2=1.67 $Y2=1.217
r87 46 47 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.217
+ $X2=1.46 $Y2=1.217
r88 45 46 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=0.99 $Y=1.217
+ $X2=1.435 $Y2=1.217
r89 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.217
+ $X2=0.99 $Y2=1.217
r90 43 44 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.217
+ $X2=0.965 $Y2=1.217
r91 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.217
+ $X2=0.52 $Y2=1.217
r92 37 42 16.3472 $w=3.27e-07 $l=1.253e-07 $layer=POLY_cond $X=0.395 $Y=1.16
+ $X2=0.495 $Y2=1.217
r93 37 39 26.6608 $w=2.7e-07 $l=1.2e-07 $layer=POLY_cond $X=0.395 $Y=1.16
+ $X2=0.275 $Y2=1.16
r94 32 62 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=1.62 $Y=1.175
+ $X2=1.615 $Y2=1.175
r95 32 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.67
+ $Y=1.16 $X2=1.67 $Y2=1.16
r96 31 62 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=1.16 $Y=1.175
+ $X2=1.615 $Y2=1.175
r97 31 59 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=1.16 $Y=1.175
+ $X2=1.155 $Y2=1.175
r98 30 59 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=1.155 $Y2=1.175
r99 29 30 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r100 29 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r101 25 52 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r102 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r103 22 51 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r104 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r105 18 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.217
r106 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r107 15 46 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.217
r108 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r109 11 45 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=1.217
r110 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=0.56
r111 8 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.217
r112 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r113 4 43 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=1.217
r114 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=0.56
r115 1 42 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.217
r116 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_4%B 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 32 49 52 56 59 64
c85 49 0 1.98913e-19 $X=3.785 $Y=1.217
r86 49 50 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.217
+ $X2=3.81 $Y2=1.217
r87 47 49 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=3.55 $Y=1.217
+ $X2=3.785 $Y2=1.217
r88 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.16 $X2=3.55 $Y2=1.16
r89 45 47 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=3.315 $Y=1.217
+ $X2=3.55 $Y2=1.217
r90 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.217
+ $X2=3.315 $Y2=1.217
r91 43 44 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=3.29 $Y2=1.217
r92 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.217
+ $X2=2.845 $Y2=1.217
r93 40 42 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=2.61 $Y=1.217
+ $X2=2.82 $Y2=1.217
r94 38 40 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.61 $Y2=1.217
r95 37 38 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r96 32 64 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=3.91 $Y=1.175 $X2=3.93
+ $Y2=1.175
r97 32 48 19.9636 $w=1.98e-07 $l=3.6e-07 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=3.55 $Y2=1.175
r98 31 48 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=3.46 $Y=1.175 $X2=3.55
+ $Y2=1.175
r99 31 59 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=3.46 $Y=1.175 $X2=3.41
+ $Y2=1.175
r100 30 59 23.5682 $w=1.98e-07 $l=4.25e-07 $layer=LI1_cond $X=2.985 $Y=1.175
+ $X2=3.41 $Y2=1.175
r101 30 56 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.985 $Y=1.175
+ $X2=2.97 $Y2=1.175
r102 29 56 24.4 $w=1.98e-07 $l=4.4e-07 $layer=LI1_cond $X=2.53 $Y=1.175 $X2=2.97
+ $Y2=1.175
r103 29 52 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=2.53 $Y=1.175
+ $X2=2.525 $Y2=1.175
r104 29 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.16 $X2=2.61 $Y2=1.16
r105 25 50 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=1.217
r106 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=0.56
r107 22 49 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.217
r108 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r109 19 45 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r110 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r111 15 44 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r112 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r113 12 43 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r114 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r115 8 42 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=1.217
r116 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.82 $Y=1.025
+ $X2=2.82 $Y2=0.56
r117 5 38 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r118 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r119 1 37 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r120 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 37 51 58 62 66
r78 51 52 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.185 $Y=1.217
+ $X2=6.21 $Y2=1.217
r79 50 62 10.8136 $w=1.98e-07 $l=1.95e-07 $layer=LI1_cond $X=5.95 $Y=1.175
+ $X2=5.755 $Y2=1.175
r80 49 51 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=5.95 $Y=1.217
+ $X2=6.185 $Y2=1.217
r81 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.95
+ $Y=1.16 $X2=5.95 $Y2=1.16
r82 47 49 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=5.74 $Y=1.217
+ $X2=5.95 $Y2=1.217
r83 46 47 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.715 $Y=1.217
+ $X2=5.74 $Y2=1.217
r84 45 46 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=5.27 $Y=1.217
+ $X2=5.715 $Y2=1.217
r85 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.245 $Y=1.217
+ $X2=5.27 $Y2=1.217
r86 43 44 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=4.8 $Y=1.217
+ $X2=5.245 $Y2=1.217
r87 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.217
+ $X2=4.8 $Y2=1.217
r88 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.51
+ $Y=1.16 $X2=4.51 $Y2=1.16
r89 37 42 16.3472 $w=3.27e-07 $l=1.253e-07 $layer=POLY_cond $X=4.675 $Y=1.16
+ $X2=4.775 $Y2=1.217
r90 37 39 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.675 $Y=1.16
+ $X2=4.51 $Y2=1.16
r91 32 66 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=6.215 $Y=1.175
+ $X2=6.235 $Y2=1.175
r92 32 50 14.6955 $w=1.98e-07 $l=2.65e-07 $layer=LI1_cond $X=6.215 $Y=1.175
+ $X2=5.95 $Y2=1.175
r93 31 62 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=5.75 $Y=1.175
+ $X2=5.755 $Y2=1.175
r94 30 31 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=5.295 $Y=1.175
+ $X2=5.75 $Y2=1.175
r95 30 58 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=5.295 $Y=1.175
+ $X2=5.29 $Y2=1.175
r96 29 58 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=4.835 $Y=1.175
+ $X2=5.29 $Y2=1.175
r97 29 40 18.0227 $w=1.98e-07 $l=3.25e-07 $layer=LI1_cond $X=4.835 $Y=1.175
+ $X2=4.51 $Y2=1.175
r98 25 52 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.21 $Y=1.025
+ $X2=6.21 $Y2=1.217
r99 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.21 $Y=1.025
+ $X2=6.21 $Y2=0.56
r100 22 51 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.217
r101 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r102 18 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.74 $Y=1.025
+ $X2=5.74 $Y2=1.217
r103 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.74 $Y=1.025
+ $X2=5.74 $Y2=0.56
r104 15 46 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.217
r105 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r106 11 45 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.27 $Y=1.025
+ $X2=5.27 $Y2=1.217
r107 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.27 $Y=1.025
+ $X2=5.27 $Y2=0.56
r108 8 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.217
r109 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r110 4 43 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.8 $Y=1.025
+ $X2=4.8 $Y2=1.217
r111 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.8 $Y=1.025 $X2=4.8
+ $Y2=0.56
r112 1 42 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.217
r113 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_4%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 37 41 45
+ 49 54 58 61 62 64 65 67 68 69 75 87 88 94 97 100
r107 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r108 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r109 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r110 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r111 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r112 85 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r113 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r114 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r115 82 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r116 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r117 79 100 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.28 $Y2=2.72
r118 79 81 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=5.29 $Y2=2.72
r119 78 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r120 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r121 75 100 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=4.28 $Y2=2.72
r122 75 77 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=3.91 $Y2=2.72
r123 74 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r124 74 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r125 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r126 71 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.14 $Y2=2.72
r127 71 73 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.99 $Y2=2.72
r128 69 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r129 69 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r130 67 84 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=2.72
+ $X2=6.21 $Y2=2.72
r131 67 68 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=6.335 $Y=2.72
+ $X2=6.467 $Y2=2.72
r132 66 87 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.6 $Y=2.72 $X2=6.67
+ $Y2=2.72
r133 66 68 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=6.6 $Y=2.72
+ $X2=6.467 $Y2=2.72
r134 64 81 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=2.72
+ $X2=5.29 $Y2=2.72
r135 64 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=2.72
+ $X2=5.48 $Y2=2.72
r136 63 84 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=2.72
+ $X2=6.21 $Y2=2.72
r137 63 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=2.72
+ $X2=5.48 $Y2=2.72
r138 61 73 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=2.99 $Y2=2.72
r139 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=3.08 $Y2=2.72
r140 60 77 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.91 $Y2=2.72
r141 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.08 $Y2=2.72
r142 56 68 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=6.467 $Y=2.635
+ $X2=6.467 $Y2=2.72
r143 56 58 27.6151 $w=2.63e-07 $l=6.35e-07 $layer=LI1_cond $X=6.467 $Y=2.635
+ $X2=6.467 $Y2=2
r144 52 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r145 52 54 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2
r146 47 100 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=2.635
+ $X2=4.28 $Y2=2.72
r147 47 49 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=4.28 $Y=2.635
+ $X2=4.28 $Y2=2
r148 43 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r149 43 45 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r150 39 97 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r151 39 41 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r152 38 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.2 $Y2=2.72
r153 37 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.14 $Y2=2.72
r154 37 38 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r155 33 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r156 33 35 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r157 32 91 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r158 31 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.2 $Y2=2.72
r159 31 32 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r160 27 30 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r161 25 91 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r162 25 30 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r163 8 58 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2
r164 7 54 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2
r165 6 49 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=4.415
+ $Y=1.485 $X2=4.54 $Y2=2
r166 5 49 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2
r167 4 45 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r168 3 41 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r169 2 35 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r170 1 30 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r171 1 27 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_4%Y 1 2 3 4 5 6 7 8 25 27 29 33 35 39 41 45
+ 47 49 57 59 63 65 70 72 74 76 78 79 80 81 87
r157 80 81 9.41096 $w=3.98e-07 $l=2.55e-07 $layer=LI1_cond $X=6.67 $Y=1.19
+ $X2=6.67 $Y2=1.445
r158 79 87 3.55828 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=6.67 $Y=0.78
+ $X2=6.67 $Y2=0.905
r159 79 80 13.5287 $w=2.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.67 $Y=0.92
+ $X2=6.67 $Y2=1.19
r160 79 87 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.67 $Y=0.92
+ $X2=6.67 $Y2=0.905
r161 66 78 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=6.115 $Y=1.555
+ $X2=5.925 $Y2=1.555
r162 65 81 3.48622 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=6.555 $Y=1.555
+ $X2=6.67 $Y2=1.555
r163 65 66 23.0489 $w=2.18e-07 $l=4.4e-07 $layer=LI1_cond $X=6.555 $Y=1.555
+ $X2=6.115 $Y2=1.555
r164 61 78 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=5.925 $Y=1.665
+ $X2=5.925 $Y2=1.555
r165 61 63 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=5.925 $Y=1.665
+ $X2=5.925 $Y2=2.34
r166 60 76 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=1.555
+ $X2=4.985 $Y2=1.555
r167 59 78 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.735 $Y=1.555
+ $X2=5.925 $Y2=1.555
r168 59 60 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=5.735 $Y=1.555
+ $X2=5.175 $Y2=1.555
r169 55 76 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=4.985 $Y=1.665
+ $X2=4.985 $Y2=1.555
r170 55 57 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.985 $Y=1.665
+ $X2=4.985 $Y2=2.34
r171 51 54 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.01 $Y=0.78
+ $X2=5.95 $Y2=0.78
r172 49 79 3.27362 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=6.555 $Y=0.78
+ $X2=6.67 $Y2=0.78
r173 49 54 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=6.555 $Y=0.78
+ $X2=5.95 $Y2=0.78
r174 48 74 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=1.555
+ $X2=3.525 $Y2=1.555
r175 47 76 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.795 $Y=1.555
+ $X2=4.985 $Y2=1.555
r176 47 48 56.5745 $w=2.18e-07 $l=1.08e-06 $layer=LI1_cond $X=4.795 $Y=1.555
+ $X2=3.715 $Y2=1.555
r177 43 74 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=1.555
r178 43 45 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=2.34
r179 42 72 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=1.555
+ $X2=2.585 $Y2=1.555
r180 41 74 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=1.555
+ $X2=3.525 $Y2=1.555
r181 41 42 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=3.335 $Y=1.555
+ $X2=2.775 $Y2=1.555
r182 37 72 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=2.585 $Y=1.665
+ $X2=2.585 $Y2=1.555
r183 37 39 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.585 $Y=1.665
+ $X2=2.585 $Y2=2.34
r184 36 70 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.555
+ $X2=1.645 $Y2=1.555
r185 35 72 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=1.555
+ $X2=2.585 $Y2=1.555
r186 35 36 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=2.395 $Y=1.555
+ $X2=1.835 $Y2=1.555
r187 31 70 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=1.555
r188 31 33 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=2.34
r189 30 68 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.555
+ $X2=0.705 $Y2=1.555
r190 29 70 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=1.645 $Y2=1.555
r191 29 30 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=0.895 $Y2=1.555
r192 25 68 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.555
r193 25 27 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r194 8 78 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.66
r195 8 63 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=2.34
r196 7 76 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.66
r197 7 57 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.34
r198 6 74 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.66
r199 6 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.34
r200 5 72 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r201 5 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r202 4 70 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r203 4 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r204 3 68 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r205 3 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r206 2 54 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.235 $X2=5.95 $Y2=0.74
r207 1 51 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_4%A_27_47# 1 2 3 4 5 18 20 21 24 32 35 36 39
+ 40 42 43
r80 42 43 11.0982 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=4.02 $Y=0.78
+ $X2=3.805 $Y2=0.78
r81 40 43 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.245 $Y=0.82
+ $X2=3.805 $Y2=0.82
r82 38 40 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=0.78
+ $X2=3.245 $Y2=0.78
r83 38 39 11.0982 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=3.08 $Y=0.78
+ $X2=2.865 $Y2=0.78
r84 36 39 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.305 $Y=0.82
+ $X2=2.865 $Y2=0.82
r85 34 36 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=0.78
+ $X2=2.305 $Y2=0.78
r86 34 35 11.0982 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=2.14 $Y=0.78
+ $X2=1.925 $Y2=0.78
r87 27 32 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0.82
+ $X2=1.175 $Y2=0.82
r88 27 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.365 $Y=0.82
+ $X2=1.925 $Y2=0.82
r89 22 32 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=0.735
+ $X2=1.175 $Y2=0.82
r90 22 24 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.175 $Y=0.735
+ $X2=1.175 $Y2=0.4
r91 20 32 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0.82
+ $X2=1.175 $Y2=0.82
r92 20 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.82
+ $X2=0.425 $Y2=0.82
r93 16 21 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.425 $Y2=0.82
r94 16 18 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.4
r95 5 42 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.74
r96 4 38 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.74
r97 3 34 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.74
r98 2 24 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.4
r99 1 18 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_4%VGND 1 2 11 13 17 19 26 27 30 33 36
r71 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r72 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r73 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r74 26 27 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r75 24 27 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=6.67
+ $Y2=0
r76 24 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r77 23 26 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=6.67
+ $Y2=0
r78 23 24 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r79 21 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.67
+ $Y2=0
r80 21 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.755 $Y=0 $X2=2.07
+ $Y2=0
r81 19 31 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r82 19 36 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r83 15 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r84 15 17 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.4
r85 14 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r86 13 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.67
+ $Y2=0
r87 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=0.815
+ $Y2=0
r88 9 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085 $X2=0.73
+ $Y2=0
r89 9 11 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.4
r90 2 17 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.4
r91 1 11 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_4%A_485_47# 1 2 3 4 5 26
r34 24 26 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=5.48 $Y=0.37
+ $X2=6.42 $Y2=0.37
r35 22 24 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=4.54 $Y=0.37
+ $X2=5.48 $Y2=0.37
r36 20 22 49.6052 $w=2.28e-07 $l=9.9e-07 $layer=LI1_cond $X=3.55 $Y=0.37
+ $X2=4.54 $Y2=0.37
r37 17 20 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=2.61 $Y=0.37
+ $X2=3.55 $Y2=0.37
r38 5 26 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.235 $X2=6.42 $Y2=0.4
r39 4 24 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.235 $X2=5.48 $Y2=0.4
r40 3 22 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=4.415
+ $Y=0.235 $X2=4.54 $Y2=0.4
r41 2 20 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.4
r42 1 17 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.4
.ends

