* File: sky130_fd_sc_hdll__buf_6.pxi.spice
* Created: Wed Sep  2 08:24:30 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUF_6%A N_A_c_75_n N_A_M1001_g N_A_M1007_g N_A_c_76_n
+ N_A_M1002_g N_A_M1009_g A A N_A_c_73_n N_A_c_74_n A
+ PM_SKY130_FD_SC_HDLL__BUF_6%A
x_PM_SKY130_FD_SC_HDLL__BUF_6%A_169_297# N_A_169_297#_M1007_s
+ N_A_169_297#_M1001_s N_A_169_297#_M1000_g N_A_169_297#_c_131_n
+ N_A_169_297#_M1003_g N_A_169_297#_M1004_g N_A_169_297#_c_132_n
+ N_A_169_297#_M1008_g N_A_169_297#_M1005_g N_A_169_297#_c_133_n
+ N_A_169_297#_M1010_g N_A_169_297#_M1006_g N_A_169_297#_c_134_n
+ N_A_169_297#_M1013_g N_A_169_297#_M1011_g N_A_169_297#_c_135_n
+ N_A_169_297#_M1014_g N_A_169_297#_c_136_n N_A_169_297#_M1015_g
+ N_A_169_297#_M1012_g N_A_169_297#_c_142_n N_A_169_297#_c_137_n
+ N_A_169_297#_c_147_n N_A_169_297#_c_125_n N_A_169_297#_c_126_n
+ N_A_169_297#_c_154_n N_A_169_297#_c_127_n N_A_169_297#_c_128_n
+ N_A_169_297#_c_206_p N_A_169_297#_c_129_n N_A_169_297#_c_130_n
+ PM_SKY130_FD_SC_HDLL__BUF_6%A_169_297#
x_PM_SKY130_FD_SC_HDLL__BUF_6%VPWR N_VPWR_M1001_d N_VPWR_M1002_d N_VPWR_M1008_d
+ N_VPWR_M1013_d N_VPWR_M1015_d N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n
+ N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n
+ N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n
+ N_VPWR_c_284_n VPWR VPWR N_VPWR_c_285_n N_VPWR_c_270_n
+ PM_SKY130_FD_SC_HDLL__BUF_6%VPWR
x_PM_SKY130_FD_SC_HDLL__BUF_6%X N_X_M1000_s N_X_M1005_s N_X_M1011_s N_X_M1003_s
+ N_X_M1010_s N_X_M1014_s N_X_c_358_n N_X_c_359_n N_X_c_352_n N_X_c_353_n
+ N_X_c_355_n N_X_c_356_n N_X_c_375_n N_X_c_377_n N_X_c_380_n N_X_c_383_n X X
+ N_X_c_354_n PM_SKY130_FD_SC_HDLL__BUF_6%X
x_PM_SKY130_FD_SC_HDLL__BUF_6%VGND N_VGND_M1007_d N_VGND_M1009_d N_VGND_M1004_d
+ N_VGND_M1006_d N_VGND_M1012_d N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n
+ N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n
+ N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_455_n
+ N_VGND_c_456_n VGND VGND N_VGND_c_457_n N_VGND_c_458_n
+ PM_SKY130_FD_SC_HDLL__BUF_6%VGND
cc_1 VNB N_A_M1007_g 0.0248167f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.56
cc_2 VNB N_A_M1009_g 0.01806f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=0.56
cc_3 VNB A 0.0109395f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.105
cc_4 VNB N_A_c_73_n 0.040848f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_5 VNB N_A_c_74_n 0.0392529f $X=-0.19 $Y=-0.24 $X2=1.225 $Y2=1.217
cc_6 VNB N_A_169_297#_M1000_g 0.0174966f $X=-0.19 $Y=-0.24 $X2=1.225 $Y2=1.985
cc_7 VNB N_A_169_297#_M1004_g 0.0181101f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.105
cc_8 VNB N_A_169_297#_M1005_g 0.017151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_169_297#_M1006_g 0.017151f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.217
cc_10 VNB N_A_169_297#_M1011_g 0.0176309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_169_297#_M1012_g 0.0241263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_169_297#_c_125_n 0.00196295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_169_297#_c_126_n 0.00233388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_169_297#_c_127_n 0.00157323f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_169_297#_c_128_n 3.60034e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_169_297#_c_129_n 0.00104338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_169_297#_c_130_n 0.15487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_270_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_352_n 0.00265585f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.16
cc_20 VNB N_X_c_353_n 0.00143033f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.16
cc_21 VNB N_X_c_354_n 0.00257172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_443_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_444_n 0.0041632f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_24 VNB N_VGND_c_445_n 3.32195e-19 $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.217
cc_25 VNB N_VGND_c_446_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.217
cc_26 VNB N_VGND_c_447_n 0.0129158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_448_n 0.0321553f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.195
cc_28 VNB N_VGND_c_449_n 0.0159859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_450_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_451_n 0.0199309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_452_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_453_n 0.0167592f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_454_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_455_n 0.0126629f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_456_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_457_n 0.0132691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_458_n 0.252158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_A_c_75_n 0.021061f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.41
cc_39 VPB N_A_c_76_n 0.0163655f $X=-0.19 $Y=1.305 $X2=1.225 $Y2=1.41
cc_40 VPB A 0.0118256f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.105
cc_41 VPB N_A_c_74_n 0.0161045f $X=-0.19 $Y=1.305 $X2=1.225 $Y2=1.217
cc_42 VPB N_A_169_297#_c_131_n 0.015821f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=1.025
cc_43 VPB N_A_169_297#_c_132_n 0.0154384f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_169_297#_c_133_n 0.0154273f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.217
cc_45 VPB N_A_169_297#_c_134_n 0.015148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_169_297#_c_135_n 0.0154273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_169_297#_c_136_n 0.0198847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_169_297#_c_137_n 0.00109065f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_169_297#_c_128_n 0.00165083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_169_297#_c_130_n 0.0388785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_271_n 0.00573847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_272_n 0.00234463f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.217
cc_53 VPB N_VPWR_c_273_n 3.21306e-19 $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.16
cc_54 VPB N_VPWR_c_274_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_275_n 0.0129491f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.195
cc_56 VPB N_VPWR_c_276_n 0.0461502f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=1.195
cc_57 VPB N_VPWR_c_277_n 0.0159859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_278_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_279_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_280_n 0.00346606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_281_n 0.0144008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_282_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_283_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_284_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_285_n 0.0140698f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_270_n 0.0581173f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_X_c_355_n 0.00168548f $X=-0.19 $Y=1.305 $X2=1.225 $Y2=1.217
cc_68 VPB N_X_c_356_n 0.00148018f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=1.217
cc_69 VPB N_X_c_354_n 0.00296714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 N_A_M1009_g N_A_169_297#_M1000_g 0.0219275f $X=1.25 $Y=0.56 $X2=0 $Y2=0
cc_71 N_A_c_76_n N_A_169_297#_c_131_n 0.0223825f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_M1007_g N_A_169_297#_c_142_n 0.0132993f $X=0.78 $Y=0.56 $X2=0 $Y2=0
cc_73 N_A_c_75_n N_A_169_297#_c_137_n 0.00347232f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_76_n N_A_169_297#_c_137_n 5.79575e-19 $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_75 A N_A_169_297#_c_137_n 0.0263123f $X=0.94 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_c_74_n N_A_169_297#_c_137_n 0.00174157f $X=1.225 $Y=1.217 $X2=0 $Y2=0
cc_77 N_A_c_75_n N_A_169_297#_c_147_n 0.0123129f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_c_76_n N_A_169_297#_c_147_n 0.0108994f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_M1009_g N_A_169_297#_c_125_n 0.0110972f $X=1.25 $Y=0.56 $X2=0 $Y2=0
cc_80 A N_A_169_297#_c_125_n 0.00769632f $X=0.94 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A_M1007_g N_A_169_297#_c_126_n 0.0101476f $X=0.78 $Y=0.56 $X2=0 $Y2=0
cc_82 A N_A_169_297#_c_126_n 0.0308888f $X=0.94 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A_c_74_n N_A_169_297#_c_126_n 0.00332f $X=1.225 $Y=1.217 $X2=0 $Y2=0
cc_84 N_A_c_76_n N_A_169_297#_c_154_n 0.0143733f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_85 A N_A_169_297#_c_154_n 0.00762487f $X=0.94 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_M1009_g N_A_169_297#_c_127_n 0.0037087f $X=1.25 $Y=0.56 $X2=0 $Y2=0
cc_87 N_A_c_76_n N_A_169_297#_c_128_n 0.00160748f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_88 A N_A_169_297#_c_128_n 0.00503213f $X=0.94 $Y=1.105 $X2=0 $Y2=0
cc_89 N_A_c_74_n N_A_169_297#_c_128_n 0.00259641f $X=1.225 $Y=1.217 $X2=0 $Y2=0
cc_90 A N_A_169_297#_c_129_n 0.0135589f $X=0.94 $Y=1.105 $X2=0 $Y2=0
cc_91 N_A_c_74_n N_A_169_297#_c_129_n 0.00144938f $X=1.225 $Y=1.217 $X2=0 $Y2=0
cc_92 A N_A_169_297#_c_130_n 2.17837e-19 $X=0.94 $Y=1.105 $X2=0 $Y2=0
cc_93 N_A_c_74_n N_A_169_297#_c_130_n 0.0219275f $X=1.225 $Y=1.217 $X2=0 $Y2=0
cc_94 N_A_c_75_n N_VPWR_c_271_n 0.00739257f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_95 A N_VPWR_c_271_n 0.0142331f $X=0.94 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A_c_73_n N_VPWR_c_271_n 0.00126394f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_c_76_n N_VPWR_c_272_n 0.00551021f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_c_75_n N_VPWR_c_279_n 0.00597712f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_c_76_n N_VPWR_c_279_n 0.00673617f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_c_75_n N_VPWR_c_270_n 0.0110738f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_76_n N_VPWR_c_270_n 0.011869f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_M1007_g N_VGND_c_443_n 0.00512729f $X=0.78 $Y=0.56 $X2=0 $Y2=0
cc_103 A N_VGND_c_443_n 0.00575903f $X=0.94 $Y=1.105 $X2=0 $Y2=0
cc_104 N_A_c_73_n N_VGND_c_443_n 0.0031817f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_M1009_g N_VGND_c_444_n 0.00268723f $X=1.25 $Y=0.56 $X2=0 $Y2=0
cc_106 N_A_M1007_g N_VGND_c_451_n 0.00465454f $X=0.78 $Y=0.56 $X2=0 $Y2=0
cc_107 N_A_M1009_g N_VGND_c_451_n 0.00439206f $X=1.25 $Y=0.56 $X2=0 $Y2=0
cc_108 N_A_M1007_g N_VGND_c_458_n 0.00904947f $X=0.78 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A_M1009_g N_VGND_c_458_n 0.00606547f $X=1.25 $Y=0.56 $X2=0 $Y2=0
cc_110 N_A_169_297#_c_154_n N_VPWR_M1002_d 0.00340529f $X=1.455 $Y=1.57 $X2=0
+ $Y2=0
cc_111 N_A_169_297#_c_137_n N_VPWR_c_271_n 0.0133617f $X=0.965 $Y=1.655 $X2=0
+ $Y2=0
cc_112 N_A_169_297#_c_147_n N_VPWR_c_271_n 0.0604323f $X=0.99 $Y=2.31 $X2=0
+ $Y2=0
cc_113 N_A_169_297#_c_131_n N_VPWR_c_272_n 0.010617f $X=1.695 $Y=1.41 $X2=0
+ $Y2=0
cc_114 N_A_169_297#_c_132_n N_VPWR_c_272_n 6.4992e-19 $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_115 N_A_169_297#_c_147_n N_VPWR_c_272_n 0.0395636f $X=0.99 $Y=2.31 $X2=0
+ $Y2=0
cc_116 N_A_169_297#_c_154_n N_VPWR_c_272_n 0.0148423f $X=1.455 $Y=1.57 $X2=0
+ $Y2=0
cc_117 N_A_169_297#_c_131_n N_VPWR_c_273_n 7.03572e-19 $X=1.695 $Y=1.41 $X2=0
+ $Y2=0
cc_118 N_A_169_297#_c_132_n N_VPWR_c_273_n 0.0154767f $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_169_297#_c_133_n N_VPWR_c_273_n 0.0117385f $X=2.635 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_A_169_297#_c_134_n N_VPWR_c_273_n 6.61031e-19 $X=3.105 $Y=1.41 $X2=0
+ $Y2=0
cc_121 N_A_169_297#_c_130_n N_VPWR_c_273_n 4.16178e-19 $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_122 N_A_169_297#_c_133_n N_VPWR_c_274_n 6.99539e-19 $X=2.635 $Y=1.41 $X2=0
+ $Y2=0
cc_123 N_A_169_297#_c_134_n N_VPWR_c_274_n 0.0154534f $X=3.105 $Y=1.41 $X2=0
+ $Y2=0
cc_124 N_A_169_297#_c_135_n N_VPWR_c_274_n 0.0117392f $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_125 N_A_169_297#_c_136_n N_VPWR_c_274_n 6.61031e-19 $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_126 N_A_169_297#_c_130_n N_VPWR_c_274_n 9.18523e-19 $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_127 N_A_169_297#_c_135_n N_VPWR_c_276_n 8.37274e-19 $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A_169_297#_c_136_n N_VPWR_c_276_n 0.022204f $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_129 N_A_169_297#_c_147_n N_VPWR_c_279_n 0.0223557f $X=0.99 $Y=2.31 $X2=0
+ $Y2=0
cc_130 N_A_169_297#_c_131_n N_VPWR_c_281_n 0.00661659f $X=1.695 $Y=1.41 $X2=0
+ $Y2=0
cc_131 N_A_169_297#_c_132_n N_VPWR_c_281_n 0.00427505f $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_132 N_A_169_297#_c_133_n N_VPWR_c_283_n 0.00622633f $X=2.635 $Y=1.41 $X2=0
+ $Y2=0
cc_133 N_A_169_297#_c_134_n N_VPWR_c_283_n 0.00427505f $X=3.105 $Y=1.41 $X2=0
+ $Y2=0
cc_134 N_A_169_297#_c_135_n N_VPWR_c_285_n 0.00622633f $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_135 N_A_169_297#_c_136_n N_VPWR_c_285_n 0.00427505f $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_136 N_A_169_297#_M1001_s N_VPWR_c_270_n 0.00231261f $X=0.845 $Y=1.485 $X2=0
+ $Y2=0
cc_137 N_A_169_297#_c_131_n N_VPWR_c_270_n 0.0110933f $X=1.695 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_A_169_297#_c_132_n N_VPWR_c_270_n 0.00740765f $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_169_297#_c_133_n N_VPWR_c_270_n 0.010479f $X=2.635 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_169_297#_c_134_n N_VPWR_c_270_n 0.00740765f $X=3.105 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_169_297#_c_135_n N_VPWR_c_270_n 0.010479f $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_169_297#_c_136_n N_VPWR_c_270_n 0.00740765f $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_143 N_A_169_297#_c_147_n N_VPWR_c_270_n 0.0140101f $X=0.99 $Y=2.31 $X2=0
+ $Y2=0
cc_144 N_A_169_297#_M1000_g N_X_c_358_n 0.00494213f $X=1.67 $Y=0.56 $X2=0 $Y2=0
cc_145 N_A_169_297#_c_131_n N_X_c_359_n 0.00649064f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_169_297#_c_132_n N_X_c_359_n 0.00657309f $X=2.165 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_169_297#_c_154_n N_X_c_359_n 0.00254387f $X=1.455 $Y=1.57 $X2=0 $Y2=0
cc_148 N_A_169_297#_M1004_g N_X_c_352_n 0.0132715f $X=2.14 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A_169_297#_c_130_n N_X_c_352_n 0.00282955f $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_150 N_A_169_297#_M1000_g N_X_c_353_n 0.0014017f $X=1.67 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A_169_297#_c_125_n N_X_c_353_n 0.012198f $X=1.455 $Y=0.82 $X2=0 $Y2=0
cc_152 N_A_169_297#_c_206_p N_X_c_353_n 0.0104474f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_169_297#_c_130_n N_X_c_353_n 0.00308294f $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_154 N_A_169_297#_c_132_n N_X_c_355_n 0.0164347f $X=2.165 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_169_297#_c_130_n N_X_c_355_n 0.00621759f $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_156 N_A_169_297#_c_131_n N_X_c_356_n 0.00133484f $X=1.695 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_169_297#_c_154_n N_X_c_356_n 0.0092999f $X=1.455 $Y=1.57 $X2=0 $Y2=0
cc_158 N_A_169_297#_c_128_n N_X_c_356_n 0.00263405f $X=1.54 $Y=1.485 $X2=0 $Y2=0
cc_159 N_A_169_297#_c_206_p N_X_c_356_n 0.00928734f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_169_297#_c_130_n N_X_c_356_n 0.00438538f $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_161 N_A_169_297#_M1005_g N_X_c_375_n 0.00464678f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A_169_297#_c_130_n N_X_c_375_n 4.53201e-19 $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_163 N_A_169_297#_c_133_n N_X_c_377_n 0.00704883f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_169_297#_c_134_n N_X_c_377_n 0.00659264f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_169_297#_c_130_n N_X_c_377_n 5.47843e-19 $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_166 N_A_169_297#_M1011_g N_X_c_380_n 0.00471006f $X=3.55 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A_169_297#_M1012_g N_X_c_380_n 0.0017519f $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A_169_297#_c_130_n N_X_c_380_n 5.90215e-19 $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_169 N_A_169_297#_c_135_n N_X_c_383_n 0.00704883f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_169_297#_c_136_n N_X_c_383_n 0.00289674f $X=4.045 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_169_297#_c_130_n N_X_c_383_n 5.50932e-19 $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_172 N_A_169_297#_M1004_g N_X_c_354_n 0.00192326f $X=2.14 $Y=0.56 $X2=0 $Y2=0
cc_173 N_A_169_297#_M1005_g N_X_c_354_n 0.0145245f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A_169_297#_c_133_n N_X_c_354_n 0.0163637f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_169_297#_M1006_g N_X_c_354_n 0.0149351f $X=3.08 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_169_297#_c_134_n N_X_c_354_n 0.014573f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_169_297#_M1011_g N_X_c_354_n 0.014543f $X=3.55 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A_169_297#_c_135_n N_X_c_354_n 0.015948f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_169_297#_c_136_n N_X_c_354_n 0.00320702f $X=4.045 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_169_297#_M1012_g N_X_c_354_n 0.00549657f $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A_169_297#_c_206_p N_X_c_354_n 0.00648218f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_169_297#_c_130_n N_X_c_354_n 0.108842f $X=4.045 $Y=1.217 $X2=0 $Y2=0
cc_183 N_A_169_297#_c_125_n N_VGND_M1009_d 0.00164499f $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_184 N_A_169_297#_c_142_n N_VGND_c_443_n 0.0231432f $X=0.99 $Y=0.38 $X2=0
+ $Y2=0
cc_185 N_A_169_297#_M1000_g N_VGND_c_444_n 0.00143136f $X=1.67 $Y=0.56 $X2=0
+ $Y2=0
cc_186 N_A_169_297#_c_125_n N_VGND_c_444_n 0.0128905f $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_187 N_A_169_297#_M1000_g N_VGND_c_445_n 5.94926e-19 $X=1.67 $Y=0.56 $X2=0
+ $Y2=0
cc_188 N_A_169_297#_M1004_g N_VGND_c_445_n 0.00824127f $X=2.14 $Y=0.56 $X2=0
+ $Y2=0
cc_189 N_A_169_297#_M1005_g N_VGND_c_445_n 0.00842493f $X=2.61 $Y=0.56 $X2=0
+ $Y2=0
cc_190 N_A_169_297#_M1006_g N_VGND_c_445_n 5.8773e-19 $X=3.08 $Y=0.56 $X2=0
+ $Y2=0
cc_191 N_A_169_297#_M1005_g N_VGND_c_446_n 5.66132e-19 $X=2.61 $Y=0.56 $X2=0
+ $Y2=0
cc_192 N_A_169_297#_M1006_g N_VGND_c_446_n 0.00806522f $X=3.08 $Y=0.56 $X2=0
+ $Y2=0
cc_193 N_A_169_297#_M1011_g N_VGND_c_446_n 0.00845883f $X=3.55 $Y=0.56 $X2=0
+ $Y2=0
cc_194 N_A_169_297#_M1012_g N_VGND_c_446_n 5.50819e-19 $X=4.07 $Y=0.56 $X2=0
+ $Y2=0
cc_195 N_A_169_297#_c_130_n N_VGND_c_446_n 5.8778e-19 $X=4.045 $Y=1.217 $X2=0
+ $Y2=0
cc_196 N_A_169_297#_M1011_g N_VGND_c_448_n 7.5279e-19 $X=3.55 $Y=0.56 $X2=0
+ $Y2=0
cc_197 N_A_169_297#_M1012_g N_VGND_c_448_n 0.0177043f $X=4.07 $Y=0.56 $X2=0
+ $Y2=0
cc_198 N_A_169_297#_c_142_n N_VGND_c_451_n 0.023074f $X=0.99 $Y=0.38 $X2=0 $Y2=0
cc_199 N_A_169_297#_c_125_n N_VGND_c_451_n 0.00248202f $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_200 N_A_169_297#_M1000_g N_VGND_c_453_n 0.00556122f $X=1.67 $Y=0.56 $X2=0
+ $Y2=0
cc_201 N_A_169_297#_M1004_g N_VGND_c_453_n 0.00350562f $X=2.14 $Y=0.56 $X2=0
+ $Y2=0
cc_202 N_A_169_297#_c_125_n N_VGND_c_453_n 8.04923e-19 $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_203 N_A_169_297#_M1005_g N_VGND_c_455_n 0.00350522f $X=2.61 $Y=0.56 $X2=0
+ $Y2=0
cc_204 N_A_169_297#_M1006_g N_VGND_c_455_n 0.00350562f $X=3.08 $Y=0.56 $X2=0
+ $Y2=0
cc_205 N_A_169_297#_M1011_g N_VGND_c_457_n 0.00350562f $X=3.55 $Y=0.56 $X2=0
+ $Y2=0
cc_206 N_A_169_297#_M1012_g N_VGND_c_457_n 0.00271402f $X=4.07 $Y=0.56 $X2=0
+ $Y2=0
cc_207 N_A_169_297#_M1007_s N_VGND_c_458_n 0.00264276f $X=0.855 $Y=0.235 $X2=0
+ $Y2=0
cc_208 N_A_169_297#_M1000_g N_VGND_c_458_n 0.00986515f $X=1.67 $Y=0.56 $X2=0
+ $Y2=0
cc_209 N_A_169_297#_M1004_g N_VGND_c_458_n 0.00431759f $X=2.14 $Y=0.56 $X2=0
+ $Y2=0
cc_210 N_A_169_297#_M1005_g N_VGND_c_458_n 0.00431683f $X=2.61 $Y=0.56 $X2=0
+ $Y2=0
cc_211 N_A_169_297#_M1006_g N_VGND_c_458_n 0.00431759f $X=3.08 $Y=0.56 $X2=0
+ $Y2=0
cc_212 N_A_169_297#_M1011_g N_VGND_c_458_n 0.00443737f $X=3.55 $Y=0.56 $X2=0
+ $Y2=0
cc_213 N_A_169_297#_M1012_g N_VGND_c_458_n 0.00522073f $X=4.07 $Y=0.56 $X2=0
+ $Y2=0
cc_214 N_A_169_297#_c_142_n N_VGND_c_458_n 0.0141066f $X=0.99 $Y=0.38 $X2=0
+ $Y2=0
cc_215 N_A_169_297#_c_125_n N_VGND_c_458_n 0.00764515f $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_216 N_VPWR_c_270_n N_X_M1003_s 0.00656398f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_217 N_VPWR_c_270_n N_X_M1010_s 0.00656398f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_c_270_n N_X_M1014_s 0.00656398f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_c_272_n N_X_c_359_n 0.0359797f $X=1.46 $Y=2 $X2=0 $Y2=0
cc_220 N_VPWR_c_273_n N_X_c_359_n 0.0470327f $X=2.4 $Y=2 $X2=0 $Y2=0
cc_221 N_VPWR_c_281_n N_X_c_359_n 0.0118139f $X=2.185 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_c_270_n N_X_c_359_n 0.00646998f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_223 N_VPWR_M1008_d N_X_c_355_n 0.00115412f $X=2.255 $Y=1.485 $X2=0 $Y2=0
cc_224 N_VPWR_c_273_n N_X_c_355_n 0.0107908f $X=2.4 $Y=2 $X2=0 $Y2=0
cc_225 N_VPWR_c_273_n N_X_c_377_n 0.0385613f $X=2.4 $Y=2 $X2=0 $Y2=0
cc_226 N_VPWR_c_274_n N_X_c_377_n 0.0470327f $X=3.34 $Y=2 $X2=0 $Y2=0
cc_227 N_VPWR_c_283_n N_X_c_377_n 0.0118139f $X=3.125 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_c_270_n N_X_c_377_n 0.00646998f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_274_n N_X_c_383_n 0.0385613f $X=3.34 $Y=2 $X2=0 $Y2=0
cc_230 N_VPWR_c_276_n N_X_c_383_n 0.0634568f $X=4.28 $Y=1.66 $X2=0 $Y2=0
cc_231 N_VPWR_c_285_n N_X_c_383_n 0.0118139f $X=4.065 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_c_270_n N_X_c_383_n 0.00646998f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_233 N_VPWR_M1008_d N_X_c_354_n 9.67171e-19 $X=2.255 $Y=1.485 $X2=0 $Y2=0
cc_234 N_VPWR_M1013_d N_X_c_354_n 0.00218693f $X=3.195 $Y=1.485 $X2=0 $Y2=0
cc_235 N_VPWR_c_273_n N_X_c_354_n 0.00707165f $X=2.4 $Y=2 $X2=0 $Y2=0
cc_236 N_VPWR_c_274_n N_X_c_354_n 0.0190013f $X=3.34 $Y=2 $X2=0 $Y2=0
cc_237 N_VPWR_c_276_n N_X_c_354_n 0.0107588f $X=4.28 $Y=1.66 $X2=0 $Y2=0
cc_238 N_VPWR_c_276_n N_VGND_c_448_n 0.0109366f $X=4.28 $Y=1.66 $X2=0 $Y2=0
cc_239 N_X_c_352_n N_VGND_M1004_d 0.00142274f $X=2.41 $Y=0.82 $X2=0 $Y2=0
cc_240 N_X_c_354_n N_VGND_M1004_d 7.35111e-19 $X=3.81 $Y=1.175 $X2=0 $Y2=0
cc_241 N_X_c_354_n N_VGND_M1006_d 0.00223254f $X=3.81 $Y=1.175 $X2=0 $Y2=0
cc_242 N_X_c_352_n N_VGND_c_445_n 0.0128838f $X=2.41 $Y=0.82 $X2=0 $Y2=0
cc_243 N_X_c_375_n N_VGND_c_445_n 0.0189749f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_244 N_X_c_354_n N_VGND_c_445_n 0.00821393f $X=3.81 $Y=1.175 $X2=0 $Y2=0
cc_245 N_X_c_380_n N_VGND_c_446_n 0.0189749f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_246 N_X_c_354_n N_VGND_c_446_n 0.0223861f $X=3.81 $Y=1.175 $X2=0 $Y2=0
cc_247 N_X_c_380_n N_VGND_c_448_n 0.0358347f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_248 N_X_c_354_n N_VGND_c_448_n 0.0124269f $X=3.81 $Y=1.175 $X2=0 $Y2=0
cc_249 N_X_c_358_n N_VGND_c_453_n 0.0115672f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_250 N_X_c_352_n N_VGND_c_453_n 0.00193763f $X=2.41 $Y=0.82 $X2=0 $Y2=0
cc_251 N_X_c_375_n N_VGND_c_455_n 0.0113207f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_252 N_X_c_354_n N_VGND_c_455_n 0.00494169f $X=3.81 $Y=1.175 $X2=0 $Y2=0
cc_253 N_X_c_380_n N_VGND_c_457_n 0.0115192f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_254 N_X_c_354_n N_VGND_c_457_n 0.00285443f $X=3.81 $Y=1.175 $X2=0 $Y2=0
cc_255 N_X_M1000_s N_VGND_c_458_n 0.00632385f $X=1.745 $Y=0.235 $X2=0 $Y2=0
cc_256 N_X_M1005_s N_VGND_c_458_n 0.00334789f $X=2.685 $Y=0.235 $X2=0 $Y2=0
cc_257 N_X_M1011_s N_VGND_c_458_n 0.00697884f $X=3.625 $Y=0.235 $X2=0 $Y2=0
cc_258 N_X_c_358_n N_VGND_c_458_n 0.0064623f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_259 N_X_c_352_n N_VGND_c_458_n 0.00470226f $X=2.41 $Y=0.82 $X2=0 $Y2=0
cc_260 N_X_c_375_n N_VGND_c_458_n 0.00641247f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_261 N_X_c_380_n N_VGND_c_458_n 0.00641247f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_262 N_X_c_354_n N_VGND_c_458_n 0.0175972f $X=3.81 $Y=1.175 $X2=0 $Y2=0
