* File: sky130_fd_sc_hdll__o21ba_1.pxi.spice
* Created: Thu Aug 27 19:19:34 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21BA_1%A_79_199# N_A_79_199#_M1009_s
+ N_A_79_199#_M1000_d N_A_79_199#_c_60_n N_A_79_199#_M1005_g N_A_79_199#_c_61_n
+ N_A_79_199#_M1007_g N_A_79_199#_c_65_n N_A_79_199#_c_106_p N_A_79_199#_c_62_n
+ N_A_79_199#_c_80_p N_A_79_199#_c_63_n N_A_79_199#_c_68_n N_A_79_199#_c_69_n
+ PM_SKY130_FD_SC_HDLL__O21BA_1%A_79_199#
x_PM_SKY130_FD_SC_HDLL__O21BA_1%B1_N N_B1_N_c_136_n N_B1_N_M1002_g
+ N_B1_N_c_137_n N_B1_N_M1001_g B1_N B1_N PM_SKY130_FD_SC_HDLL__O21BA_1%B1_N
x_PM_SKY130_FD_SC_HDLL__O21BA_1%A_222_93# N_A_222_93#_M1002_d
+ N_A_222_93#_M1001_d N_A_222_93#_c_170_n N_A_222_93#_M1000_g
+ N_A_222_93#_c_165_n N_A_222_93#_M1009_g N_A_222_93#_c_166_n
+ N_A_222_93#_c_167_n N_A_222_93#_c_173_n N_A_222_93#_c_168_n
+ N_A_222_93#_c_169_n PM_SKY130_FD_SC_HDLL__O21BA_1%A_222_93#
x_PM_SKY130_FD_SC_HDLL__O21BA_1%A2 N_A2_c_215_n N_A2_M1008_g N_A2_c_216_n
+ N_A2_M1004_g A2 A2 PM_SKY130_FD_SC_HDLL__O21BA_1%A2
x_PM_SKY130_FD_SC_HDLL__O21BA_1%A1 N_A1_c_243_n N_A1_M1003_g N_A1_c_244_n
+ N_A1_M1006_g A1 A1 PM_SKY130_FD_SC_HDLL__O21BA_1%A1
x_PM_SKY130_FD_SC_HDLL__O21BA_1%X N_X_M1007_s N_X_M1005_s N_X_c_262_n
+ N_X_c_264_n N_X_c_263_n X PM_SKY130_FD_SC_HDLL__O21BA_1%X
x_PM_SKY130_FD_SC_HDLL__O21BA_1%VPWR N_VPWR_M1005_d N_VPWR_M1000_s
+ N_VPWR_M1006_d N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n
+ VPWR N_VPWR_c_287_n N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_290_n
+ N_VPWR_c_291_n N_VPWR_c_282_n PM_SKY130_FD_SC_HDLL__O21BA_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O21BA_1%VGND N_VGND_M1007_d N_VGND_M1004_d
+ N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n VGND
+ N_VGND_c_334_n N_VGND_c_335_n N_VGND_c_336_n
+ PM_SKY130_FD_SC_HDLL__O21BA_1%VGND
x_PM_SKY130_FD_SC_HDLL__O21BA_1%A_460_47# N_A_460_47#_M1009_d
+ N_A_460_47#_M1003_d N_A_460_47#_c_376_n N_A_460_47#_c_373_n
+ N_A_460_47#_c_374_n N_A_460_47#_c_375_n
+ PM_SKY130_FD_SC_HDLL__O21BA_1%A_460_47#
cc_1 VNB N_A_79_199#_c_60_n 0.0285098f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A_79_199#_c_61_n 0.0223891f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_3 VNB N_A_79_199#_c_62_n 0.00195733f $X=-0.19 $Y=-0.24 $X2=1.975 $Y2=0.57
cc_4 VNB N_A_79_199#_c_63_n 0.00348049f $X=-0.19 $Y=-0.24 $X2=0.752 $Y2=1.16
cc_5 VNB N_B1_N_c_136_n 0.0216295f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.235
cc_6 VNB N_B1_N_c_137_n 0.0235766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB B1_N 0.00714238f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_A_222_93#_c_165_n 0.019846f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_9 VNB N_A_222_93#_c_166_n 0.0468258f $X=-0.19 $Y=-0.24 $X2=0.752 $Y2=1.325
cc_10 VNB N_A_222_93#_c_167_n 0.0131694f $X=-0.19 $Y=-0.24 $X2=0.752 $Y2=1.865
cc_11 VNB N_A_222_93#_c_168_n 0.00322048f $X=-0.19 $Y=-0.24 $X2=2.432 $Y2=2.3
cc_12 VNB N_A_222_93#_c_169_n 0.0123648f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_13 VNB N_A2_c_215_n 0.0202073f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.235
cc_14 VNB N_A2_c_216_n 0.0167691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB A2 0.00827309f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_16 VNB N_A1_c_243_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.235
cc_17 VNB N_A1_c_244_n 0.027445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB A1 0.0170438f $X=-0.19 $Y=-0.24 $X2=1.89 $Y2=1.95
cc_19 VNB N_X_c_262_n 0.0172248f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_20 VNB N_X_c_263_n 0.0242325f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.95
cc_21 VNB N_VPWR_c_282_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_330_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_23 VNB N_VGND_c_331_n 0.00471543f $X=-0.19 $Y=-0.24 $X2=1.89 $Y2=1.95
cc_24 VNB N_VGND_c_332_n 0.0549554f $X=-0.19 $Y=-0.24 $X2=1.975 $Y2=0.57
cc_25 VNB N_VGND_c_333_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=1.975 $Y2=0.57
cc_26 VNB N_VGND_c_334_n 0.0199212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_335_n 0.222409f $X=-0.19 $Y=-0.24 $X2=1.975 $Y2=1.745
cc_28 VNB N_VGND_c_336_n 0.0245951f $X=-0.19 $Y=-0.24 $X2=2.445 $Y2=1.745
cc_29 VNB N_A_460_47#_c_373_n 0.0170716f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_30 VNB N_A_460_47#_c_374_n 0.00256037f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_31 VNB N_A_460_47#_c_375_n 0.0181301f $X=-0.19 $Y=-0.24 $X2=1.89 $Y2=1.95
cc_32 VPB N_A_79_199#_c_60_n 0.0347953f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_33 VPB N_A_79_199#_c_65_n 0.00301754f $X=-0.19 $Y=1.305 $X2=0.752 $Y2=1.865
cc_34 VPB N_A_79_199#_c_62_n 0.0028515f $X=-0.19 $Y=1.305 $X2=1.975 $Y2=0.57
cc_35 VPB N_A_79_199#_c_63_n 4.80651e-19 $X=-0.19 $Y=1.305 $X2=0.752 $Y2=1.16
cc_36 VPB N_A_79_199#_c_68_n 0.0156878f $X=-0.19 $Y=1.305 $X2=1.89 $Y2=1.745
cc_37 VPB N_A_79_199#_c_69_n 0.00401354f $X=-0.19 $Y=1.305 $X2=2.445 $Y2=1.62
cc_38 VPB N_B1_N_c_137_n 0.0302624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB B1_N 0.00226922f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_40 VPB N_A_222_93#_c_170_n 0.0193484f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_41 VPB N_A_222_93#_c_166_n 0.0187712f $X=-0.19 $Y=1.305 $X2=0.752 $Y2=1.325
cc_42 VPB N_A_222_93#_c_167_n 0.00655548f $X=-0.19 $Y=1.305 $X2=0.752 $Y2=1.865
cc_43 VPB N_A_222_93#_c_173_n 0.00804367f $X=-0.19 $Y=1.305 $X2=1.89 $Y2=1.95
cc_44 VPB N_A_222_93#_c_168_n 0.00377215f $X=-0.19 $Y=1.305 $X2=2.432 $Y2=2.3
cc_45 VPB N_A2_c_215_n 0.0256007f $X=-0.19 $Y=1.305 $X2=1.85 $Y2=0.235
cc_46 VPB N_A1_c_244_n 0.0321628f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_X_c_264_n 0.00759142f $X=-0.19 $Y=1.305 $X2=1.89 $Y2=1.95
cc_48 VPB N_X_c_263_n 0.00838059f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.95
cc_49 VPB X 0.0322798f $X=-0.19 $Y=1.305 $X2=1.975 $Y2=1.455
cc_50 VPB N_VPWR_c_283_n 0.0188196f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.56
cc_51 VPB N_VPWR_c_284_n 0.0163315f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.95
cc_52 VPB N_VPWR_c_285_n 0.0121516f $X=-0.19 $Y=1.305 $X2=1.975 $Y2=0.57
cc_53 VPB N_VPWR_c_286_n 0.0396463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_287_n 0.0177751f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_55 VPB N_VPWR_c_288_n 0.0212115f $X=-0.19 $Y=1.305 $X2=1.975 $Y2=1.745
cc_56 VPB N_VPWR_c_289_n 0.0292293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_290_n 0.00785178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_291_n 0.00631679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_282_n 0.0539226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 N_A_79_199#_c_61_n N_B1_N_c_136_n 0.0144197f $X=0.55 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_61 N_A_79_199#_c_60_n N_B1_N_c_137_n 0.0348729f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_62 N_A_79_199#_c_65_n N_B1_N_c_137_n 0.0105947f $X=0.752 $Y=1.865 $X2=0 $Y2=0
cc_63 N_A_79_199#_c_63_n N_B1_N_c_137_n 0.00222541f $X=0.752 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_79_199#_c_68_n N_B1_N_c_137_n 0.0162558f $X=1.89 $Y=1.745 $X2=0 $Y2=0
cc_65 N_A_79_199#_c_60_n B1_N 2.89974e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_79_199#_c_63_n B1_N 0.0263171f $X=0.752 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_79_199#_c_68_n B1_N 0.00122077f $X=1.89 $Y=1.745 $X2=0 $Y2=0
cc_68 N_A_79_199#_c_68_n N_A_222_93#_M1001_d 0.00265291f $X=1.89 $Y=1.745 $X2=0
+ $Y2=0
cc_69 N_A_79_199#_c_62_n N_A_222_93#_c_170_n 0.0017729f $X=1.975 $Y=0.57 $X2=0
+ $Y2=0
cc_70 N_A_79_199#_c_80_p N_A_222_93#_c_170_n 0.0103214f $X=2.445 $Y=2.3 $X2=0
+ $Y2=0
cc_71 N_A_79_199#_c_69_n N_A_222_93#_c_170_n 0.0328633f $X=2.445 $Y=1.62 $X2=0
+ $Y2=0
cc_72 N_A_79_199#_c_62_n N_A_222_93#_c_165_n 0.0102549f $X=1.975 $Y=0.57 $X2=0
+ $Y2=0
cc_73 N_A_79_199#_c_62_n N_A_222_93#_c_166_n 0.0212186f $X=1.975 $Y=0.57 $X2=0
+ $Y2=0
cc_74 N_A_79_199#_c_68_n N_A_222_93#_c_166_n 0.00495661f $X=1.89 $Y=1.745 $X2=0
+ $Y2=0
cc_75 N_A_79_199#_c_69_n N_A_222_93#_c_166_n 0.00278379f $X=2.445 $Y=1.62 $X2=0
+ $Y2=0
cc_76 N_A_79_199#_c_62_n N_A_222_93#_c_167_n 0.00346625f $X=1.975 $Y=0.57 $X2=0
+ $Y2=0
cc_77 N_A_79_199#_c_69_n N_A_222_93#_c_167_n 8.22352e-19 $X=2.445 $Y=1.62 $X2=0
+ $Y2=0
cc_78 N_A_79_199#_c_65_n N_A_222_93#_c_173_n 0.0111419f $X=0.752 $Y=1.865 $X2=0
+ $Y2=0
cc_79 N_A_79_199#_c_68_n N_A_222_93#_c_173_n 0.0445768f $X=1.89 $Y=1.745 $X2=0
+ $Y2=0
cc_80 N_A_79_199#_c_69_n N_A_222_93#_c_173_n 0.0155901f $X=2.445 $Y=1.62 $X2=0
+ $Y2=0
cc_81 N_A_79_199#_c_62_n N_A_222_93#_c_168_n 0.0448396f $X=1.975 $Y=0.57 $X2=0
+ $Y2=0
cc_82 N_A_79_199#_c_69_n N_A_222_93#_c_168_n 0.00572925f $X=2.445 $Y=1.62 $X2=0
+ $Y2=0
cc_83 N_A_79_199#_c_62_n N_A_222_93#_c_169_n 0.02043f $X=1.975 $Y=0.57 $X2=0
+ $Y2=0
cc_84 N_A_79_199#_c_62_n N_A2_c_215_n 6.39012e-19 $X=1.975 $Y=0.57 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_79_199#_c_69_n N_A2_c_215_n 0.00279562f $X=2.445 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_79_199#_c_62_n A2 0.0157222f $X=1.975 $Y=0.57 $X2=0 $Y2=0
cc_87 N_A_79_199#_c_69_n A2 0.0290673f $X=2.445 $Y=1.62 $X2=0 $Y2=0
cc_88 N_A_79_199#_c_60_n N_X_c_262_n 0.00135005f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_79_199#_c_60_n N_X_c_264_n 0.002856f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_79_199#_c_65_n N_X_c_264_n 0.0237219f $X=0.752 $Y=1.865 $X2=0 $Y2=0
cc_91 N_A_79_199#_c_60_n N_X_c_263_n 0.0125168f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_79_199#_c_61_n N_X_c_263_n 0.00578113f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_79_199#_c_65_n N_X_c_263_n 0.00812237f $X=0.752 $Y=1.865 $X2=0 $Y2=0
cc_94 N_A_79_199#_c_63_n N_X_c_263_n 0.0256678f $X=0.752 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_79_199#_c_60_n X 0.0149429f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_79_199#_c_106_p X 0.0115315f $X=0.86 $Y=1.95 $X2=0 $Y2=0
cc_97 N_A_79_199#_c_65_n N_VPWR_M1005_d 0.0109535f $X=0.752 $Y=1.865 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A_79_199#_c_106_p N_VPWR_M1005_d 0.00524855f $X=0.86 $Y=1.95 $X2=-0.19
+ $Y2=-0.24
cc_99 N_A_79_199#_c_68_n N_VPWR_M1005_d 0.00223163f $X=1.89 $Y=1.745 $X2=-0.19
+ $Y2=-0.24
cc_100 N_A_79_199#_c_68_n N_VPWR_M1000_s 0.00282833f $X=1.89 $Y=1.745 $X2=0
+ $Y2=0
cc_101 N_A_79_199#_c_69_n N_VPWR_M1000_s 0.0129734f $X=2.445 $Y=1.62 $X2=0 $Y2=0
cc_102 N_A_79_199#_c_60_n N_VPWR_c_283_n 0.00503427f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_103 N_A_79_199#_c_106_p N_VPWR_c_283_n 0.0183673f $X=0.86 $Y=1.95 $X2=0 $Y2=0
cc_104 N_A_79_199#_c_68_n N_VPWR_c_283_n 0.0113507f $X=1.89 $Y=1.745 $X2=0 $Y2=0
cc_105 N_A_79_199#_c_68_n N_VPWR_c_284_n 0.0218908f $X=1.89 $Y=1.745 $X2=0 $Y2=0
cc_106 N_A_79_199#_c_60_n N_VPWR_c_287_n 0.00673617f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_107 N_A_79_199#_c_68_n N_VPWR_c_288_n 0.0123218f $X=1.89 $Y=1.745 $X2=0 $Y2=0
cc_108 N_A_79_199#_c_80_p N_VPWR_c_289_n 0.0170491f $X=2.445 $Y=2.3 $X2=0 $Y2=0
cc_109 N_A_79_199#_c_69_n N_VPWR_c_289_n 0.0027968f $X=2.445 $Y=1.62 $X2=0 $Y2=0
cc_110 N_A_79_199#_M1000_d N_VPWR_c_282_n 0.00235276f $X=2.29 $Y=1.485 $X2=0
+ $Y2=0
cc_111 N_A_79_199#_c_60_n N_VPWR_c_282_n 0.0139121f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_79_199#_c_106_p N_VPWR_c_282_n 9.92431e-19 $X=0.86 $Y=1.95 $X2=0
+ $Y2=0
cc_113 N_A_79_199#_c_80_p N_VPWR_c_282_n 0.0114213f $X=2.445 $Y=2.3 $X2=0 $Y2=0
cc_114 N_A_79_199#_c_68_n N_VPWR_c_282_n 0.0228085f $X=1.89 $Y=1.745 $X2=0 $Y2=0
cc_115 N_A_79_199#_c_69_n N_VPWR_c_282_n 0.00432231f $X=2.445 $Y=1.62 $X2=0
+ $Y2=0
cc_116 N_A_79_199#_c_60_n N_VGND_c_330_n 0.00123968f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_117 N_A_79_199#_c_61_n N_VGND_c_330_n 0.00694531f $X=0.55 $Y=0.995 $X2=0
+ $Y2=0
cc_118 N_A_79_199#_c_63_n N_VGND_c_330_n 0.0140728f $X=0.752 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_79_199#_c_62_n N_VGND_c_332_n 0.0118139f $X=1.975 $Y=0.57 $X2=0 $Y2=0
cc_120 N_A_79_199#_M1009_s N_VGND_c_335_n 0.00701161f $X=1.85 $Y=0.235 $X2=0
+ $Y2=0
cc_121 N_A_79_199#_c_61_n N_VGND_c_335_n 0.0131276f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_79_199#_c_62_n N_VGND_c_335_n 0.00646998f $X=1.975 $Y=0.57 $X2=0
+ $Y2=0
cc_123 N_A_79_199#_c_61_n N_VGND_c_336_n 0.00585385f $X=0.55 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_A_79_199#_c_62_n N_A_460_47#_c_376_n 0.0290299f $X=1.975 $Y=0.57 $X2=0
+ $Y2=0
cc_125 N_A_79_199#_c_62_n N_A_460_47#_c_374_n 0.0109673f $X=1.975 $Y=0.57 $X2=0
+ $Y2=0
cc_126 N_B1_N_c_137_n N_A_222_93#_c_166_n 0.0193112f $X=1.06 $Y=1.41 $X2=0 $Y2=0
cc_127 B1_N N_A_222_93#_c_166_n 0.00240381f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_128 N_B1_N_c_137_n N_A_222_93#_c_173_n 0.00536327f $X=1.06 $Y=1.41 $X2=0
+ $Y2=0
cc_129 B1_N N_A_222_93#_c_173_n 0.0182918f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_130 N_B1_N_c_136_n N_A_222_93#_c_168_n 0.0039709f $X=1.035 $Y=0.995 $X2=0
+ $Y2=0
cc_131 N_B1_N_c_137_n N_A_222_93#_c_168_n 0.00526795f $X=1.06 $Y=1.41 $X2=0
+ $Y2=0
cc_132 B1_N N_A_222_93#_c_168_n 0.0250383f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_133 N_B1_N_c_136_n N_A_222_93#_c_169_n 0.00238949f $X=1.035 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_B1_N_c_137_n N_A_222_93#_c_169_n 4.49744e-19 $X=1.06 $Y=1.41 $X2=0
+ $Y2=0
cc_135 B1_N N_A_222_93#_c_169_n 0.0138303f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_136 N_B1_N_c_137_n N_VPWR_c_283_n 9.21934e-19 $X=1.06 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B1_N_c_137_n N_VPWR_c_288_n 0.00250363f $X=1.06 $Y=1.41 $X2=0 $Y2=0
cc_138 N_B1_N_c_137_n N_VPWR_c_282_n 0.00406356f $X=1.06 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B1_N_c_136_n N_VGND_c_330_n 0.00606311f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B1_N_c_136_n N_VGND_c_332_n 0.00510437f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B1_N_c_136_n N_VGND_c_335_n 0.00512902f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_222_93#_c_170_n N_A2_c_215_n 0.00917729f $X=2.2 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_143 N_A_222_93#_c_167_n N_A2_c_215_n 0.0267053f $X=2.2 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_144 N_A_222_93#_c_165_n N_A2_c_216_n 0.00969055f $X=2.225 $Y=0.995 $X2=0
+ $Y2=0
cc_145 N_A_222_93#_c_167_n A2 0.00973885f $X=2.2 $Y=1.202 $X2=0 $Y2=0
cc_146 N_A_222_93#_c_170_n N_VPWR_c_284_n 0.00496378f $X=2.2 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_222_93#_c_170_n N_VPWR_c_289_n 0.00514296f $X=2.2 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_222_93#_c_170_n N_VPWR_c_282_n 0.00796532f $X=2.2 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_222_93#_c_169_n N_VGND_c_330_n 0.0162021f $X=1.295 $Y=0.66 $X2=0
+ $Y2=0
cc_150 N_A_222_93#_c_165_n N_VGND_c_332_n 0.0055654f $X=2.225 $Y=0.995 $X2=0
+ $Y2=0
cc_151 N_A_222_93#_c_169_n N_VGND_c_332_n 0.0114543f $X=1.295 $Y=0.66 $X2=0
+ $Y2=0
cc_152 N_A_222_93#_c_165_n N_VGND_c_335_n 0.0116149f $X=2.225 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_222_93#_c_169_n N_VGND_c_335_n 0.0154915f $X=1.295 $Y=0.66 $X2=0
+ $Y2=0
cc_154 N_A_222_93#_c_165_n N_A_460_47#_c_376_n 0.00571573f $X=2.225 $Y=0.995
+ $X2=0 $Y2=0
cc_155 N_A_222_93#_c_165_n N_A_460_47#_c_374_n 0.00251094f $X=2.225 $Y=0.995
+ $X2=0 $Y2=0
cc_156 N_A2_c_216_n N_A1_c_243_n 0.0237539f $X=2.705 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_157 N_A2_c_215_n N_A1_c_244_n 0.0743723f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_158 A2 N_A1_c_244_n 7.46909e-19 $X=2.515 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A2_c_215_n A1 6.65775e-19 $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_160 A2 A1 0.019043f $X=2.515 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A2_c_215_n N_VPWR_c_286_n 0.00413089f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A2_c_215_n N_VPWR_c_289_n 0.00702461f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A2_c_215_n N_VPWR_c_282_n 0.0127602f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A2_c_216_n N_VGND_c_331_n 0.00268723f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A2_c_216_n N_VGND_c_332_n 0.00439206f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A2_c_216_n N_VGND_c_335_n 0.0061063f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A2_c_215_n N_A_460_47#_c_373_n 5.76324e-19 $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A2_c_216_n N_A_460_47#_c_373_n 0.0103662f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_169 A2 N_A_460_47#_c_373_n 0.0171072f $X=2.515 $Y=1.105 $X2=0 $Y2=0
cc_170 N_A2_c_215_n N_A_460_47#_c_374_n 0.00265731f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_171 A2 N_A_460_47#_c_374_n 0.0276188f $X=2.515 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A1_c_244_n N_VPWR_c_286_n 0.0308786f $X=3.15 $Y=1.41 $X2=0 $Y2=0
cc_173 A1 N_VPWR_c_286_n 0.0213068f $X=3.37 $Y=1.19 $X2=0 $Y2=0
cc_174 N_A1_c_244_n N_VPWR_c_289_n 0.00427505f $X=3.15 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A1_c_244_n N_VPWR_c_282_n 0.00743383f $X=3.15 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A1_c_243_n N_VGND_c_331_n 0.00268723f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A1_c_243_n N_VGND_c_334_n 0.00439206f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A1_c_243_n N_VGND_c_335_n 0.00704893f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A1_c_243_n N_A_460_47#_c_373_n 0.0137032f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A1_c_244_n N_A_460_47#_c_373_n 0.00321782f $X=3.15 $Y=1.41 $X2=0 $Y2=0
cc_181 A1 N_A_460_47#_c_373_n 0.0429268f $X=3.37 $Y=1.19 $X2=0 $Y2=0
cc_182 X N_VPWR_c_287_n 0.0217765f $X=0.145 $Y=2.125 $X2=0 $Y2=0
cc_183 N_X_M1005_s N_VPWR_c_282_n 0.00217517f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_184 X N_VPWR_c_282_n 0.0128576f $X=0.145 $Y=2.125 $X2=0 $Y2=0
cc_185 N_X_M1007_s N_VGND_c_335_n 0.00346044f $X=0.215 $Y=0.235 $X2=0 $Y2=0
cc_186 N_X_c_262_n N_VGND_c_335_n 0.0122067f $X=0.34 $Y=0.66 $X2=0 $Y2=0
cc_187 N_X_c_262_n N_VGND_c_336_n 0.0106755f $X=0.34 $Y=0.66 $X2=0 $Y2=0
cc_188 N_VPWR_c_282_n A_554_297# 0.0123962f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_189 N_VGND_c_335_n N_A_460_47#_M1009_d 0.00272306f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_190 N_VGND_c_335_n N_A_460_47#_M1003_d 0.00285244f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_191 N_VGND_c_332_n N_A_460_47#_c_376_n 0.0196975f $X=2.83 $Y=0 $X2=0 $Y2=0
cc_192 N_VGND_c_335_n N_A_460_47#_c_376_n 0.0124576f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_193 N_VGND_M1004_d N_A_460_47#_c_373_n 0.00165819f $X=2.78 $Y=0.235 $X2=0
+ $Y2=0
cc_194 N_VGND_c_331_n N_A_460_47#_c_373_n 0.0116529f $X=2.915 $Y=0.39 $X2=0
+ $Y2=0
cc_195 N_VGND_c_332_n N_A_460_47#_c_373_n 0.00248202f $X=2.83 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_c_334_n N_A_460_47#_c_373_n 0.00260097f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_197 N_VGND_c_335_n N_A_460_47#_c_373_n 0.0109399f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_334_n N_A_460_47#_c_375_n 0.020323f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_335_n N_A_460_47#_c_375_n 0.0125178f $X=3.45 $Y=0 $X2=0 $Y2=0
