* File: sky130_fd_sc_hdll__muxb8to1_4.pxi.spice
* Created: Wed Sep  2 08:36:14 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[0] N_S[0]_c_904_n N_S[0]_c_905_n
+ N_S[0]_M1001_g N_S[0]_c_906_n N_S[0]_M1043_g N_S[0]_c_907_n N_S[0]_c_908_n
+ N_S[0]_M1067_g N_S[0]_c_909_n N_S[0]_c_929_n N_S[0]_M1040_g N_S[0]_c_910_n
+ N_S[0]_c_911_n N_S[0]_c_912_n N_S[0]_c_913_n N_S[0]_c_914_n N_S[0]_M1003_g
+ N_S[0]_c_915_n N_S[0]_c_916_n N_S[0]_M1100_g N_S[0]_c_917_n N_S[0]_c_918_n
+ N_S[0]_M1109_g N_S[0]_c_919_n N_S[0]_c_920_n N_S[0]_M1133_g N_S[0]_c_921_n
+ N_S[0]_c_922_n N_S[0]_c_923_n N_S[0]_c_924_n S[0] N_S[0]_c_925_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[0]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[1] N_S[1]_c_1016_n N_S[1]_c_1038_n
+ N_S[1]_M1052_g N_S[1]_c_1017_n N_S[1]_M1084_g N_S[1]_c_1018_n N_S[1]_c_1040_n
+ N_S[1]_c_1019_n N_S[1]_c_1020_n N_S[1]_M1138_g N_S[1]_c_1042_n N_S[1]_M1088_g
+ N_S[1]_c_1021_n N_S[1]_c_1022_n N_S[1]_c_1023_n N_S[1]_c_1024_n
+ N_S[1]_c_1025_n N_S[1]_M1029_g N_S[1]_c_1026_n N_S[1]_c_1027_n N_S[1]_M1058_g
+ N_S[1]_c_1028_n N_S[1]_c_1029_n N_S[1]_M1083_g N_S[1]_c_1030_n N_S[1]_c_1031_n
+ N_S[1]_M1102_g N_S[1]_c_1032_n N_S[1]_c_1033_n N_S[1]_c_1034_n N_S[1]_c_1035_n
+ S[1] N_S[1]_c_1036_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[1]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_142_325# N_A_142_325#_M1043_s
+ N_A_142_325#_M1001_s N_A_142_325#_c_1141_n N_A_142_325#_M1010_g
+ N_A_142_325#_c_1142_n N_A_142_325#_c_1134_n N_A_142_325#_c_1144_n
+ N_A_142_325#_M1019_g N_A_142_325#_c_1145_n N_A_142_325#_c_1146_n
+ N_A_142_325#_M1051_g N_A_142_325#_c_1147_n N_A_142_325#_c_1148_n
+ N_A_142_325#_M1147_g N_A_142_325#_c_1149_n N_A_142_325#_c_1150_n
+ N_A_142_325#_c_1151_n N_A_142_325#_c_1135_n N_A_142_325#_c_1136_n
+ N_A_142_325#_c_1137_n N_A_142_325#_c_1153_n N_A_142_325#_c_1138_n
+ N_A_142_325#_c_1139_n N_A_142_325#_c_1140_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_142_325#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_142_599# N_A_142_599#_M1084_d
+ N_A_142_599#_M1052_s N_A_142_599#_c_1253_n N_A_142_599#_M1054_g
+ N_A_142_599#_c_1254_n N_A_142_599#_c_1246_n N_A_142_599#_c_1256_n
+ N_A_142_599#_M1080_g N_A_142_599#_c_1257_n N_A_142_599#_c_1258_n
+ N_A_142_599#_M1092_g N_A_142_599#_c_1259_n N_A_142_599#_c_1260_n
+ N_A_142_599#_M1123_g N_A_142_599#_c_1261_n N_A_142_599#_c_1262_n
+ N_A_142_599#_c_1263_n N_A_142_599#_c_1247_n N_A_142_599#_c_1248_n
+ N_A_142_599#_c_1264_n N_A_142_599#_c_1249_n N_A_142_599#_c_1266_n
+ N_A_142_599#_c_1250_n N_A_142_599#_c_1251_n N_A_142_599#_c_1252_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_142_599#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[0] N_D[0]_M1012_g N_D[0]_M1065_g
+ N_D[0]_M1097_g N_D[0]_M1049_g N_D[0]_M1086_g N_D[0]_M1151_g N_D[0]_M1156_g
+ N_D[0]_M1137_g D[0] N_D[0]_c_1372_n N_D[0]_c_1373_n N_D[0]_c_1374_n
+ N_D[0]_c_1375_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[0]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[1] N_D[1]_M1017_g N_D[1]_M1030_g
+ N_D[1]_M1059_g N_D[1]_M1055_g N_D[1]_M1093_g N_D[1]_M1068_g N_D[1]_M1157_g
+ N_D[1]_M1141_g D[1] N_D[1]_c_1471_n N_D[1]_c_1472_n N_D[1]_c_1473_n
+ N_D[1]_c_1474_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[1]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[2] N_D[2]_M1071_g N_D[2]_M1013_g
+ N_D[2]_M1037_g N_D[2]_M1090_g N_D[2]_M1118_g N_D[2]_M1069_g N_D[2]_M1150_g
+ N_D[2]_M1158_g D[2] N_D[2]_c_1568_n N_D[2]_c_1569_n N_D[2]_c_1570_n
+ N_D[2]_c_1571_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[2]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[3] N_D[3]_M1000_g N_D[3]_M1015_g
+ N_D[3]_M1047_g N_D[3]_M1076_g N_D[3]_M1095_g N_D[3]_M1104_g N_D[3]_M1136_g
+ N_D[3]_M1120_g D[3] N_D[3]_c_1669_n N_D[3]_c_1670_n N_D[3]_c_1671_n
+ N_D[3]_c_1672_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[3]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1755_265# N_A_1755_265#_M1094_s
+ N_A_1755_265#_M1072_s N_A_1755_265#_c_1765_n N_A_1755_265#_M1050_g
+ N_A_1755_265#_c_1766_n N_A_1755_265#_c_1767_n N_A_1755_265#_c_1768_n
+ N_A_1755_265#_M1073_g N_A_1755_265#_c_1769_n N_A_1755_265#_c_1770_n
+ N_A_1755_265#_M1116_g N_A_1755_265#_c_1771_n N_A_1755_265#_c_1772_n
+ N_A_1755_265#_M1126_g N_A_1755_265#_c_1773_n N_A_1755_265#_c_1774_n
+ N_A_1755_265#_c_1758_n N_A_1755_265#_c_1759_n N_A_1755_265#_c_1760_n
+ N_A_1755_265#_c_1761_n N_A_1755_265#_c_1777_n N_A_1755_265#_c_1762_n
+ N_A_1755_265#_c_1763_n N_A_1755_265#_c_1779_n N_A_1755_265#_c_1764_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1755_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1755_793# N_A_1755_793#_M1060_s
+ N_A_1755_793#_M1007_d N_A_1755_793#_c_1884_n N_A_1755_793#_M1031_g
+ N_A_1755_793#_c_1885_n N_A_1755_793#_c_1886_n N_A_1755_793#_c_1887_n
+ N_A_1755_793#_M1036_g N_A_1755_793#_c_1888_n N_A_1755_793#_c_1889_n
+ N_A_1755_793#_M1124_g N_A_1755_793#_c_1890_n N_A_1755_793#_c_1891_n
+ N_A_1755_793#_M1152_g N_A_1755_793#_c_1892_n N_A_1755_793#_c_1893_n
+ N_A_1755_793#_c_1877_n N_A_1755_793#_c_1878_n N_A_1755_793#_c_1896_n
+ N_A_1755_793#_c_1897_n N_A_1755_793#_c_1879_n N_A_1755_793#_c_1880_n
+ N_A_1755_793#_c_1898_n N_A_1755_793#_c_1881_n N_A_1755_793#_c_1882_n
+ N_A_1755_793#_c_1883_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1755_793#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[2] N_S[2]_c_2002_n N_S[2]_M1024_g
+ N_S[2]_c_2003_n N_S[2]_c_2004_n N_S[2]_c_2005_n N_S[2]_M1028_g N_S[2]_c_2006_n
+ N_S[2]_c_2007_n N_S[2]_M1044_g N_S[2]_c_2008_n N_S[2]_c_2009_n N_S[2]_M1057_g
+ N_S[2]_c_2010_n N_S[2]_c_2011_n N_S[2]_c_2012_n N_S[2]_c_2013_n
+ N_S[2]_c_2014_n N_S[2]_c_2025_n N_S[2]_M1072_g N_S[2]_c_2015_n N_S[2]_M1094_g
+ N_S[2]_c_2016_n N_S[2]_c_2017_n N_S[2]_M1103_g N_S[2]_c_2018_n N_S[2]_M1115_g
+ N_S[2]_c_2019_n N_S[2]_c_2020_n N_S[2]_c_2021_n N_S[2]_c_2022_n S[2]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[2]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[3] N_S[3]_c_2119_n N_S[3]_M1016_g
+ N_S[3]_c_2120_n N_S[3]_c_2121_n N_S[3]_c_2122_n N_S[3]_M1020_g N_S[3]_c_2123_n
+ N_S[3]_c_2124_n N_S[3]_M1048_g N_S[3]_c_2125_n N_S[3]_c_2126_n N_S[3]_M1135_g
+ N_S[3]_c_2127_n N_S[3]_c_2128_n N_S[3]_c_2129_n N_S[3]_c_2130_n
+ N_S[3]_c_2140_n N_S[3]_c_2131_n N_S[3]_c_2142_n N_S[3]_M1007_g N_S[3]_c_2132_n
+ N_S[3]_M1060_g N_S[3]_c_2133_n N_S[3]_c_2134_n N_S[3]_M1140_g N_S[3]_c_2144_n
+ N_S[3]_M1125_g N_S[3]_c_2135_n N_S[3]_c_2136_n N_S[3]_c_2137_n N_S[3]_c_2138_n
+ S[3] PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[3]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[4] N_S[4]_c_2244_n N_S[4]_c_2245_n
+ N_S[4]_M1128_g N_S[4]_c_2246_n N_S[4]_M1121_g N_S[4]_c_2247_n N_S[4]_c_2248_n
+ N_S[4]_M1129_g N_S[4]_c_2249_n N_S[4]_c_2269_n N_S[4]_M1155_g N_S[4]_c_2250_n
+ N_S[4]_c_2251_n N_S[4]_c_2252_n N_S[4]_c_2253_n N_S[4]_c_2254_n N_S[4]_M1006_g
+ N_S[4]_c_2255_n N_S[4]_c_2256_n N_S[4]_M1022_g N_S[4]_c_2257_n N_S[4]_c_2258_n
+ N_S[4]_M1035_g N_S[4]_c_2259_n N_S[4]_c_2260_n N_S[4]_M1066_g N_S[4]_c_2261_n
+ N_S[4]_c_2262_n N_S[4]_c_2263_n N_S[4]_c_2264_n S[4] N_S[4]_c_2265_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[4]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[5] N_S[5]_c_2364_n N_S[5]_c_2386_n
+ N_S[5]_M1018_g N_S[5]_c_2365_n N_S[5]_M1074_g N_S[5]_c_2366_n N_S[5]_c_2388_n
+ N_S[5]_c_2367_n N_S[5]_c_2368_n N_S[5]_M1154_g N_S[5]_c_2390_n N_S[5]_M1039_g
+ N_S[5]_c_2369_n N_S[5]_c_2370_n N_S[5]_c_2371_n N_S[5]_c_2372_n
+ N_S[5]_c_2373_n N_S[5]_M1009_g N_S[5]_c_2374_n N_S[5]_c_2375_n N_S[5]_M1038_g
+ N_S[5]_c_2376_n N_S[5]_c_2377_n N_S[5]_M1112_g N_S[5]_c_2378_n N_S[5]_c_2379_n
+ N_S[5]_M1142_g N_S[5]_c_2380_n N_S[5]_c_2381_n N_S[5]_c_2382_n N_S[5]_c_2383_n
+ S[5] N_S[5]_c_2384_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[5]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2626_325# N_A_2626_325#_M1121_s
+ N_A_2626_325#_M1128_s N_A_2626_325#_c_2499_n N_A_2626_325#_M1004_g
+ N_A_2626_325#_c_2500_n N_A_2626_325#_c_2492_n N_A_2626_325#_c_2502_n
+ N_A_2626_325#_M1110_g N_A_2626_325#_c_2503_n N_A_2626_325#_c_2504_n
+ N_A_2626_325#_M1131_g N_A_2626_325#_c_2505_n N_A_2626_325#_c_2506_n
+ N_A_2626_325#_M1146_g N_A_2626_325#_c_2507_n N_A_2626_325#_c_2508_n
+ N_A_2626_325#_c_2509_n N_A_2626_325#_c_2493_n N_A_2626_325#_c_2494_n
+ N_A_2626_325#_c_2495_n N_A_2626_325#_c_2511_n N_A_2626_325#_c_2496_n
+ N_A_2626_325#_c_2497_n N_A_2626_325#_c_2498_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2626_325#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2626_599# N_A_2626_599#_M1074_s
+ N_A_2626_599#_M1018_s N_A_2626_599#_c_2615_n N_A_2626_599#_M1021_g
+ N_A_2626_599#_c_2616_n N_A_2626_599#_c_2608_n N_A_2626_599#_c_2618_n
+ N_A_2626_599#_M1041_g N_A_2626_599#_c_2619_n N_A_2626_599#_c_2620_n
+ N_A_2626_599#_M1056_g N_A_2626_599#_c_2621_n N_A_2626_599#_c_2622_n
+ N_A_2626_599#_M1078_g N_A_2626_599#_c_2623_n N_A_2626_599#_c_2624_n
+ N_A_2626_599#_c_2625_n N_A_2626_599#_c_2609_n N_A_2626_599#_c_2610_n
+ N_A_2626_599#_c_2626_n N_A_2626_599#_c_2611_n N_A_2626_599#_c_2628_n
+ N_A_2626_599#_c_2612_n N_A_2626_599#_c_2613_n N_A_2626_599#_c_2614_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2626_599#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[4] N_D[4]_M1042_g N_D[4]_M1027_g
+ N_D[4]_M1034_g N_D[4]_M1062_g N_D[4]_M1105_g N_D[4]_M1045_g N_D[4]_M1079_g
+ N_D[4]_M1127_g D[4] N_D[4]_c_2738_n N_D[4]_c_2739_n N_D[4]_c_2740_n
+ N_D[4]_c_2741_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[4]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[5] N_D[5]_M1046_g N_D[5]_M1033_g
+ N_D[5]_M1077_g N_D[5]_M1070_g N_D[5]_M1113_g N_D[5]_M1106_g N_D[5]_M1107_g
+ N_D[5]_M1134_g D[5] N_D[5]_c_2837_n N_D[5]_c_2838_n N_D[5]_c_2839_n
+ N_D[5]_c_2840_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[5]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[6] N_D[6]_M1082_g N_D[6]_M1005_g
+ N_D[6]_M1081_g N_D[6]_M1108_g N_D[6]_M1130_g N_D[6]_M1111_g N_D[6]_M1159_g
+ N_D[6]_M1145_g D[6] N_D[6]_c_2934_n N_D[6]_c_2935_n N_D[6]_c_2936_n
+ N_D[6]_c_2937_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[6]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[7] N_D[7]_M1087_g N_D[7]_M1014_g
+ N_D[7]_M1025_g N_D[7]_M1117_g N_D[7]_M1139_g N_D[7]_M1026_g N_D[7]_M1098_g
+ N_D[7]_M1153_g D[7] N_D[7]_c_3035_n N_D[7]_c_3036_n N_D[7]_c_3037_n
+ N_D[7]_c_3038_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[7]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_4239_265# N_A_4239_265#_M1032_d
+ N_A_4239_265#_M1064_s N_A_4239_265#_c_3131_n N_A_4239_265#_M1002_g
+ N_A_4239_265#_c_3132_n N_A_4239_265#_c_3133_n N_A_4239_265#_c_3134_n
+ N_A_4239_265#_M1023_g N_A_4239_265#_c_3135_n N_A_4239_265#_c_3136_n
+ N_A_4239_265#_M1099_g N_A_4239_265#_c_3137_n N_A_4239_265#_c_3138_n
+ N_A_4239_265#_M1143_g N_A_4239_265#_c_3139_n N_A_4239_265#_c_3140_n
+ N_A_4239_265#_c_3124_n N_A_4239_265#_c_3125_n N_A_4239_265#_c_3126_n
+ N_A_4239_265#_c_3127_n N_A_4239_265#_c_3143_n N_A_4239_265#_c_3128_n
+ N_A_4239_265#_c_3129_n N_A_4239_265#_c_3145_n N_A_4239_265#_c_3130_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_4239_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_4239_793# N_A_4239_793#_M1114_d
+ N_A_4239_793#_M1119_s N_A_4239_793#_c_3246_n N_A_4239_793#_M1011_g
+ N_A_4239_793#_c_3247_n N_A_4239_793#_c_3248_n N_A_4239_793#_c_3249_n
+ N_A_4239_793#_M1053_g N_A_4239_793#_c_3250_n N_A_4239_793#_c_3251_n
+ N_A_4239_793#_M1075_g N_A_4239_793#_c_3252_n N_A_4239_793#_c_3253_n
+ N_A_4239_793#_M1096_g N_A_4239_793#_c_3254_n N_A_4239_793#_c_3255_n
+ N_A_4239_793#_c_3239_n N_A_4239_793#_c_3240_n N_A_4239_793#_c_3258_n
+ N_A_4239_793#_c_3259_n N_A_4239_793#_c_3241_n N_A_4239_793#_c_3242_n
+ N_A_4239_793#_c_3260_n N_A_4239_793#_c_3243_n N_A_4239_793#_c_3244_n
+ N_A_4239_793#_c_3245_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_4239_793#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[6] N_S[6]_c_3360_n N_S[6]_M1089_g
+ N_S[6]_c_3361_n N_S[6]_c_3362_n N_S[6]_c_3363_n N_S[6]_M1101_g N_S[6]_c_3364_n
+ N_S[6]_c_3365_n N_S[6]_M1122_g N_S[6]_c_3366_n N_S[6]_c_3367_n N_S[6]_M1132_g
+ N_S[6]_c_3368_n N_S[6]_c_3369_n N_S[6]_c_3370_n N_S[6]_c_3371_n
+ N_S[6]_c_3372_n N_S[6]_c_3383_n N_S[6]_M1064_g N_S[6]_c_3373_n N_S[6]_M1032_g
+ N_S[6]_c_3374_n N_S[6]_c_3375_n N_S[6]_M1061_g N_S[6]_c_3376_n N_S[6]_M1085_g
+ N_S[6]_c_3377_n N_S[6]_c_3378_n N_S[6]_c_3379_n N_S[6]_c_3380_n S[6]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[6]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[7] N_S[7]_c_3470_n N_S[7]_M1008_g
+ N_S[7]_c_3471_n N_S[7]_c_3472_n N_S[7]_c_3473_n N_S[7]_M1063_g N_S[7]_c_3474_n
+ N_S[7]_c_3475_n N_S[7]_M1091_g N_S[7]_c_3476_n N_S[7]_c_3477_n N_S[7]_M1144_g
+ N_S[7]_c_3478_n N_S[7]_c_3479_n N_S[7]_c_3480_n N_S[7]_c_3481_n
+ N_S[7]_c_3491_n N_S[7]_c_3482_n N_S[7]_c_3493_n N_S[7]_M1119_g N_S[7]_c_3483_n
+ N_S[7]_M1114_g N_S[7]_c_3484_n N_S[7]_c_3485_n N_S[7]_M1149_g N_S[7]_c_3495_n
+ N_S[7]_M1148_g N_S[7]_c_3486_n N_S[7]_c_3487_n N_S[7]_c_3488_n N_S[7]_c_3489_n
+ S[7] PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[7]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%VPWR N_VPWR_M1001_d N_VPWR_M1052_d
+ N_VPWR_M1040_d N_VPWR_M1088_d N_VPWR_M1012_s N_VPWR_M1017_s N_VPWR_M1049_s
+ N_VPWR_M1055_s N_VPWR_M1137_s N_VPWR_M1141_s N_VPWR_M1090_d N_VPWR_M1076_s
+ N_VPWR_M1158_d N_VPWR_M1120_s N_VPWR_M1072_d N_VPWR_M1007_s N_VPWR_M1115_d
+ N_VPWR_M1125_s N_VPWR_M1128_d N_VPWR_M1018_d N_VPWR_M1155_d N_VPWR_M1039_d
+ N_VPWR_M1042_d N_VPWR_M1046_d N_VPWR_M1062_d N_VPWR_M1070_d N_VPWR_M1127_d
+ N_VPWR_M1134_d N_VPWR_M1108_s N_VPWR_M1117_s N_VPWR_M1145_s N_VPWR_M1153_s
+ N_VPWR_M1064_d N_VPWR_M1119_d N_VPWR_M1085_d N_VPWR_M1148_d N_VPWR_c_3586_n
+ N_VPWR_c_3587_n N_VPWR_c_3588_n N_VPWR_c_3589_n N_VPWR_c_3590_n
+ N_VPWR_c_3591_n N_VPWR_c_3592_n N_VPWR_c_3593_n N_VPWR_c_3594_n
+ N_VPWR_c_3595_n N_VPWR_c_3596_n N_VPWR_c_3597_n N_VPWR_c_3598_n
+ N_VPWR_c_3599_n N_VPWR_c_3600_n N_VPWR_c_3601_n N_VPWR_c_3602_n
+ N_VPWR_c_3603_n N_VPWR_c_3604_n N_VPWR_c_3605_n N_VPWR_c_3606_n
+ N_VPWR_c_3607_n N_VPWR_c_3608_n N_VPWR_c_3609_n N_VPWR_c_3610_n
+ N_VPWR_c_3611_n N_VPWR_c_3612_n N_VPWR_c_3613_n N_VPWR_c_3614_n
+ N_VPWR_c_3615_n N_VPWR_c_3616_n N_VPWR_c_3617_n N_VPWR_c_3618_n
+ N_VPWR_c_3619_n N_VPWR_c_3620_n N_VPWR_c_3621_n N_VPWR_c_3622_n
+ N_VPWR_c_3623_n N_VPWR_c_3624_n N_VPWR_c_3625_n N_VPWR_c_3626_n
+ N_VPWR_c_3627_n N_VPWR_c_3628_n N_VPWR_c_3629_n N_VPWR_c_3630_n
+ N_VPWR_c_3631_n N_VPWR_c_3632_n N_VPWR_c_3633_n N_VPWR_c_3634_n
+ N_VPWR_c_3635_n N_VPWR_c_3636_n N_VPWR_c_3637_n N_VPWR_c_3638_n
+ N_VPWR_c_3639_n N_VPWR_c_3640_n VPWR VPWR VPWR N_VPWR_c_3641_n N_VPWR_c_3642_n
+ N_VPWR_c_3643_n N_VPWR_c_3644_n N_VPWR_c_3645_n N_VPWR_c_3646_n
+ N_VPWR_c_3647_n N_VPWR_c_3648_n N_VPWR_c_3649_n N_VPWR_c_3650_n
+ N_VPWR_c_3651_n N_VPWR_c_3652_n N_VPWR_c_3653_n N_VPWR_c_3654_n
+ N_VPWR_c_3655_n N_VPWR_c_3656_n N_VPWR_c_3657_n N_VPWR_c_3658_n
+ N_VPWR_c_3659_n N_VPWR_c_3660_n N_VPWR_c_3661_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%VPWR
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_355_311# N_A_355_311#_M1010_d
+ N_A_355_311#_M1019_d N_A_355_311#_M1147_d N_A_355_311#_M1012_d
+ N_A_355_311#_M1086_d N_A_355_311#_c_4334_n N_A_355_311#_c_4335_n
+ N_A_355_311#_c_4356_n N_A_355_311#_c_4360_n N_A_355_311#_c_4364_n
+ N_A_355_311#_c_4343_n N_A_355_311#_c_4385_n N_A_355_311#_c_4345_n
+ N_A_355_311#_c_4388_n N_A_355_311#_c_4336_n N_A_355_311#_c_4393_n
+ N_A_355_311#_c_4369_n N_A_355_311#_c_4399_n N_A_355_311#_c_4371_n
+ N_A_355_311#_c_4406_n N_A_355_311#_c_4374_n N_A_355_311#_c_4337_n
+ N_A_355_311#_c_4338_n N_A_355_311#_c_4339_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_355_311#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_355_613# N_A_355_613#_M1054_d
+ N_A_355_613#_M1080_d N_A_355_613#_M1123_d N_A_355_613#_M1017_d
+ N_A_355_613#_M1093_d N_A_355_613#_c_4461_n N_A_355_613#_c_4462_n
+ N_A_355_613#_c_4483_n N_A_355_613#_c_4487_n N_A_355_613#_c_4491_n
+ N_A_355_613#_c_4470_n N_A_355_613#_c_4512_n N_A_355_613#_c_4472_n
+ N_A_355_613#_c_4515_n N_A_355_613#_c_4463_n N_A_355_613#_c_4520_n
+ N_A_355_613#_c_4496_n N_A_355_613#_c_4526_n N_A_355_613#_c_4529_n
+ N_A_355_613#_c_4464_n N_A_355_613#_c_4465_n N_A_355_613#_c_4466_n
+ N_A_355_613#_c_4499_n N_A_355_613#_c_4502_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_355_613#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%Z N_Z_M1003_s N_Z_M1029_s N_Z_M1109_s
+ N_Z_M1083_s N_Z_M1024_d N_Z_M1016_d N_Z_M1044_d N_Z_M1048_d N_Z_M1006_s
+ N_Z_M1009_d N_Z_M1035_s N_Z_M1112_d N_Z_M1089_s N_Z_M1008_d N_Z_M1122_s
+ N_Z_M1091_d N_Z_M1010_s N_Z_M1054_s N_Z_M1051_s N_Z_M1092_s N_Z_M1050_d
+ N_Z_M1031_d N_Z_M1116_d N_Z_M1124_d N_Z_M1004_d N_Z_M1021_s N_Z_M1131_d
+ N_Z_M1056_s N_Z_M1002_s N_Z_M1011_s N_Z_M1099_s N_Z_M1075_s N_Z_c_4588_n
+ N_Z_c_4589_n N_Z_c_4590_n N_Z_c_4591_n N_Z_c_4592_n N_Z_c_4593_n N_Z_c_4594_n
+ N_Z_c_4595_n N_Z_c_4596_n N_Z_c_4597_n N_Z_c_4598_n N_Z_c_4599_n N_Z_c_4600_n
+ N_Z_c_4601_n N_Z_c_4602_n N_Z_c_4603_n N_Z_c_4604_n N_Z_c_4605_n N_Z_c_4606_n
+ N_Z_c_4607_n N_Z_c_4608_n N_Z_c_4609_n N_Z_c_4610_n N_Z_c_4611_n N_Z_c_4612_n
+ N_Z_c_4613_n N_Z_c_4614_n N_Z_c_4615_n N_Z_c_4616_n N_Z_c_4617_n N_Z_c_4618_n
+ N_Z_c_4619_n N_Z_c_4620_n N_Z_c_4621_n N_Z_c_4622_n N_Z_c_4623_n N_Z_c_4624_n
+ N_Z_c_4625_n N_Z_c_4626_n N_Z_c_4627_n N_Z_c_4628_n N_Z_c_4629_n N_Z_c_4630_n
+ N_Z_c_4631_n N_Z_c_4632_n N_Z_c_4633_n N_Z_c_4634_n N_Z_c_4635_n N_Z_c_4644_n
+ N_Z_c_5128_n N_Z_c_4645_n N_Z_c_5164_n N_Z_c_4646_n N_Z_c_5203_p N_Z_c_4647_n
+ N_Z_c_5243_p N_Z_c_4648_n N_Z_c_5279_p N_Z_c_4649_n N_Z_c_5319_p N_Z_c_4693_n
+ N_Z_c_4718_n N_Z_c_5197_p N_Z_c_5237_p N_Z_c_4895_n N_Z_c_4924_n N_Z_c_5356_p
+ N_Z_c_5390_p Z Z Z Z Z Z Z Z N_Z_c_4650_n N_Z_c_4651_n N_Z_c_4652_n
+ N_Z_c_4653_n N_Z_c_4654_n N_Z_c_4655_n N_Z_c_4656_n N_Z_c_4657_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%Z
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1313_297# N_A_1313_297#_M1071_s
+ N_A_1313_297#_M1118_s N_A_1313_297#_M1050_s N_A_1313_297#_M1073_s
+ N_A_1313_297#_M1126_s N_A_1313_297#_c_5507_n N_A_1313_297#_c_5502_n
+ N_A_1313_297#_c_5512_n N_A_1313_297#_c_5516_n N_A_1313_297#_c_5520_n
+ N_A_1313_297#_c_5555_n N_A_1313_297#_c_5503_n N_A_1313_297#_c_5562_n
+ N_A_1313_297#_c_5531_n N_A_1313_297#_c_5566_n N_A_1313_297#_c_5533_n
+ N_A_1313_297#_c_5569_n N_A_1313_297#_c_5523_n N_A_1313_297#_c_5526_n
+ N_A_1313_297#_c_5578_n N_A_1313_297#_c_5504_n N_A_1313_297#_c_5505_n
+ N_A_1313_297#_c_5506_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1313_297#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1313_591# N_A_1313_591#_M1000_d
+ N_A_1313_591#_M1095_d N_A_1313_591#_M1031_s N_A_1313_591#_M1036_s
+ N_A_1313_591#_M1152_s N_A_1313_591#_c_5635_n N_A_1313_591#_c_5630_n
+ N_A_1313_591#_c_5640_n N_A_1313_591#_c_5644_n N_A_1313_591#_c_5648_n
+ N_A_1313_591#_c_5683_n N_A_1313_591#_c_5631_n N_A_1313_591#_c_5690_n
+ N_A_1313_591#_c_5659_n N_A_1313_591#_c_5694_n N_A_1313_591#_c_5661_n
+ N_A_1313_591#_c_5697_n N_A_1313_591#_c_5698_n N_A_1313_591#_c_5651_n
+ N_A_1313_591#_c_5654_n N_A_1313_591#_c_5632_n N_A_1313_591#_c_5633_n
+ N_A_1313_591#_c_5634_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1313_591#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2839_311# N_A_2839_311#_M1004_s
+ N_A_2839_311#_M1110_s N_A_2839_311#_M1146_s N_A_2839_311#_M1042_s
+ N_A_2839_311#_M1105_s N_A_2839_311#_c_5758_n N_A_2839_311#_c_5759_n
+ N_A_2839_311#_c_5780_n N_A_2839_311#_c_5784_n N_A_2839_311#_c_5788_n
+ N_A_2839_311#_c_5767_n N_A_2839_311#_c_5809_n N_A_2839_311#_c_5769_n
+ N_A_2839_311#_c_5812_n N_A_2839_311#_c_5760_n N_A_2839_311#_c_5817_n
+ N_A_2839_311#_c_5793_n N_A_2839_311#_c_5823_n N_A_2839_311#_c_5795_n
+ N_A_2839_311#_c_5830_n N_A_2839_311#_c_5798_n N_A_2839_311#_c_5761_n
+ N_A_2839_311#_c_5762_n N_A_2839_311#_c_5763_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2839_311#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2839_613# N_A_2839_613#_M1021_d
+ N_A_2839_613#_M1041_d N_A_2839_613#_M1078_d N_A_2839_613#_M1046_s
+ N_A_2839_613#_M1113_s N_A_2839_613#_c_5889_n N_A_2839_613#_c_5890_n
+ N_A_2839_613#_c_5911_n N_A_2839_613#_c_5915_n N_A_2839_613#_c_5919_n
+ N_A_2839_613#_c_5898_n N_A_2839_613#_c_5940_n N_A_2839_613#_c_5900_n
+ N_A_2839_613#_c_5943_n N_A_2839_613#_c_5891_n N_A_2839_613#_c_5948_n
+ N_A_2839_613#_c_5924_n N_A_2839_613#_c_5954_n N_A_2839_613#_c_5957_n
+ N_A_2839_613#_c_5892_n N_A_2839_613#_c_5893_n N_A_2839_613#_c_5894_n
+ N_A_2839_613#_c_5927_n N_A_2839_613#_c_5930_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2839_613#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3797_297# N_A_3797_297#_M1082_d
+ N_A_3797_297#_M1130_d N_A_3797_297#_M1002_d N_A_3797_297#_M1023_d
+ N_A_3797_297#_M1143_d N_A_3797_297#_c_6025_n N_A_3797_297#_c_6020_n
+ N_A_3797_297#_c_6030_n N_A_3797_297#_c_6034_n N_A_3797_297#_c_6038_n
+ N_A_3797_297#_c_6073_n N_A_3797_297#_c_6021_n N_A_3797_297#_c_6080_n
+ N_A_3797_297#_c_6049_n N_A_3797_297#_c_6084_n N_A_3797_297#_c_6051_n
+ N_A_3797_297#_c_6087_n N_A_3797_297#_c_6041_n N_A_3797_297#_c_6044_n
+ N_A_3797_297#_c_6096_n N_A_3797_297#_c_6022_n N_A_3797_297#_c_6023_n
+ N_A_3797_297#_c_6024_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3797_297#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3797_591# N_A_3797_591#_M1087_d
+ N_A_3797_591#_M1139_d N_A_3797_591#_M1011_d N_A_3797_591#_M1053_d
+ N_A_3797_591#_M1096_d N_A_3797_591#_c_6147_n N_A_3797_591#_c_6142_n
+ N_A_3797_591#_c_6152_n N_A_3797_591#_c_6156_n N_A_3797_591#_c_6160_n
+ N_A_3797_591#_c_6195_n N_A_3797_591#_c_6143_n N_A_3797_591#_c_6202_n
+ N_A_3797_591#_c_6171_n N_A_3797_591#_c_6206_n N_A_3797_591#_c_6173_n
+ N_A_3797_591#_c_6209_n N_A_3797_591#_c_6210_n N_A_3797_591#_c_6163_n
+ N_A_3797_591#_c_6166_n N_A_3797_591#_c_6144_n N_A_3797_591#_c_6145_n
+ N_A_3797_591#_c_6146_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3797_591#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%VGND N_VGND_M1043_d N_VGND_M1084_s
+ N_VGND_M1067_d N_VGND_M1138_s N_VGND_M1065_s N_VGND_M1030_s N_VGND_M1097_s
+ N_VGND_M1059_s N_VGND_M1156_s N_VGND_M1157_s N_VGND_M1037_d N_VGND_M1047_s
+ N_VGND_M1150_d N_VGND_M1136_s N_VGND_M1094_d N_VGND_M1060_d N_VGND_M1103_d
+ N_VGND_M1140_d N_VGND_M1121_d N_VGND_M1074_d N_VGND_M1129_d N_VGND_M1154_d
+ N_VGND_M1027_d N_VGND_M1033_d N_VGND_M1034_d N_VGND_M1077_d N_VGND_M1079_d
+ N_VGND_M1107_d N_VGND_M1081_s N_VGND_M1025_d N_VGND_M1159_s N_VGND_M1098_d
+ N_VGND_M1032_s N_VGND_M1114_s N_VGND_M1061_s N_VGND_M1149_s N_VGND_c_6264_n
+ N_VGND_c_6265_n N_VGND_c_6266_n N_VGND_c_6267_n N_VGND_c_6268_n
+ N_VGND_c_6269_n N_VGND_c_6270_n N_VGND_c_6271_n N_VGND_c_6272_n
+ N_VGND_c_6273_n N_VGND_c_6274_n N_VGND_c_6275_n N_VGND_c_6276_n
+ N_VGND_c_6277_n N_VGND_c_6278_n N_VGND_c_6279_n N_VGND_c_6280_n
+ N_VGND_c_6281_n N_VGND_c_6282_n N_VGND_c_6283_n N_VGND_c_6284_n
+ N_VGND_c_6285_n N_VGND_c_6286_n N_VGND_c_6287_n N_VGND_c_6288_n
+ N_VGND_c_6289_n N_VGND_c_6290_n N_VGND_c_6291_n N_VGND_c_6292_n
+ N_VGND_c_6293_n N_VGND_c_6294_n N_VGND_c_6295_n N_VGND_c_6296_n
+ N_VGND_c_6297_n N_VGND_c_6298_n N_VGND_c_6299_n N_VGND_c_6300_n
+ N_VGND_c_6301_n N_VGND_c_6302_n N_VGND_c_6303_n N_VGND_c_6304_n
+ N_VGND_c_6305_n N_VGND_c_6306_n N_VGND_c_6307_n N_VGND_c_6308_n
+ N_VGND_c_6309_n N_VGND_c_6310_n N_VGND_c_6311_n N_VGND_c_6312_n
+ N_VGND_c_6313_n N_VGND_c_6314_n N_VGND_c_6315_n N_VGND_c_6316_n
+ N_VGND_c_6317_n N_VGND_c_6318_n N_VGND_c_6319_n N_VGND_c_6320_n
+ N_VGND_c_6321_n N_VGND_c_6322_n N_VGND_c_6323_n N_VGND_c_6324_n
+ N_VGND_c_6325_n N_VGND_c_6326_n N_VGND_c_6327_n N_VGND_c_6328_n
+ N_VGND_c_6329_n N_VGND_c_6330_n N_VGND_c_6331_n N_VGND_c_6332_n
+ N_VGND_c_6333_n N_VGND_c_6334_n N_VGND_c_6335_n N_VGND_c_6336_n
+ N_VGND_c_6337_n N_VGND_c_6338_n N_VGND_c_6339_n VGND VGND VGND VGND VGND VGND
+ N_VGND_c_6340_n N_VGND_c_6341_n N_VGND_c_6342_n N_VGND_c_6343_n
+ N_VGND_c_6344_n N_VGND_c_6345_n N_VGND_c_6346_n N_VGND_c_6347_n
+ N_VGND_c_6348_n N_VGND_c_6349_n N_VGND_c_6350_n N_VGND_c_6351_n
+ N_VGND_c_6352_n N_VGND_c_6353_n N_VGND_c_6354_n N_VGND_c_6355_n
+ N_VGND_c_6356_n N_VGND_c_6357_n N_VGND_c_6358_n N_VGND_c_6359_n
+ N_VGND_c_6360_n N_VGND_c_6361_n N_VGND_c_6362_n N_VGND_c_6363_n
+ N_VGND_c_6364_n N_VGND_c_6365_n N_VGND_c_6366_n N_VGND_c_6367_n
+ N_VGND_c_6368_n N_VGND_c_6369_n N_VGND_c_6370_n N_VGND_c_6371_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%VGND
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_405_66# N_A_405_66#_M1003_d
+ N_A_405_66#_M1100_d N_A_405_66#_M1133_d N_A_405_66#_M1065_d
+ N_A_405_66#_M1151_d N_A_405_66#_c_6926_n N_A_405_66#_c_6927_n
+ N_A_405_66#_c_6928_n N_A_405_66#_c_6948_n N_A_405_66#_c_6929_n
+ N_A_405_66#_c_6930_n N_A_405_66#_c_6931_n N_A_405_66#_c_6932_n
+ N_A_405_66#_c_6951_n N_A_405_66#_c_6933_n N_A_405_66#_c_6960_n
+ N_A_405_66#_c_6945_n N_A_405_66#_c_6934_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_405_66#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_405_918# N_A_405_918#_M1029_d
+ N_A_405_918#_M1058_d N_A_405_918#_M1102_d N_A_405_918#_M1030_d
+ N_A_405_918#_M1068_d N_A_405_918#_c_7010_n N_A_405_918#_c_7011_n
+ N_A_405_918#_c_7012_n N_A_405_918#_c_7032_n N_A_405_918#_c_7013_n
+ N_A_405_918#_c_7014_n N_A_405_918#_c_7015_n N_A_405_918#_c_7016_n
+ N_A_405_918#_c_7035_n N_A_405_918#_c_7029_n N_A_405_918#_c_7017_n
+ N_A_405_918#_c_7018_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_405_918#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1315_47# N_A_1315_47#_M1013_s
+ N_A_1315_47#_M1069_s N_A_1315_47#_M1024_s N_A_1315_47#_M1028_s
+ N_A_1315_47#_M1057_s N_A_1315_47#_c_7100_n N_A_1315_47#_c_7103_n
+ N_A_1315_47#_c_7092_n N_A_1315_47#_c_7111_n N_A_1315_47#_c_7093_n
+ N_A_1315_47#_c_7094_n N_A_1315_47#_c_7095_n N_A_1315_47#_c_7096_n
+ N_A_1315_47#_c_7120_n N_A_1315_47#_c_7097_n N_A_1315_47#_c_7098_n
+ N_A_1315_47#_c_7099_n N_A_1315_47#_c_7133_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1315_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1315_911# N_A_1315_911#_M1015_d
+ N_A_1315_911#_M1104_d N_A_1315_911#_M1016_s N_A_1315_911#_M1020_s
+ N_A_1315_911#_M1135_s N_A_1315_911#_c_7183_n N_A_1315_911#_c_7175_n
+ N_A_1315_911#_c_7176_n N_A_1315_911#_c_7177_n N_A_1315_911#_c_7178_n
+ N_A_1315_911#_c_7199_n N_A_1315_911#_c_7179_n N_A_1315_911#_c_7180_n
+ N_A_1315_911#_c_7181_n N_A_1315_911#_c_7182_n N_A_1315_911#_c_7212_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1315_911#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2889_66# N_A_2889_66#_M1006_d
+ N_A_2889_66#_M1022_d N_A_2889_66#_M1066_d N_A_2889_66#_M1027_s
+ N_A_2889_66#_M1045_s N_A_2889_66#_c_7254_n N_A_2889_66#_c_7255_n
+ N_A_2889_66#_c_7256_n N_A_2889_66#_c_7276_n N_A_2889_66#_c_7257_n
+ N_A_2889_66#_c_7258_n N_A_2889_66#_c_7259_n N_A_2889_66#_c_7260_n
+ N_A_2889_66#_c_7279_n N_A_2889_66#_c_7261_n N_A_2889_66#_c_7288_n
+ N_A_2889_66#_c_7273_n N_A_2889_66#_c_7262_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2889_66#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2889_918# N_A_2889_918#_M1009_s
+ N_A_2889_918#_M1038_s N_A_2889_918#_M1142_s N_A_2889_918#_M1033_s
+ N_A_2889_918#_M1106_s N_A_2889_918#_c_7338_n N_A_2889_918#_c_7339_n
+ N_A_2889_918#_c_7340_n N_A_2889_918#_c_7360_n N_A_2889_918#_c_7341_n
+ N_A_2889_918#_c_7342_n N_A_2889_918#_c_7343_n N_A_2889_918#_c_7344_n
+ N_A_2889_918#_c_7363_n N_A_2889_918#_c_7357_n N_A_2889_918#_c_7345_n
+ N_A_2889_918#_c_7346_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2889_918#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3799_47# N_A_3799_47#_M1005_d
+ N_A_3799_47#_M1111_d N_A_3799_47#_M1089_d N_A_3799_47#_M1101_d
+ N_A_3799_47#_M1132_d N_A_3799_47#_c_7428_n N_A_3799_47#_c_7431_n
+ N_A_3799_47#_c_7420_n N_A_3799_47#_c_7439_n N_A_3799_47#_c_7421_n
+ N_A_3799_47#_c_7422_n N_A_3799_47#_c_7423_n N_A_3799_47#_c_7424_n
+ N_A_3799_47#_c_7448_n N_A_3799_47#_c_7425_n N_A_3799_47#_c_7426_n
+ N_A_3799_47#_c_7427_n N_A_3799_47#_c_7461_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3799_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3799_911# N_A_3799_911#_M1014_s
+ N_A_3799_911#_M1026_s N_A_3799_911#_M1008_s N_A_3799_911#_M1063_s
+ N_A_3799_911#_M1144_s N_A_3799_911#_c_7511_n N_A_3799_911#_c_7503_n
+ N_A_3799_911#_c_7504_n N_A_3799_911#_c_7505_n N_A_3799_911#_c_7506_n
+ N_A_3799_911#_c_7527_n N_A_3799_911#_c_7507_n N_A_3799_911#_c_7508_n
+ N_A_3799_911#_c_7509_n N_A_3799_911#_c_7510_n N_A_3799_911#_c_7540_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3799_911#
cc_1 VNB N_S[0]_c_904_n 0.0378855f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_2 VNB N_S[0]_c_905_n 0.0330319f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_3 VNB N_S[0]_c_906_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.735
cc_4 VNB N_S[0]_c_907_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.81
cc_5 VNB N_S[0]_c_908_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_6 VNB N_S[0]_c_909_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_7 VNB N_S[0]_c_910_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_8 VNB N_S[0]_c_911_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_9 VNB N_S[0]_c_912_n 0.046608f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_10 VNB N_S[0]_c_913_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=0.18
cc_11 VNB N_S[0]_c_914_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.255
cc_12 VNB N_S[0]_c_915_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.18
cc_13 VNB N_S[0]_c_916_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.255
cc_14 VNB N_S[0]_c_917_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_15 VNB N_S[0]_c_918_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_16 VNB N_S[0]_c_919_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=3.545 $Y2=0.18
cc_17 VNB N_S[0]_c_920_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.255
cc_18 VNB N_S[0]_c_921_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_19 VNB N_S[0]_c_922_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_20 VNB N_S[0]_c_923_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_21 VNB N_S[0]_c_924_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.18
cc_22 VNB N_S[0]_c_925_n 0.0131272f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_23 VNB N_S[1]_c_1016_n 0.0378855f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_24 VNB N_S[1]_c_1017_n 0.0525882f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.735
cc_25 VNB N_S[1]_c_1018_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.81
cc_26 VNB N_S[1]_c_1019_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.445
cc_27 VNB N_S[1]_c_1020_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.445
cc_28 VNB N_S[1]_c_1021_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_29 VNB N_S[1]_c_1022_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_30 VNB N_S[1]_c_1023_n 0.046608f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_31 VNB N_S[1]_c_1024_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=0.18
cc_32 VNB N_S[1]_c_1025_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.255
cc_33 VNB N_S[1]_c_1026_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.18
cc_34 VNB N_S[1]_c_1027_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.255
cc_35 VNB N_S[1]_c_1028_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_36 VNB N_S[1]_c_1029_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_37 VNB N_S[1]_c_1030_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=3.545 $Y2=0.18
cc_38 VNB N_S[1]_c_1031_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.255
cc_39 VNB N_S[1]_c_1032_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_40 VNB N_S[1]_c_1033_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_41 VNB N_S[1]_c_1034_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_42 VNB N_S[1]_c_1035_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.18
cc_43 VNB N_S[1]_c_1036_n 0.0131272f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_44 VNB N_A_142_325#_c_1134_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_45 VNB N_A_142_325#_c_1135_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_46 VNB N_A_142_325#_c_1136_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_47 VNB N_A_142_325#_c_1137_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_48 VNB N_A_142_325#_c_1138_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_142_325#_c_1139_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=0.81
cc_50 VNB N_A_142_325#_c_1140_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_51 VNB N_A_142_599#_c_1246_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_52 VNB N_A_142_599#_c_1247_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_53 VNB N_A_142_599#_c_1248_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_54 VNB N_A_142_599#_c_1249_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_55 VNB N_A_142_599#_c_1250_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_142_599#_c_1251_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=0.81
cc_57 VNB N_A_142_599#_c_1252_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_58 VNB N_D[0]_M1012_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_59 VNB N_D[0]_M1065_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.445
cc_60 VNB N_D[0]_M1097_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_61 VNB N_D[0]_M1049_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_62 VNB N_D[0]_M1086_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_63 VNB N_D[0]_M1151_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_64 VNB N_D[0]_M1156_g 0.0199741f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_65 VNB N_D[0]_M1137_g 4.3907e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_66 VNB N_D[0]_c_1372_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_67 VNB N_D[0]_c_1373_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_68 VNB N_D[0]_c_1374_n 0.00220429f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_69 VNB N_D[0]_c_1375_n 0.0314703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_D[1]_M1017_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_71 VNB N_D[1]_M1030_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.445
cc_72 VNB N_D[1]_M1059_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_73 VNB N_D[1]_M1055_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_74 VNB N_D[1]_M1093_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_75 VNB N_D[1]_M1068_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_76 VNB N_D[1]_M1157_g 0.0199741f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_77 VNB N_D[1]_M1141_g 4.3907e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_78 VNB N_D[1]_c_1471_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_79 VNB N_D[1]_c_1472_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_80 VNB N_D[1]_c_1473_n 0.00220429f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_81 VNB N_D[1]_c_1474_n 0.0314703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_D[2]_M1071_g 4.3907e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_83 VNB N_D[2]_M1013_g 0.0199741f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.445
cc_84 VNB N_D[2]_M1037_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_85 VNB N_D[2]_M1090_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_86 VNB N_D[2]_M1118_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_87 VNB N_D[2]_M1069_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_88 VNB N_D[2]_M1150_g 0.024303f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_89 VNB N_D[2]_M1158_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_90 VNB N_D[2]_c_1568_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_91 VNB N_D[2]_c_1569_n 0.0314703f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_92 VNB N_D[2]_c_1570_n 0.00220429f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_93 VNB N_D[2]_c_1571_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_94 VNB N_D[3]_M1000_g 4.3907e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_95 VNB N_D[3]_M1015_g 0.0199741f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.445
cc_96 VNB N_D[3]_M1047_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_97 VNB N_D[3]_M1076_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_98 VNB N_D[3]_M1095_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_99 VNB N_D[3]_M1104_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_100 VNB N_D[3]_M1136_g 0.024303f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_101 VNB N_D[3]_M1120_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_102 VNB N_D[3]_c_1669_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_103 VNB N_D[3]_c_1670_n 0.0314703f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_104 VNB N_D[3]_c_1671_n 0.00220429f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_105 VNB N_D[3]_c_1672_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_106 VNB N_A_1755_265#_c_1758_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_107 VNB N_A_1755_265#_c_1759_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=2.855
+ $Y2=0.18
cc_108 VNB N_A_1755_265#_c_1760_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_109 VNB N_A_1755_265#_c_1761_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=3.62
+ $Y2=0.255
cc_110 VNB N_A_1755_265#_c_1762_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_111 VNB N_A_1755_265#_c_1763_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_A_1755_265#_c_1764_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_113 VNB N_A_1755_793#_c_1877_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_114 VNB N_A_1755_793#_c_1878_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=2.855
+ $Y2=0.18
cc_115 VNB N_A_1755_793#_c_1879_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_116 VNB N_A_1755_793#_c_1880_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_117 VNB N_A_1755_793#_c_1881_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_A_1755_793#_c_1882_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0.62
+ $Y2=0.81
cc_119 VNB N_A_1755_793#_c_1883_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_120 VNB N_S[2]_c_2002_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_121 VNB N_S[2]_c_2003_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=2.035
cc_122 VNB N_S[2]_c_2004_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=2.035
cc_123 VNB N_S[2]_c_2005_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.735
cc_124 VNB N_S[2]_c_2006_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.81
cc_125 VNB N_S[2]_c_2007_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_126 VNB N_S[2]_c_2008_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.885
cc_127 VNB N_S[2]_c_2009_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.55
cc_128 VNB N_S[2]_c_2010_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_129 VNB N_S[2]_c_2011_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_130 VNB N_S[2]_c_2012_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_131 VNB N_S[2]_c_2013_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=0.18
cc_132 VNB N_S[2]_c_2014_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_133 VNB N_S[2]_c_2015_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.255
cc_134 VNB N_S[2]_c_2016_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_135 VNB N_S[2]_c_2017_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_136 VNB N_S[2]_c_2018_n 0.065295f $X=-0.19 $Y=-0.24 $X2=3.545 $Y2=0.18
cc_137 VNB N_S[2]_c_2019_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_138 VNB N_S[2]_c_2020_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_139 VNB N_S[2]_c_2021_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_140 VNB N_S[2]_c_2022_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_141 VNB S[2] 0.00265247f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_142 VNB N_S[3]_c_2119_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_143 VNB N_S[3]_c_2120_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=2.035
cc_144 VNB N_S[3]_c_2121_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=2.035
cc_145 VNB N_S[3]_c_2122_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.735
cc_146 VNB N_S[3]_c_2123_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.81
cc_147 VNB N_S[3]_c_2124_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_148 VNB N_S[3]_c_2125_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.885
cc_149 VNB N_S[3]_c_2126_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.55
cc_150 VNB N_S[3]_c_2127_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_151 VNB N_S[3]_c_2128_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_152 VNB N_S[3]_c_2129_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_153 VNB N_S[3]_c_2130_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=0.18
cc_154 VNB N_S[3]_c_2131_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_155 VNB N_S[3]_c_2132_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.255
cc_156 VNB N_S[3]_c_2133_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_157 VNB N_S[3]_c_2134_n 0.0848512f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_158 VNB N_S[3]_c_2135_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_159 VNB N_S[3]_c_2136_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_160 VNB N_S[3]_c_2137_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_161 VNB N_S[3]_c_2138_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_162 VNB S[3] 0.00265247f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_163 VNB N_S[4]_c_2244_n 0.032202f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_164 VNB N_S[4]_c_2245_n 0.0330319f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_165 VNB N_S[4]_c_2246_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.735
cc_166 VNB N_S[4]_c_2247_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.81
cc_167 VNB N_S[4]_c_2248_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_168 VNB N_S[4]_c_2249_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_169 VNB N_S[4]_c_2250_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_170 VNB N_S[4]_c_2251_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_171 VNB N_S[4]_c_2252_n 0.046608f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_172 VNB N_S[4]_c_2253_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=0.18
cc_173 VNB N_S[4]_c_2254_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.255
cc_174 VNB N_S[4]_c_2255_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.18
cc_175 VNB N_S[4]_c_2256_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.255
cc_176 VNB N_S[4]_c_2257_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_177 VNB N_S[4]_c_2258_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_178 VNB N_S[4]_c_2259_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=3.545 $Y2=0.18
cc_179 VNB N_S[4]_c_2260_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.255
cc_180 VNB N_S[4]_c_2261_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_181 VNB N_S[4]_c_2262_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_182 VNB N_S[4]_c_2263_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_183 VNB N_S[4]_c_2264_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.18
cc_184 VNB N_S[4]_c_2265_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_185 VNB N_S[5]_c_2364_n 0.032202f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_186 VNB N_S[5]_c_2365_n 0.0525882f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.735
cc_187 VNB N_S[5]_c_2366_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.81
cc_188 VNB N_S[5]_c_2367_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.445
cc_189 VNB N_S[5]_c_2368_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.445
cc_190 VNB N_S[5]_c_2369_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_191 VNB N_S[5]_c_2370_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_192 VNB N_S[5]_c_2371_n 0.046608f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_193 VNB N_S[5]_c_2372_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=0.18
cc_194 VNB N_S[5]_c_2373_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.255
cc_195 VNB N_S[5]_c_2374_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.18
cc_196 VNB N_S[5]_c_2375_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.255
cc_197 VNB N_S[5]_c_2376_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_198 VNB N_S[5]_c_2377_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_199 VNB N_S[5]_c_2378_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=3.545 $Y2=0.18
cc_200 VNB N_S[5]_c_2379_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.255
cc_201 VNB N_S[5]_c_2380_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_202 VNB N_S[5]_c_2381_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_203 VNB N_S[5]_c_2382_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_204 VNB N_S[5]_c_2383_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.18
cc_205 VNB N_S[5]_c_2384_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_206 VNB N_A_2626_325#_c_2492_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=1.065
+ $Y2=0.735
cc_207 VNB N_A_2626_325#_c_2493_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=3.125
+ $Y2=0.18
cc_208 VNB N_A_2626_325#_c_2494_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_209 VNB N_A_2626_325#_c_2495_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_210 VNB N_A_2626_325#_c_2496_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_211 VNB N_A_2626_325#_c_2497_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0.62
+ $Y2=0.81
cc_212 VNB N_A_2626_325#_c_2498_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_213 VNB N_A_2626_599#_c_2608_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=1.065
+ $Y2=0.735
cc_214 VNB N_A_2626_599#_c_2609_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_215 VNB N_A_2626_599#_c_2610_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=3.125
+ $Y2=0.18
cc_216 VNB N_A_2626_599#_c_2611_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_217 VNB N_A_2626_599#_c_2612_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_218 VNB N_A_2626_599#_c_2613_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0.62
+ $Y2=0.81
cc_219 VNB N_A_2626_599#_c_2614_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_220 VNB N_D[4]_M1042_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_221 VNB N_D[4]_M1027_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.445
cc_222 VNB N_D[4]_M1034_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_223 VNB N_D[4]_M1062_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_224 VNB N_D[4]_M1105_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_225 VNB N_D[4]_M1045_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_226 VNB N_D[4]_M1079_g 0.0199741f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_227 VNB N_D[4]_M1127_g 4.3907e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_228 VNB N_D[4]_c_2738_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_229 VNB N_D[4]_c_2739_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_230 VNB N_D[4]_c_2740_n 0.00220429f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_231 VNB N_D[4]_c_2741_n 0.0314703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_232 VNB N_D[5]_M1046_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_233 VNB N_D[5]_M1033_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.445
cc_234 VNB N_D[5]_M1077_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_235 VNB N_D[5]_M1070_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_236 VNB N_D[5]_M1113_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_237 VNB N_D[5]_M1106_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_238 VNB N_D[5]_M1107_g 0.0199741f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_239 VNB N_D[5]_M1134_g 4.3907e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_240 VNB N_D[5]_c_2837_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_241 VNB N_D[5]_c_2838_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_242 VNB N_D[5]_c_2839_n 0.00220429f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_243 VNB N_D[5]_c_2840_n 0.0314703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_244 VNB N_D[6]_M1082_g 4.3907e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_245 VNB N_D[6]_M1005_g 0.0199741f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.445
cc_246 VNB N_D[6]_M1081_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_247 VNB N_D[6]_M1108_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_248 VNB N_D[6]_M1130_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_249 VNB N_D[6]_M1111_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_250 VNB N_D[6]_M1159_g 0.024303f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_251 VNB N_D[6]_M1145_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_252 VNB N_D[6]_c_2934_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_253 VNB N_D[6]_c_2935_n 0.0314703f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_254 VNB N_D[6]_c_2936_n 0.00220429f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_255 VNB N_D[6]_c_2937_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_256 VNB N_D[7]_M1087_g 4.3907e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.55
cc_257 VNB N_D[7]_M1014_g 0.0199741f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.445
cc_258 VNB N_D[7]_M1025_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_259 VNB N_D[7]_M1117_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.45
cc_260 VNB N_D[7]_M1139_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_261 VNB N_D[7]_M1026_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_262 VNB N_D[7]_M1098_g 0.024303f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_263 VNB N_D[7]_M1153_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_264 VNB N_D[7]_c_3035_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_265 VNB N_D[7]_c_3036_n 0.0314703f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_266 VNB N_D[7]_c_3037_n 0.00220429f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_267 VNB N_D[7]_c_3038_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_268 VNB N_A_4239_265#_c_3124_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_269 VNB N_A_4239_265#_c_3125_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=2.855
+ $Y2=0.18
cc_270 VNB N_A_4239_265#_c_3126_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.59
cc_271 VNB N_A_4239_265#_c_3127_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=3.62
+ $Y2=0.255
cc_272 VNB N_A_4239_265#_c_3128_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_273 VNB N_A_4239_265#_c_3129_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_274 VNB N_A_4239_265#_c_3130_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_275 VNB N_A_4239_793#_c_3239_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_276 VNB N_A_4239_793#_c_3240_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=2.855
+ $Y2=0.18
cc_277 VNB N_A_4239_793#_c_3241_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_278 VNB N_A_4239_793#_c_3242_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_279 VNB N_A_4239_793#_c_3243_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_280 VNB N_A_4239_793#_c_3244_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0.62
+ $Y2=0.81
cc_281 VNB N_A_4239_793#_c_3245_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_282 VNB N_S[6]_c_3360_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_283 VNB N_S[6]_c_3361_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=2.035
cc_284 VNB N_S[6]_c_3362_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=2.035
cc_285 VNB N_S[6]_c_3363_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.735
cc_286 VNB N_S[6]_c_3364_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.81
cc_287 VNB N_S[6]_c_3365_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_288 VNB N_S[6]_c_3366_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.885
cc_289 VNB N_S[6]_c_3367_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.55
cc_290 VNB N_S[6]_c_3368_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_291 VNB N_S[6]_c_3369_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_292 VNB N_S[6]_c_3370_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_293 VNB N_S[6]_c_3371_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=0.18
cc_294 VNB N_S[6]_c_3372_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_295 VNB N_S[6]_c_3373_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.255
cc_296 VNB N_S[6]_c_3374_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_297 VNB N_S[6]_c_3375_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_298 VNB N_S[6]_c_3376_n 0.0709784f $X=-0.19 $Y=-0.24 $X2=3.545 $Y2=0.18
cc_299 VNB N_S[6]_c_3377_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_300 VNB N_S[6]_c_3378_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_301 VNB N_S[6]_c_3379_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_302 VNB N_S[6]_c_3380_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_303 VNB S[6] 0.0131272f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_304 VNB N_S[7]_c_3470_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_305 VNB N_S[7]_c_3471_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=2.035
cc_306 VNB N_S[7]_c_3472_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=2.035
cc_307 VNB N_S[7]_c_3473_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.735
cc_308 VNB N_S[7]_c_3474_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.81
cc_309 VNB N_S[7]_c_3475_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.735
cc_310 VNB N_S[7]_c_3476_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.885
cc_311 VNB N_S[7]_c_3477_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.55
cc_312 VNB N_S[7]_c_3478_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.81
cc_313 VNB N_S[7]_c_3479_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_314 VNB N_S[7]_c_3480_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.18
cc_315 VNB N_S[7]_c_3481_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=0.18
cc_316 VNB N_S[7]_c_3482_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_317 VNB N_S[7]_c_3483_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.255
cc_318 VNB N_S[7]_c_3484_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_319 VNB N_S[7]_c_3485_n 0.0905347f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=0.255
cc_320 VNB N_S[7]_c_3486_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_321 VNB N_S[7]_c_3487_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_322 VNB N_S[7]_c_3488_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=0.81
cc_323 VNB N_S[7]_c_3489_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_324 VNB S[7] 0.0131272f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_325 VNB N_Z_c_4588_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_326 VNB N_Z_c_4589_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_327 VNB N_Z_c_4590_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_328 VNB N_Z_c_4591_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_329 VNB N_Z_c_4592_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_330 VNB N_Z_c_4593_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_331 VNB N_Z_c_4594_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_332 VNB N_Z_c_4595_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_333 VNB N_Z_c_4596_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_334 VNB N_Z_c_4597_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_335 VNB N_Z_c_4598_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_336 VNB N_Z_c_4599_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_337 VNB N_Z_c_4600_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_338 VNB N_Z_c_4601_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_339 VNB N_Z_c_4602_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_340 VNB N_Z_c_4603_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_341 VNB N_Z_c_4604_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_342 VNB N_Z_c_4605_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_343 VNB N_Z_c_4606_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_344 VNB N_Z_c_4607_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_345 VNB N_Z_c_4608_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_346 VNB N_Z_c_4609_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_347 VNB N_Z_c_4610_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_348 VNB N_Z_c_4611_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_349 VNB N_Z_c_4612_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_350 VNB N_Z_c_4613_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_351 VNB N_Z_c_4614_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_352 VNB N_Z_c_4615_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_353 VNB N_Z_c_4616_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_354 VNB N_Z_c_4617_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_355 VNB N_Z_c_4618_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_356 VNB N_Z_c_4619_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_357 VNB N_Z_c_4620_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_358 VNB N_Z_c_4621_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_359 VNB N_Z_c_4622_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_360 VNB N_Z_c_4623_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_361 VNB N_Z_c_4624_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_362 VNB N_Z_c_4625_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_363 VNB N_Z_c_4626_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_364 VNB N_Z_c_4627_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_365 VNB N_Z_c_4628_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_366 VNB N_Z_c_4629_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_367 VNB N_Z_c_4630_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_368 VNB N_Z_c_4631_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_369 VNB N_Z_c_4632_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_370 VNB N_Z_c_4633_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_371 VNB N_Z_c_4634_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_372 VNB N_Z_c_4635_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_373 VNB N_VGND_c_6264_n 0.0163664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_374 VNB N_VGND_c_6265_n 0.0193722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_375 VNB N_VGND_c_6266_n 0.0163664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_376 VNB N_VGND_c_6267_n 0.0193722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_377 VNB N_VGND_c_6268_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_378 VNB N_VGND_c_6269_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_379 VNB N_VGND_c_6270_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_380 VNB N_VGND_c_6271_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_381 VNB N_VGND_c_6272_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_382 VNB N_VGND_c_6273_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_383 VNB N_VGND_c_6274_n 0.00968695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_384 VNB N_VGND_c_6275_n 0.00968695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_385 VNB N_VGND_c_6276_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_386 VNB N_VGND_c_6277_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_387 VNB N_VGND_c_6278_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_388 VNB N_VGND_c_6279_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_389 VNB N_VGND_c_6280_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_390 VNB N_VGND_c_6281_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_391 VNB N_VGND_c_6282_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_392 VNB N_VGND_c_6283_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_393 VNB N_VGND_c_6284_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_394 VNB N_VGND_c_6285_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_395 VNB N_VGND_c_6286_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_396 VNB N_VGND_c_6287_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_397 VNB N_VGND_c_6288_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_398 VNB N_VGND_c_6289_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_399 VNB N_VGND_c_6290_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_400 VNB N_VGND_c_6291_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_401 VNB N_VGND_c_6292_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_402 VNB N_VGND_c_6293_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_403 VNB N_VGND_c_6294_n 0.00968695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_404 VNB N_VGND_c_6295_n 0.00968695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_405 VNB N_VGND_c_6296_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_406 VNB N_VGND_c_6297_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_407 VNB N_VGND_c_6298_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_408 VNB N_VGND_c_6299_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_409 VNB N_VGND_c_6300_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_410 VNB N_VGND_c_6301_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_411 VNB N_VGND_c_6302_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_412 VNB N_VGND_c_6303_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_413 VNB N_VGND_c_6304_n 0.0163664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_414 VNB N_VGND_c_6305_n 0.0193722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_415 VNB N_VGND_c_6306_n 0.0163664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_416 VNB N_VGND_c_6307_n 0.0193722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_417 VNB N_VGND_c_6308_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_418 VNB N_VGND_c_6309_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_419 VNB N_VGND_c_6310_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_420 VNB N_VGND_c_6311_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_421 VNB N_VGND_c_6312_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_422 VNB N_VGND_c_6313_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_423 VNB N_VGND_c_6314_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_424 VNB N_VGND_c_6315_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_425 VNB N_VGND_c_6316_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_426 VNB N_VGND_c_6317_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_427 VNB N_VGND_c_6318_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_428 VNB N_VGND_c_6319_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_429 VNB N_VGND_c_6320_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_430 VNB N_VGND_c_6321_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_431 VNB N_VGND_c_6322_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_432 VNB N_VGND_c_6323_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_433 VNB N_VGND_c_6324_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_434 VNB N_VGND_c_6325_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_435 VNB N_VGND_c_6326_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_436 VNB N_VGND_c_6327_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_437 VNB N_VGND_c_6328_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_438 VNB N_VGND_c_6329_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_439 VNB N_VGND_c_6330_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_440 VNB N_VGND_c_6331_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_441 VNB N_VGND_c_6332_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_442 VNB N_VGND_c_6333_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_443 VNB N_VGND_c_6334_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_444 VNB N_VGND_c_6335_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_445 VNB N_VGND_c_6336_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_446 VNB N_VGND_c_6337_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_447 VNB N_VGND_c_6338_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_448 VNB N_VGND_c_6339_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_449 VNB N_VGND_c_6340_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_450 VNB N_VGND_c_6341_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_451 VNB N_VGND_c_6342_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_452 VNB N_VGND_c_6343_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_453 VNB N_VGND_c_6344_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_454 VNB N_VGND_c_6345_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_455 VNB N_VGND_c_6346_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_456 VNB N_VGND_c_6347_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_457 VNB N_VGND_c_6348_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_458 VNB N_VGND_c_6349_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_459 VNB N_VGND_c_6350_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_460 VNB N_VGND_c_6351_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_461 VNB N_VGND_c_6352_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_462 VNB N_VGND_c_6353_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_463 VNB N_VGND_c_6354_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_464 VNB N_VGND_c_6355_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_465 VNB N_VGND_c_6356_n 0.00634081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_466 VNB N_VGND_c_6357_n 0.00631492f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_467 VNB N_VGND_c_6358_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_468 VNB N_VGND_c_6359_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_469 VNB N_VGND_c_6360_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_470 VNB N_VGND_c_6361_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_471 VNB N_VGND_c_6362_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_472 VNB N_VGND_c_6363_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_473 VNB N_VGND_c_6364_n 0.00634081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_474 VNB N_VGND_c_6365_n 0.00631492f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_475 VNB N_VGND_c_6366_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_476 VNB N_VGND_c_6367_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_477 VNB N_VGND_c_6368_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_478 VNB N_VGND_c_6369_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_479 VNB N_VGND_c_6370_n 1.13682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_480 VNB N_VGND_c_6371_n 1.13682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_481 VNB N_A_405_66#_c_6926_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=2.035
cc_482 VNB N_A_405_66#_c_6927_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=1.19 $Y2=0.81
cc_483 VNB N_A_405_66#_c_6928_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.255
cc_484 VNB N_A_405_66#_c_6929_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_485 VNB N_A_405_66#_c_6930_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_486 VNB N_A_405_66#_c_6931_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_487 VNB N_A_405_66#_c_6932_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.18
cc_488 VNB N_A_405_66#_c_6933_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=3.545 $Y2=0.18
cc_489 VNB N_A_405_66#_c_6934_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_490 VNB N_A_405_918#_c_7010_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=2.035
cc_491 VNB N_A_405_918#_c_7011_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=1.19 $Y2=0.81
cc_492 VNB N_A_405_918#_c_7012_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.255
cc_493 VNB N_A_405_918#_c_7013_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_494 VNB N_A_405_918#_c_7014_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_495 VNB N_A_405_918#_c_7015_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_496 VNB N_A_405_918#_c_7016_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=3.125
+ $Y2=0.18
cc_497 VNB N_A_405_918#_c_7017_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_498 VNB N_A_405_918#_c_7018_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_499 VNB N_A_1315_47#_c_7092_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.255
cc_500 VNB N_A_1315_47#_c_7093_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_501 VNB N_A_1315_47#_c_7094_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_502 VNB N_A_1315_47#_c_7095_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_503 VNB N_A_1315_47#_c_7096_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=3.125
+ $Y2=0.18
cc_504 VNB N_A_1315_47#_c_7097_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=3.545
+ $Y2=0.18
cc_505 VNB N_A_1315_47#_c_7098_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_506 VNB N_A_1315_47#_c_7099_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_507 VNB N_A_1315_911#_c_7175_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_508 VNB N_A_1315_911#_c_7176_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=2.36
+ $Y2=0.59
cc_509 VNB N_A_1315_911#_c_7177_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=2.705
+ $Y2=0.18
cc_510 VNB N_A_1315_911#_c_7178_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=2.435
+ $Y2=0.18
cc_511 VNB N_A_1315_911#_c_7179_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=2.855
+ $Y2=0.18
cc_512 VNB N_A_1315_911#_c_7180_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=3.545
+ $Y2=0.18
cc_513 VNB N_A_1315_911#_c_7181_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=3.62
+ $Y2=0.59
cc_514 VNB N_A_1315_911#_c_7182_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.09
+ $Y2=0.81
cc_515 VNB N_A_2889_66#_c_7254_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=2.035
cc_516 VNB N_A_2889_66#_c_7255_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=1.19 $Y2=0.81
cc_517 VNB N_A_2889_66#_c_7256_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.255
cc_518 VNB N_A_2889_66#_c_7257_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_519 VNB N_A_2889_66#_c_7258_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_520 VNB N_A_2889_66#_c_7259_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_521 VNB N_A_2889_66#_c_7260_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=3.125
+ $Y2=0.18
cc_522 VNB N_A_2889_66#_c_7261_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=3.545
+ $Y2=0.18
cc_523 VNB N_A_2889_66#_c_7262_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.18
cc_524 VNB N_A_2889_918#_c_7338_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=1.09
+ $Y2=2.035
cc_525 VNB N_A_2889_918#_c_7339_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=1.19
+ $Y2=0.81
cc_526 VNB N_A_2889_918#_c_7340_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=1.6
+ $Y2=0.255
cc_527 VNB N_A_2889_918#_c_7341_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_528 VNB N_A_2889_918#_c_7342_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=2.78
+ $Y2=0.59
cc_529 VNB N_A_2889_918#_c_7343_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=2.78
+ $Y2=0.59
cc_530 VNB N_A_2889_918#_c_7344_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=3.125
+ $Y2=0.18
cc_531 VNB N_A_2889_918#_c_7345_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=3.62
+ $Y2=0.59
cc_532 VNB N_A_2889_918#_c_7346_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=2.36
+ $Y2=0.18
cc_533 VNB N_A_3799_47#_c_7420_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.255
cc_534 VNB N_A_3799_47#_c_7421_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.59
cc_535 VNB N_A_3799_47#_c_7422_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_536 VNB N_A_3799_47#_c_7423_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.59
cc_537 VNB N_A_3799_47#_c_7424_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=3.125
+ $Y2=0.18
cc_538 VNB N_A_3799_47#_c_7425_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=3.545
+ $Y2=0.18
cc_539 VNB N_A_3799_47#_c_7426_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.59
cc_540 VNB N_A_3799_47#_c_7427_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.18
cc_541 VNB N_A_3799_911#_c_7503_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.735
cc_542 VNB N_A_3799_911#_c_7504_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=2.36
+ $Y2=0.59
cc_543 VNB N_A_3799_911#_c_7505_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=2.705
+ $Y2=0.18
cc_544 VNB N_A_3799_911#_c_7506_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=2.435
+ $Y2=0.18
cc_545 VNB N_A_3799_911#_c_7507_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=2.855
+ $Y2=0.18
cc_546 VNB N_A_3799_911#_c_7508_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=3.545
+ $Y2=0.18
cc_547 VNB N_A_3799_911#_c_7509_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=3.62
+ $Y2=0.59
cc_548 VNB N_A_3799_911#_c_7510_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.09
+ $Y2=0.81
cc_549 VPB N_S[0]_c_904_n 0.0150835f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_550 VPB N_S[0]_c_905_n 0.0395631f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_551 VPB N_S[0]_c_909_n 0.00781808f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_552 VPB N_S[0]_c_929_n 0.0262387f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.55
cc_553 VPB N_S[0]_c_925_n 0.00150672f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_554 VPB N_S[1]_c_1016_n 0.0150835f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_555 VPB N_S[1]_c_1038_n 0.0185487f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_556 VPB N_S[1]_c_1017_n 0.0210144f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=0.735
cc_557 VPB N_S[1]_c_1040_n 0.00863542f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=0.735
cc_558 VPB N_S[1]_c_1019_n 0.00781808f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=0.445
cc_559 VPB N_S[1]_c_1042_n 0.0176033f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.55
cc_560 VPB N_S[1]_c_1036_n 0.00150672f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_561 VPB N_A_142_325#_c_1141_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=0.445
cc_562 VPB N_A_142_325#_c_1142_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0.72 $Y2=0.81
cc_563 VPB N_A_142_325#_c_1134_n 0.0216727f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.735
cc_564 VPB N_A_142_325#_c_1144_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.445
cc_565 VPB N_A_142_325#_c_1145_n 0.013221f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_566 VPB N_A_142_325#_c_1146_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=2.035
cc_567 VPB N_A_142_325#_c_1147_n 0.0312612f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=0.81
cc_568 VPB N_A_142_325#_c_1148_n 0.0215147f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=0.735
cc_569 VPB N_A_142_325#_c_1149_n 0.00800249f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.255
cc_570 VPB N_A_142_325#_c_1150_n 0.00747525f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_571 VPB N_A_142_325#_c_1151_n 0.00751381f $X=-0.19 $Y=1.305 $X2=2.435
+ $Y2=0.18
cc_572 VPB N_A_142_325#_c_1137_n 0.0136355f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.18
cc_573 VPB N_A_142_325#_c_1153_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_574 VPB N_A_142_325#_c_1139_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0.62 $Y2=0.81
cc_575 VPB N_A_142_325#_c_1140_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_576 VPB N_A_142_599#_c_1253_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=0.445
cc_577 VPB N_A_142_599#_c_1254_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0.72 $Y2=0.81
cc_578 VPB N_A_142_599#_c_1246_n 0.0216727f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.735
cc_579 VPB N_A_142_599#_c_1256_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.445
cc_580 VPB N_A_142_599#_c_1257_n 0.013221f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_581 VPB N_A_142_599#_c_1258_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=2.035
cc_582 VPB N_A_142_599#_c_1259_n 0.0312612f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=0.81
cc_583 VPB N_A_142_599#_c_1260_n 0.0215147f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=0.735
cc_584 VPB N_A_142_599#_c_1261_n 0.00800249f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.255
cc_585 VPB N_A_142_599#_c_1262_n 0.00747525f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_586 VPB N_A_142_599#_c_1263_n 0.0021116f $X=-0.19 $Y=1.305 $X2=2.435 $Y2=0.18
cc_587 VPB N_A_142_599#_c_1264_n 0.00195069f $X=-0.19 $Y=1.305 $X2=3.2 $Y2=0.59
cc_588 VPB N_A_142_599#_c_1249_n 0.0136355f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.18
cc_589 VPB N_A_142_599#_c_1266_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_590 VPB N_A_142_599#_c_1251_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0.62 $Y2=0.81
cc_591 VPB N_A_142_599#_c_1252_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_592 VPB N_D[0]_M1012_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_593 VPB N_D[0]_M1049_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_594 VPB N_D[0]_M1086_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.81
cc_595 VPB N_D[0]_M1137_g 0.0187623f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_596 VPB N_D[0]_c_1374_n 0.00769922f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_597 VPB N_D[1]_M1017_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_598 VPB N_D[1]_M1055_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_599 VPB N_D[1]_M1093_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.81
cc_600 VPB N_D[1]_M1141_g 0.0187623f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_601 VPB N_D[1]_c_1473_n 0.00769922f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_602 VPB N_D[2]_M1071_g 0.0187623f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_603 VPB N_D[2]_M1090_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_604 VPB N_D[2]_M1118_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.81
cc_605 VPB N_D[2]_M1158_g 0.0259085f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_606 VPB N_D[2]_c_1570_n 0.00769922f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_607 VPB N_D[3]_M1000_g 0.0187623f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_608 VPB N_D[3]_M1076_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_609 VPB N_D[3]_M1095_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.81
cc_610 VPB N_D[3]_M1120_g 0.0259085f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_611 VPB N_D[3]_c_1671_n 0.00769922f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_612 VPB N_A_1755_265#_c_1765_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=0.445
cc_613 VPB N_A_1755_265#_c_1766_n 0.0145708f $X=-0.19 $Y=1.305 $X2=0.72 $Y2=0.81
cc_614 VPB N_A_1755_265#_c_1767_n 0.0166904f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.735
cc_615 VPB N_A_1755_265#_c_1768_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.445
cc_616 VPB N_A_1755_265#_c_1769_n 0.013221f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_617 VPB N_A_1755_265#_c_1770_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_618 VPB N_A_1755_265#_c_1771_n 0.0140434f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=0.81
cc_619 VPB N_A_1755_265#_c_1772_n 0.0231078f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=0.735
cc_620 VPB N_A_1755_265#_c_1773_n 0.00747525f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.255
cc_621 VPB N_A_1755_265#_c_1774_n 0.00800249f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.59
cc_622 VPB N_A_1755_265#_c_1758_n 0.00733901f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.59
cc_623 VPB N_A_1755_265#_c_1759_n 0.0150864f $X=-0.19 $Y=1.305 $X2=2.855
+ $Y2=0.18
cc_624 VPB N_A_1755_265#_c_1777_n 0.00751381f $X=-0.19 $Y=1.305 $X2=2.78
+ $Y2=0.18
cc_625 VPB N_A_1755_265#_c_1763_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_626 VPB N_A_1755_265#_c_1779_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0.62
+ $Y2=0.81
cc_627 VPB N_A_1755_265#_c_1764_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_628 VPB N_A_1755_793#_c_1884_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=0.445
cc_629 VPB N_A_1755_793#_c_1885_n 0.0145708f $X=-0.19 $Y=1.305 $X2=0.72 $Y2=0.81
cc_630 VPB N_A_1755_793#_c_1886_n 0.0166904f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.735
cc_631 VPB N_A_1755_793#_c_1887_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.445
cc_632 VPB N_A_1755_793#_c_1888_n 0.013221f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_633 VPB N_A_1755_793#_c_1889_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_634 VPB N_A_1755_793#_c_1890_n 0.0140434f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=0.81
cc_635 VPB N_A_1755_793#_c_1891_n 0.0231078f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=0.735
cc_636 VPB N_A_1755_793#_c_1892_n 0.00747525f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.255
cc_637 VPB N_A_1755_793#_c_1893_n 0.00800249f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.59
cc_638 VPB N_A_1755_793#_c_1877_n 0.00733901f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.59
cc_639 VPB N_A_1755_793#_c_1878_n 0.0150864f $X=-0.19 $Y=1.305 $X2=2.855
+ $Y2=0.18
cc_640 VPB N_A_1755_793#_c_1896_n 0.0021116f $X=-0.19 $Y=1.305 $X2=3.2 $Y2=0.59
cc_641 VPB N_A_1755_793#_c_1897_n 0.00195069f $X=-0.19 $Y=1.305 $X2=3.62
+ $Y2=0.255
cc_642 VPB N_A_1755_793#_c_1898_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_643 VPB N_A_1755_793#_c_1881_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_644 VPB N_A_1755_793#_c_1883_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_645 VPB N_S[2]_c_2014_n 0.00781808f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_646 VPB N_S[2]_c_2025_n 0.0260812f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_647 VPB N_S[2]_c_2018_n 0.0526479f $X=-0.19 $Y=1.305 $X2=3.545 $Y2=0.18
cc_648 VPB S[2] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.18
cc_649 VPB N_S[3]_c_2140_n 0.00847786f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.255
cc_650 VPB N_S[3]_c_2131_n 0.00781808f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_651 VPB N_S[3]_c_2142_n 0.0176033f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_652 VPB N_S[3]_c_2134_n 0.0340992f $X=-0.19 $Y=1.305 $X2=3.2 $Y2=0.255
cc_653 VPB N_S[3]_c_2144_n 0.0185487f $X=-0.19 $Y=1.305 $X2=3.545 $Y2=0.18
cc_654 VPB S[3] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.18
cc_655 VPB N_S[4]_c_2244_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_656 VPB N_S[4]_c_2245_n 0.0394096f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_657 VPB N_S[4]_c_2249_n 0.00781808f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_658 VPB N_S[4]_c_2269_n 0.0260812f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.55
cc_659 VPB N_S[4]_c_2265_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_660 VPB N_S[5]_c_2364_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_661 VPB N_S[5]_c_2386_n 0.0185487f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_662 VPB N_S[5]_c_2365_n 0.0208609f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=0.735
cc_663 VPB N_S[5]_c_2388_n 0.00847786f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=0.735
cc_664 VPB N_S[5]_c_2367_n 0.00781808f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=0.445
cc_665 VPB N_S[5]_c_2390_n 0.0176033f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.55
cc_666 VPB N_S[5]_c_2384_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_667 VPB N_A_2626_325#_c_2499_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=0.445
cc_668 VPB N_A_2626_325#_c_2500_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0.72 $Y2=0.81
cc_669 VPB N_A_2626_325#_c_2492_n 0.0215299f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.735
cc_670 VPB N_A_2626_325#_c_2502_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.445
cc_671 VPB N_A_2626_325#_c_2503_n 0.013221f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_672 VPB N_A_2626_325#_c_2504_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_673 VPB N_A_2626_325#_c_2505_n 0.0312612f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=0.81
cc_674 VPB N_A_2626_325#_c_2506_n 0.0215147f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=0.735
cc_675 VPB N_A_2626_325#_c_2507_n 0.00800249f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.255
cc_676 VPB N_A_2626_325#_c_2508_n 0.00747525f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.59
cc_677 VPB N_A_2626_325#_c_2509_n 0.00751381f $X=-0.19 $Y=1.305 $X2=2.435
+ $Y2=0.18
cc_678 VPB N_A_2626_325#_c_2495_n 0.00733901f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.18
cc_679 VPB N_A_2626_325#_c_2511_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_680 VPB N_A_2626_325#_c_2497_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0.62
+ $Y2=0.81
cc_681 VPB N_A_2626_325#_c_2498_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_682 VPB N_A_2626_599#_c_2615_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=0.445
cc_683 VPB N_A_2626_599#_c_2616_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0.72 $Y2=0.81
cc_684 VPB N_A_2626_599#_c_2608_n 0.0215299f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.735
cc_685 VPB N_A_2626_599#_c_2618_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.445
cc_686 VPB N_A_2626_599#_c_2619_n 0.013221f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_687 VPB N_A_2626_599#_c_2620_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_688 VPB N_A_2626_599#_c_2621_n 0.0312612f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=0.81
cc_689 VPB N_A_2626_599#_c_2622_n 0.0215147f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=0.735
cc_690 VPB N_A_2626_599#_c_2623_n 0.00800249f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.255
cc_691 VPB N_A_2626_599#_c_2624_n 0.00747525f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.59
cc_692 VPB N_A_2626_599#_c_2625_n 0.0021116f $X=-0.19 $Y=1.305 $X2=2.435
+ $Y2=0.18
cc_693 VPB N_A_2626_599#_c_2626_n 0.00195069f $X=-0.19 $Y=1.305 $X2=3.2 $Y2=0.59
cc_694 VPB N_A_2626_599#_c_2611_n 0.00733901f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.18
cc_695 VPB N_A_2626_599#_c_2628_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_696 VPB N_A_2626_599#_c_2613_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0.62
+ $Y2=0.81
cc_697 VPB N_A_2626_599#_c_2614_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_698 VPB N_D[4]_M1042_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_699 VPB N_D[4]_M1062_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_700 VPB N_D[4]_M1105_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.81
cc_701 VPB N_D[4]_M1127_g 0.0187623f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_702 VPB N_D[4]_c_2740_n 0.00769922f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_703 VPB N_D[5]_M1046_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_704 VPB N_D[5]_M1070_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_705 VPB N_D[5]_M1113_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.81
cc_706 VPB N_D[5]_M1134_g 0.0187623f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_707 VPB N_D[5]_c_2839_n 0.00769922f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_708 VPB N_D[6]_M1082_g 0.0187623f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_709 VPB N_D[6]_M1108_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_710 VPB N_D[6]_M1130_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.81
cc_711 VPB N_D[6]_M1145_g 0.0259085f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_712 VPB N_D[6]_c_2936_n 0.00769922f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_713 VPB N_D[7]_M1087_g 0.0187623f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.55
cc_714 VPB N_D[7]_M1117_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_715 VPB N_D[7]_M1139_g 0.0177422f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.81
cc_716 VPB N_D[7]_M1153_g 0.0259085f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_717 VPB N_D[7]_c_3037_n 0.00769922f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_718 VPB N_A_4239_265#_c_3131_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=0.445
cc_719 VPB N_A_4239_265#_c_3132_n 0.0145708f $X=-0.19 $Y=1.305 $X2=0.72 $Y2=0.81
cc_720 VPB N_A_4239_265#_c_3133_n 0.0166904f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.735
cc_721 VPB N_A_4239_265#_c_3134_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.445
cc_722 VPB N_A_4239_265#_c_3135_n 0.013221f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_723 VPB N_A_4239_265#_c_3136_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_724 VPB N_A_4239_265#_c_3137_n 0.0140434f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=0.81
cc_725 VPB N_A_4239_265#_c_3138_n 0.0231078f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=0.735
cc_726 VPB N_A_4239_265#_c_3139_n 0.00747525f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.255
cc_727 VPB N_A_4239_265#_c_3140_n 0.00800249f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.59
cc_728 VPB N_A_4239_265#_c_3124_n 0.0136355f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_729 VPB N_A_4239_265#_c_3125_n 0.0150864f $X=-0.19 $Y=1.305 $X2=2.855
+ $Y2=0.18
cc_730 VPB N_A_4239_265#_c_3143_n 0.00751381f $X=-0.19 $Y=1.305 $X2=2.78
+ $Y2=0.18
cc_731 VPB N_A_4239_265#_c_3129_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_732 VPB N_A_4239_265#_c_3145_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0.62
+ $Y2=0.81
cc_733 VPB N_A_4239_265#_c_3130_n 0.0216727f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_734 VPB N_A_4239_793#_c_3246_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0.645
+ $Y2=0.445
cc_735 VPB N_A_4239_793#_c_3247_n 0.0145708f $X=-0.19 $Y=1.305 $X2=0.72 $Y2=0.81
cc_736 VPB N_A_4239_793#_c_3248_n 0.0166904f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.735
cc_737 VPB N_A_4239_793#_c_3249_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.065
+ $Y2=0.445
cc_738 VPB N_A_4239_793#_c_3250_n 0.013221f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.45
cc_739 VPB N_A_4239_793#_c_3251_n 0.0174802f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_740 VPB N_A_4239_793#_c_3252_n 0.0140434f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=0.81
cc_741 VPB N_A_4239_793#_c_3253_n 0.0231078f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=0.735
cc_742 VPB N_A_4239_793#_c_3254_n 0.00747525f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.255
cc_743 VPB N_A_4239_793#_c_3255_n 0.00800249f $X=-0.19 $Y=1.305 $X2=2.36
+ $Y2=0.59
cc_744 VPB N_A_4239_793#_c_3239_n 0.0136355f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_745 VPB N_A_4239_793#_c_3240_n 0.0150864f $X=-0.19 $Y=1.305 $X2=2.855
+ $Y2=0.18
cc_746 VPB N_A_4239_793#_c_3258_n 0.0021116f $X=-0.19 $Y=1.305 $X2=3.2 $Y2=0.59
cc_747 VPB N_A_4239_793#_c_3259_n 0.00195069f $X=-0.19 $Y=1.305 $X2=3.62
+ $Y2=0.255
cc_748 VPB N_A_4239_793#_c_3260_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_749 VPB N_A_4239_793#_c_3243_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_750 VPB N_A_4239_793#_c_3245_n 0.0216727f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_751 VPB N_S[6]_c_3372_n 0.00781808f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_752 VPB N_S[6]_c_3383_n 0.0262387f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_753 VPB N_S[6]_c_3376_n 0.0546486f $X=-0.19 $Y=1.305 $X2=3.545 $Y2=0.18
cc_754 VPB S[6] 0.00150672f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.18
cc_755 VPB N_S[7]_c_3491_n 0.00863542f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.255
cc_756 VPB N_S[7]_c_3482_n 0.00781808f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_757 VPB N_S[7]_c_3493_n 0.0176033f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.59
cc_758 VPB N_S[7]_c_3485_n 0.0361f $X=-0.19 $Y=1.305 $X2=3.2 $Y2=0.255
cc_759 VPB N_S[7]_c_3495_n 0.0185487f $X=-0.19 $Y=1.305 $X2=3.545 $Y2=0.18
cc_760 VPB S[7] 0.00150672f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.18
cc_761 VPB N_VPWR_c_3586_n 0.0422729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_762 VPB N_VPWR_c_3587_n 0.0422729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_763 VPB N_VPWR_c_3588_n 0.0171933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_764 VPB N_VPWR_c_3589_n 0.0171933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_765 VPB N_VPWR_c_3590_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_766 VPB N_VPWR_c_3591_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_767 VPB N_VPWR_c_3592_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_768 VPB N_VPWR_c_3593_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_769 VPB N_VPWR_c_3594_n 0.00446796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_770 VPB N_VPWR_c_3595_n 0.00446796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_771 VPB N_VPWR_c_3596_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_772 VPB N_VPWR_c_3597_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_773 VPB N_VPWR_c_3598_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_774 VPB N_VPWR_c_3599_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_775 VPB N_VPWR_c_3600_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_776 VPB N_VPWR_c_3601_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_777 VPB N_VPWR_c_3602_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_778 VPB N_VPWR_c_3603_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_779 VPB N_VPWR_c_3604_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_780 VPB N_VPWR_c_3605_n 0.013938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_781 VPB N_VPWR_c_3606_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_782 VPB N_VPWR_c_3607_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_783 VPB N_VPWR_c_3608_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_784 VPB N_VPWR_c_3609_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_785 VPB N_VPWR_c_3610_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_786 VPB N_VPWR_c_3611_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_787 VPB N_VPWR_c_3612_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_788 VPB N_VPWR_c_3613_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_789 VPB N_VPWR_c_3614_n 0.00446796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_790 VPB N_VPWR_c_3615_n 0.00446796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_791 VPB N_VPWR_c_3616_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_792 VPB N_VPWR_c_3617_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_793 VPB N_VPWR_c_3618_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_794 VPB N_VPWR_c_3619_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_795 VPB N_VPWR_c_3620_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_796 VPB N_VPWR_c_3621_n 0.0171933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_797 VPB N_VPWR_c_3622_n 0.0171933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_798 VPB N_VPWR_c_3623_n 0.0422729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_799 VPB N_VPWR_c_3624_n 0.0422729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_800 VPB N_VPWR_c_3625_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_801 VPB N_VPWR_c_3626_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_802 VPB N_VPWR_c_3627_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_803 VPB N_VPWR_c_3628_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_804 VPB N_VPWR_c_3629_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_805 VPB N_VPWR_c_3630_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_806 VPB N_VPWR_c_3631_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_807 VPB N_VPWR_c_3632_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_808 VPB N_VPWR_c_3633_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_809 VPB N_VPWR_c_3634_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_810 VPB N_VPWR_c_3635_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_811 VPB N_VPWR_c_3636_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_812 VPB N_VPWR_c_3637_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_813 VPB N_VPWR_c_3638_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_814 VPB N_VPWR_c_3639_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_815 VPB N_VPWR_c_3640_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_816 VPB N_VPWR_c_3641_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_817 VPB N_VPWR_c_3642_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_818 VPB N_VPWR_c_3643_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_819 VPB N_VPWR_c_3644_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_820 VPB N_VPWR_c_3645_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_821 VPB N_VPWR_c_3646_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_822 VPB N_VPWR_c_3647_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_823 VPB N_VPWR_c_3648_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_824 VPB N_VPWR_c_3649_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_825 VPB N_VPWR_c_3650_n 0.0110983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_826 VPB N_VPWR_c_3651_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_827 VPB N_VPWR_c_3652_n 0.00206163f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_828 VPB N_VPWR_c_3653_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_829 VPB N_VPWR_c_3654_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_830 VPB N_VPWR_c_3655_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_831 VPB N_VPWR_c_3656_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_832 VPB N_VPWR_c_3657_n 0.00206163f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_833 VPB N_VPWR_c_3658_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_834 VPB N_VPWR_c_3659_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_835 VPB N_VPWR_c_3660_n 0.0110983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_836 VPB N_VPWR_c_3661_n 0.207817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_837 VPB N_A_355_311#_c_4334_n 0.0075016f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.55
cc_838 VPB N_A_355_311#_c_4335_n 0.00726062f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_839 VPB N_A_355_311#_c_4336_n 0.00219932f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_840 VPB N_A_355_311#_c_4337_n 0.0128471f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_841 VPB N_A_355_311#_c_4338_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_842 VPB N_A_355_311#_c_4339_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_843 VPB N_A_355_613#_c_4461_n 0.0075016f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.55
cc_844 VPB N_A_355_613#_c_4462_n 0.00726062f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_845 VPB N_A_355_613#_c_4463_n 0.00219932f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.59
cc_846 VPB N_A_355_613#_c_4464_n 0.0128471f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_847 VPB N_A_355_613#_c_4465_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_848 VPB N_A_355_613#_c_4466_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_849 VPB N_Z_c_4610_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_850 VPB N_Z_c_4611_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_851 VPB N_Z_c_4618_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_852 VPB N_Z_c_4619_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_853 VPB N_Z_c_4624_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_854 VPB N_Z_c_4625_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_855 VPB N_Z_c_4632_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_856 VPB N_Z_c_4633_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_857 VPB N_Z_c_4644_n 0.0070095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_858 VPB N_Z_c_4645_n 0.0070095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_859 VPB N_Z_c_4646_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_860 VPB N_Z_c_4647_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_861 VPB N_Z_c_4648_n 0.0070095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_862 VPB N_Z_c_4649_n 0.0070095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_863 VPB N_Z_c_4650_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_864 VPB N_Z_c_4651_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_865 VPB N_Z_c_4652_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_866 VPB N_Z_c_4653_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_867 VPB N_Z_c_4654_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_868 VPB N_Z_c_4655_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_869 VPB N_Z_c_4656_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_870 VPB N_Z_c_4657_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_871 VPB N_A_1313_297#_c_5502_n 0.0147622f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_872 VPB N_A_1313_297#_c_5503_n 0.00219932f $X=-0.19 $Y=1.305 $X2=2.435
+ $Y2=0.18
cc_873 VPB N_A_1313_297#_c_5504_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_874 VPB N_A_1313_297#_c_5505_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_875 VPB N_A_1313_297#_c_5506_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_876 VPB N_A_1313_591#_c_5630_n 0.0147622f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_877 VPB N_A_1313_591#_c_5631_n 0.00219932f $X=-0.19 $Y=1.305 $X2=2.435
+ $Y2=0.18
cc_878 VPB N_A_1313_591#_c_5632_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_879 VPB N_A_1313_591#_c_5633_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_880 VPB N_A_1313_591#_c_5634_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_881 VPB N_A_2839_311#_c_5758_n 0.0075016f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.55
cc_882 VPB N_A_2839_311#_c_5759_n 0.00726062f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_883 VPB N_A_2839_311#_c_5760_n 0.00219932f $X=-0.19 $Y=1.305 $X2=2.78
+ $Y2=0.59
cc_884 VPB N_A_2839_311#_c_5761_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_885 VPB N_A_2839_311#_c_5762_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_886 VPB N_A_2839_311#_c_5763_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_887 VPB N_A_2839_613#_c_5889_n 0.0075016f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.55
cc_888 VPB N_A_2839_613#_c_5890_n 0.00726062f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_889 VPB N_A_2839_613#_c_5891_n 0.00219932f $X=-0.19 $Y=1.305 $X2=2.78
+ $Y2=0.59
cc_890 VPB N_A_2839_613#_c_5892_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_891 VPB N_A_2839_613#_c_5893_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_892 VPB N_A_2839_613#_c_5894_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_893 VPB N_A_3797_297#_c_6020_n 0.0147622f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_894 VPB N_A_3797_297#_c_6021_n 0.00219932f $X=-0.19 $Y=1.305 $X2=2.435
+ $Y2=0.18
cc_895 VPB N_A_3797_297#_c_6022_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_896 VPB N_A_3797_297#_c_6023_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_897 VPB N_A_3797_297#_c_6024_n 0.0128471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_898 VPB N_A_3797_591#_c_6142_n 0.0147622f $X=-0.19 $Y=1.305 $X2=1.09
+ $Y2=2.035
cc_899 VPB N_A_3797_591#_c_6143_n 0.00219932f $X=-0.19 $Y=1.305 $X2=2.435
+ $Y2=0.18
cc_900 VPB N_A_3797_591#_c_6144_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_901 VPB N_A_3797_591#_c_6145_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_902 VPB N_A_3797_591#_c_6146_n 0.0128471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_903 N_S[0]_c_905_n N_S[1]_c_1038_n 0.0130744f $X=0.62 $Y=1.55 $X2=0 $Y2=0
cc_904 N_S[0]_c_929_n N_S[1]_c_1042_n 0.0130744f $X=1.09 $Y=1.55 $X2=0 $Y2=0
cc_905 N_S[0]_c_914_n N_A_142_325#_c_1142_n 0.00507688f $X=2.36 $Y=0.255 $X2=0
+ $Y2=0
cc_906 N_S[0]_c_909_n N_A_142_325#_c_1134_n 0.00262132f $X=1.09 $Y=1.45 $X2=0
+ $Y2=0
cc_907 N_S[0]_c_916_n N_A_142_325#_c_1145_n 0.00509204f $X=2.78 $Y=0.255 $X2=0
+ $Y2=0
cc_908 N_S[0]_c_920_n N_A_142_325#_c_1147_n 0.00507426f $X=3.62 $Y=0.255 $X2=0
+ $Y2=0
cc_909 N_S[0]_c_918_n N_A_142_325#_c_1150_n 0.00509391f $X=3.2 $Y=0.255 $X2=0
+ $Y2=0
cc_910 N_S[0]_c_905_n N_A_142_325#_c_1151_n 0.0133753f $X=0.62 $Y=1.55 $X2=0
+ $Y2=0
cc_911 N_S[0]_c_929_n N_A_142_325#_c_1151_n 0.0123982f $X=1.09 $Y=1.55 $X2=0
+ $Y2=0
cc_912 N_S[0]_c_906_n N_A_142_325#_c_1135_n 0.00207203f $X=0.645 $Y=0.735 $X2=0
+ $Y2=0
cc_913 N_S[0]_c_908_n N_A_142_325#_c_1135_n 0.00603996f $X=1.065 $Y=0.735 $X2=0
+ $Y2=0
cc_914 N_S[0]_c_911_n N_A_142_325#_c_1135_n 6.53442e-19 $X=1.6 $Y=0.735 $X2=0
+ $Y2=0
cc_915 N_S[0]_c_905_n N_A_142_325#_c_1136_n 0.00289358f $X=0.62 $Y=1.55 $X2=0
+ $Y2=0
cc_916 N_S[0]_c_907_n N_A_142_325#_c_1136_n 0.00429801f $X=0.99 $Y=0.81 $X2=0
+ $Y2=0
cc_917 N_S[0]_c_909_n N_A_142_325#_c_1136_n 0.0085951f $X=1.09 $Y=1.45 $X2=0
+ $Y2=0
cc_918 N_S[0]_c_921_n N_A_142_325#_c_1136_n 0.00268644f $X=1.09 $Y=0.81 $X2=0
+ $Y2=0
cc_919 N_S[0]_c_925_n N_A_142_325#_c_1136_n 0.00541767f $X=0.58 $Y=1.16 $X2=0
+ $Y2=0
cc_920 N_S[0]_c_909_n N_A_142_325#_c_1137_n 0.0250056f $X=1.09 $Y=1.45 $X2=0
+ $Y2=0
cc_921 N_S[0]_c_910_n N_A_142_325#_c_1137_n 0.0103812f $X=1.525 $Y=0.81 $X2=0
+ $Y2=0
cc_922 N_S[0]_c_905_n N_A_142_325#_c_1153_n 0.00454075f $X=0.62 $Y=1.55 $X2=0
+ $Y2=0
cc_923 N_S[0]_c_909_n N_A_142_325#_c_1153_n 0.00255921f $X=1.09 $Y=1.45 $X2=0
+ $Y2=0
cc_924 N_S[0]_c_929_n N_A_142_325#_c_1153_n 0.00762115f $X=1.09 $Y=1.55 $X2=0
+ $Y2=0
cc_925 N_S[0]_c_907_n N_A_142_325#_c_1138_n 0.0111895f $X=0.99 $Y=0.81 $X2=0
+ $Y2=0
cc_926 N_S[0]_c_908_n N_A_142_325#_c_1138_n 9.67113e-19 $X=1.065 $Y=0.735 $X2=0
+ $Y2=0
cc_927 N_S[0]_c_921_n N_A_142_325#_c_1138_n 0.00426435f $X=1.09 $Y=0.81 $X2=0
+ $Y2=0
cc_928 N_S[0]_c_905_n N_A_142_325#_c_1139_n 0.00416423f $X=0.62 $Y=1.55 $X2=0
+ $Y2=0
cc_929 N_S[0]_c_909_n N_A_142_325#_c_1139_n 0.00322131f $X=1.09 $Y=1.45 $X2=0
+ $Y2=0
cc_930 N_S[0]_c_925_n N_A_142_325#_c_1139_n 0.0228692f $X=0.58 $Y=1.16 $X2=0
+ $Y2=0
cc_931 N_S[0]_c_909_n N_A_142_325#_c_1140_n 0.0175393f $X=1.09 $Y=1.45 $X2=0
+ $Y2=0
cc_932 N_S[0]_c_910_n N_A_142_325#_c_1140_n 0.0179529f $X=1.525 $Y=0.81 $X2=0
+ $Y2=0
cc_933 N_S[0]_c_904_n N_VPWR_c_3586_n 0.00652399f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_934 N_S[0]_c_905_n N_VPWR_c_3586_n 0.00966078f $X=0.62 $Y=1.55 $X2=0 $Y2=0
cc_935 N_S[0]_c_925_n N_VPWR_c_3586_n 0.017333f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_936 N_S[0]_c_929_n N_VPWR_c_3588_n 0.00929376f $X=1.09 $Y=1.55 $X2=0 $Y2=0
cc_937 N_S[0]_c_905_n N_VPWR_c_3626_n 0.0035837f $X=0.62 $Y=1.55 $X2=0 $Y2=0
cc_938 N_S[0]_c_929_n N_VPWR_c_3626_n 0.0035837f $X=1.09 $Y=1.55 $X2=0 $Y2=0
cc_939 N_S[0]_c_905_n N_VPWR_c_3661_n 0.0114704f $X=0.62 $Y=1.55 $X2=0 $Y2=0
cc_940 N_S[0]_c_929_n N_VPWR_c_3661_n 0.0118174f $X=1.09 $Y=1.55 $X2=0 $Y2=0
cc_941 N_S[0]_c_920_n N_A_355_311#_c_4335_n 0.00168571f $X=3.62 $Y=0.255 $X2=0
+ $Y2=0
cc_942 N_S[0]_c_929_n N_A_355_311#_c_4337_n 0.00249814f $X=1.09 $Y=1.55 $X2=0
+ $Y2=0
cc_943 N_S[0]_c_914_n N_Z_c_4588_n 0.0134253f $X=2.36 $Y=0.255 $X2=0 $Y2=0
cc_944 N_S[0]_c_916_n N_Z_c_4588_n 0.0077801f $X=2.78 $Y=0.255 $X2=0 $Y2=0
cc_945 N_S[0]_c_918_n N_Z_c_4588_n 6.35774e-19 $X=3.2 $Y=0.255 $X2=0 $Y2=0
cc_946 N_S[0]_c_916_n N_Z_c_4590_n 0.00190704f $X=2.78 $Y=0.255 $X2=0 $Y2=0
cc_947 N_S[0]_c_918_n N_Z_c_4590_n 3.10191e-19 $X=3.2 $Y=0.255 $X2=0 $Y2=0
cc_948 N_S[0]_c_918_n N_Z_c_4592_n 0.00283489f $X=3.2 $Y=0.255 $X2=0 $Y2=0
cc_949 N_S[0]_c_920_n N_Z_c_4592_n 0.002324f $X=3.62 $Y=0.255 $X2=0 $Y2=0
cc_950 N_S[0]_c_914_n N_Z_c_4608_n 0.00216436f $X=2.36 $Y=0.255 $X2=0 $Y2=0
cc_951 N_S[0]_c_918_n N_Z_c_4610_n 0.00180363f $X=3.2 $Y=0.255 $X2=0 $Y2=0
cc_952 N_S[0]_c_916_n N_Z_c_4612_n 6.35664e-19 $X=2.78 $Y=0.255 $X2=0 $Y2=0
cc_953 N_S[0]_c_918_n N_Z_c_4612_n 0.00462308f $X=3.2 $Y=0.255 $X2=0 $Y2=0
cc_954 N_S[0]_c_920_n N_Z_c_4612_n 0.00443615f $X=3.62 $Y=0.255 $X2=0 $Y2=0
cc_955 N_S[0]_c_904_n N_VGND_c_6265_n 0.00576464f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_956 N_S[0]_c_906_n N_VGND_c_6265_n 0.00374526f $X=0.645 $Y=0.735 $X2=0 $Y2=0
cc_957 N_S[0]_c_925_n N_VGND_c_6265_n 0.0116218f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_958 N_S[0]_c_908_n N_VGND_c_6268_n 0.00173127f $X=1.065 $Y=0.735 $X2=0 $Y2=0
cc_959 N_S[0]_c_910_n N_VGND_c_6268_n 0.00525833f $X=1.525 $Y=0.81 $X2=0 $Y2=0
cc_960 N_S[0]_c_913_n N_VGND_c_6268_n 0.00862298f $X=1.675 $Y=0.18 $X2=0 $Y2=0
cc_961 N_S[0]_c_919_n N_VGND_c_6270_n 0.0028166f $X=3.545 $Y=0.18 $X2=0 $Y2=0
cc_962 N_S[0]_c_920_n N_VGND_c_6270_n 5.5039e-19 $X=3.62 $Y=0.255 $X2=0 $Y2=0
cc_963 N_S[0]_c_906_n N_VGND_c_6308_n 0.00585385f $X=0.645 $Y=0.735 $X2=0 $Y2=0
cc_964 N_S[0]_c_907_n N_VGND_c_6308_n 2.16067e-19 $X=0.99 $Y=0.81 $X2=0 $Y2=0
cc_965 N_S[0]_c_908_n N_VGND_c_6308_n 0.00542362f $X=1.065 $Y=0.735 $X2=0 $Y2=0
cc_966 N_S[0]_c_913_n N_VGND_c_6312_n 0.0559651f $X=1.675 $Y=0.18 $X2=0 $Y2=0
cc_967 N_S[0]_c_906_n N_VGND_c_6370_n 0.0117149f $X=0.645 $Y=0.735 $X2=0 $Y2=0
cc_968 N_S[0]_c_908_n N_VGND_c_6370_n 0.00990284f $X=1.065 $Y=0.735 $X2=0 $Y2=0
cc_969 N_S[0]_c_912_n N_VGND_c_6370_n 0.0244174f $X=2.285 $Y=0.18 $X2=0 $Y2=0
cc_970 N_S[0]_c_913_n N_VGND_c_6370_n 0.0101627f $X=1.675 $Y=0.18 $X2=0 $Y2=0
cc_971 N_S[0]_c_915_n N_VGND_c_6370_n 0.00642387f $X=2.705 $Y=0.18 $X2=0 $Y2=0
cc_972 N_S[0]_c_917_n N_VGND_c_6370_n 0.0064237f $X=3.125 $Y=0.18 $X2=0 $Y2=0
cc_973 N_S[0]_c_919_n N_VGND_c_6370_n 0.0123437f $X=3.545 $Y=0.18 $X2=0 $Y2=0
cc_974 N_S[0]_c_922_n N_VGND_c_6370_n 0.00366655f $X=2.36 $Y=0.18 $X2=0 $Y2=0
cc_975 N_S[0]_c_923_n N_VGND_c_6370_n 0.00366655f $X=2.78 $Y=0.18 $X2=0 $Y2=0
cc_976 N_S[0]_c_924_n N_VGND_c_6370_n 0.00366655f $X=3.2 $Y=0.18 $X2=0 $Y2=0
cc_977 N_S[0]_c_911_n N_A_405_66#_c_6926_n 0.00529837f $X=1.6 $Y=0.735 $X2=0
+ $Y2=0
cc_978 N_S[0]_c_914_n N_A_405_66#_c_6927_n 0.0112916f $X=2.36 $Y=0.255 $X2=0
+ $Y2=0
cc_979 N_S[0]_c_915_n N_A_405_66#_c_6927_n 0.00211351f $X=2.705 $Y=0.18 $X2=0
+ $Y2=0
cc_980 N_S[0]_c_916_n N_A_405_66#_c_6927_n 0.0106844f $X=2.78 $Y=0.255 $X2=0
+ $Y2=0
cc_981 N_S[0]_c_911_n N_A_405_66#_c_6928_n 0.00189496f $X=1.6 $Y=0.735 $X2=0
+ $Y2=0
cc_982 N_S[0]_c_912_n N_A_405_66#_c_6928_n 0.00685838f $X=2.285 $Y=0.18 $X2=0
+ $Y2=0
cc_983 N_S[0]_c_918_n N_A_405_66#_c_6929_n 0.0106826f $X=3.2 $Y=0.255 $X2=0
+ $Y2=0
cc_984 N_S[0]_c_919_n N_A_405_66#_c_6929_n 0.00211351f $X=3.545 $Y=0.18 $X2=0
+ $Y2=0
cc_985 N_S[0]_c_920_n N_A_405_66#_c_6929_n 0.0139014f $X=3.62 $Y=0.255 $X2=0
+ $Y2=0
cc_986 N_S[0]_c_920_n N_A_405_66#_c_6932_n 0.00206084f $X=3.62 $Y=0.255 $X2=0
+ $Y2=0
cc_987 N_S[0]_c_917_n N_A_405_66#_c_6945_n 0.0034777f $X=3.125 $Y=0.18 $X2=0
+ $Y2=0
cc_988 N_S[1]_c_1025_n N_A_142_599#_c_1254_n 0.00507688f $X=2.36 $Y=5.185 $X2=0
+ $Y2=0
cc_989 N_S[1]_c_1040_n N_A_142_599#_c_1246_n 0.00262132f $X=1.09 $Y=3.99 $X2=0
+ $Y2=0
cc_990 N_S[1]_c_1027_n N_A_142_599#_c_1257_n 0.00509204f $X=2.78 $Y=5.185 $X2=0
+ $Y2=0
cc_991 N_S[1]_c_1031_n N_A_142_599#_c_1259_n 0.00507426f $X=3.62 $Y=5.185 $X2=0
+ $Y2=0
cc_992 N_S[1]_c_1029_n N_A_142_599#_c_1262_n 0.00509391f $X=3.2 $Y=5.185 $X2=0
+ $Y2=0
cc_993 N_S[1]_c_1038_n N_A_142_599#_c_1263_n 0.0097833f $X=0.62 $Y=3.89 $X2=0
+ $Y2=0
cc_994 N_S[1]_c_1042_n N_A_142_599#_c_1263_n 0.010234f $X=1.09 $Y=3.89 $X2=0
+ $Y2=0
cc_995 N_S[1]_c_1017_n N_A_142_599#_c_1247_n 0.00207203f $X=0.645 $Y=4.705 $X2=0
+ $Y2=0
cc_996 N_S[1]_c_1018_n N_A_142_599#_c_1247_n 0.0111895f $X=0.99 $Y=4.63 $X2=0
+ $Y2=0
cc_997 N_S[1]_c_1020_n N_A_142_599#_c_1247_n 9.67113e-19 $X=1.065 $Y=4.705 $X2=0
+ $Y2=0
cc_998 N_S[1]_c_1022_n N_A_142_599#_c_1247_n 6.53442e-19 $X=1.6 $Y=5.185 $X2=0
+ $Y2=0
cc_999 N_S[1]_c_1032_n N_A_142_599#_c_1247_n 0.00426435f $X=1.09 $Y=4.63 $X2=0
+ $Y2=0
cc_1000 N_S[1]_c_1020_n N_A_142_599#_c_1248_n 0.00603996f $X=1.065 $Y=4.705
+ $X2=0 $Y2=0
cc_1001 N_S[1]_c_1038_n N_A_142_599#_c_1264_n 0.00117303f $X=0.62 $Y=3.89 $X2=0
+ $Y2=0
cc_1002 N_S[1]_c_1017_n N_A_142_599#_c_1264_n 0.00336772f $X=0.645 $Y=4.705
+ $X2=0 $Y2=0
cc_1003 N_S[1]_c_1040_n N_A_142_599#_c_1264_n 0.00508008f $X=1.09 $Y=3.99 $X2=0
+ $Y2=0
cc_1004 N_S[1]_c_1019_n N_A_142_599#_c_1264_n 0.00255921f $X=1.09 $Y=4.555 $X2=0
+ $Y2=0
cc_1005 N_S[1]_c_1042_n N_A_142_599#_c_1264_n 0.00254107f $X=1.09 $Y=3.89 $X2=0
+ $Y2=0
cc_1006 N_S[1]_c_1019_n N_A_142_599#_c_1249_n 0.0250056f $X=1.09 $Y=4.555 $X2=0
+ $Y2=0
cc_1007 N_S[1]_c_1021_n N_A_142_599#_c_1249_n 0.0103812f $X=1.525 $Y=4.63 $X2=0
+ $Y2=0
cc_1008 N_S[1]_c_1038_n N_A_142_599#_c_1266_n 0.00304348f $X=0.62 $Y=3.89 $X2=0
+ $Y2=0
cc_1009 N_S[1]_c_1017_n N_A_142_599#_c_1266_n 5.48523e-19 $X=0.645 $Y=4.705
+ $X2=0 $Y2=0
cc_1010 N_S[1]_c_1042_n N_A_142_599#_c_1266_n 0.00216424f $X=1.09 $Y=3.89 $X2=0
+ $Y2=0
cc_1011 N_S[1]_c_1017_n N_A_142_599#_c_1250_n 0.00289358f $X=0.645 $Y=4.705
+ $X2=0 $Y2=0
cc_1012 N_S[1]_c_1018_n N_A_142_599#_c_1250_n 0.00429801f $X=0.99 $Y=4.63 $X2=0
+ $Y2=0
cc_1013 N_S[1]_c_1019_n N_A_142_599#_c_1250_n 0.0085951f $X=1.09 $Y=4.555 $X2=0
+ $Y2=0
cc_1014 N_S[1]_c_1032_n N_A_142_599#_c_1250_n 0.00268644f $X=1.09 $Y=4.63 $X2=0
+ $Y2=0
cc_1015 N_S[1]_c_1036_n N_A_142_599#_c_1250_n 0.00541767f $X=0.58 $Y=4.28 $X2=0
+ $Y2=0
cc_1016 N_S[1]_c_1017_n N_A_142_599#_c_1251_n 0.00416423f $X=0.645 $Y=4.705
+ $X2=0 $Y2=0
cc_1017 N_S[1]_c_1019_n N_A_142_599#_c_1251_n 0.00322131f $X=1.09 $Y=4.555 $X2=0
+ $Y2=0
cc_1018 N_S[1]_c_1036_n N_A_142_599#_c_1251_n 0.0228692f $X=0.58 $Y=4.28 $X2=0
+ $Y2=0
cc_1019 N_S[1]_c_1019_n N_A_142_599#_c_1252_n 0.0175393f $X=1.09 $Y=4.555 $X2=0
+ $Y2=0
cc_1020 N_S[1]_c_1021_n N_A_142_599#_c_1252_n 0.0179529f $X=1.525 $Y=4.63 $X2=0
+ $Y2=0
cc_1021 N_S[1]_c_1016_n N_VPWR_c_3587_n 0.00652399f $X=0.52 $Y=4.28 $X2=0 $Y2=0
cc_1022 N_S[1]_c_1038_n N_VPWR_c_3587_n 0.00966078f $X=0.62 $Y=3.89 $X2=0 $Y2=0
cc_1023 N_S[1]_c_1036_n N_VPWR_c_3587_n 0.017333f $X=0.58 $Y=4.28 $X2=0 $Y2=0
cc_1024 N_S[1]_c_1042_n N_VPWR_c_3589_n 0.00929376f $X=1.09 $Y=3.89 $X2=0 $Y2=0
cc_1025 N_S[1]_c_1038_n N_VPWR_c_3626_n 0.0035837f $X=0.62 $Y=3.89 $X2=0 $Y2=0
cc_1026 N_S[1]_c_1042_n N_VPWR_c_3626_n 0.0035837f $X=1.09 $Y=3.89 $X2=0 $Y2=0
cc_1027 N_S[1]_c_1038_n N_VPWR_c_3661_n 0.0114704f $X=0.62 $Y=3.89 $X2=0 $Y2=0
cc_1028 N_S[1]_c_1042_n N_VPWR_c_3661_n 0.0118174f $X=1.09 $Y=3.89 $X2=0 $Y2=0
cc_1029 N_S[1]_c_1031_n N_A_355_613#_c_4462_n 0.00168571f $X=3.62 $Y=5.185 $X2=0
+ $Y2=0
cc_1030 N_S[1]_c_1042_n N_A_355_613#_c_4464_n 0.00249814f $X=1.09 $Y=3.89 $X2=0
+ $Y2=0
cc_1031 N_S[1]_c_1025_n N_Z_c_4589_n 0.0134253f $X=2.36 $Y=5.185 $X2=0 $Y2=0
cc_1032 N_S[1]_c_1027_n N_Z_c_4589_n 0.0077801f $X=2.78 $Y=5.185 $X2=0 $Y2=0
cc_1033 N_S[1]_c_1029_n N_Z_c_4589_n 6.35774e-19 $X=3.2 $Y=5.185 $X2=0 $Y2=0
cc_1034 N_S[1]_c_1027_n N_Z_c_4591_n 0.00190704f $X=2.78 $Y=5.185 $X2=0 $Y2=0
cc_1035 N_S[1]_c_1029_n N_Z_c_4591_n 3.10191e-19 $X=3.2 $Y=5.185 $X2=0 $Y2=0
cc_1036 N_S[1]_c_1025_n N_Z_c_4609_n 0.00216436f $X=2.36 $Y=5.185 $X2=0 $Y2=0
cc_1037 N_S[1]_c_1029_n N_Z_c_4611_n 0.00180363f $X=3.2 $Y=5.185 $X2=0 $Y2=0
cc_1038 N_S[1]_c_1029_n N_Z_c_4613_n 0.00462308f $X=3.2 $Y=5.185 $X2=0 $Y2=0
cc_1039 N_S[1]_c_1031_n N_Z_c_4613_n 0.00443615f $X=3.62 $Y=5.185 $X2=0 $Y2=0
cc_1040 N_S[1]_c_1027_n N_Z_c_4614_n 6.35664e-19 $X=2.78 $Y=5.185 $X2=0 $Y2=0
cc_1041 N_S[1]_c_1029_n N_Z_c_4614_n 0.00283489f $X=3.2 $Y=5.185 $X2=0 $Y2=0
cc_1042 N_S[1]_c_1031_n N_Z_c_4614_n 0.002324f $X=3.62 $Y=5.185 $X2=0 $Y2=0
cc_1043 N_S[1]_c_1016_n N_VGND_c_6267_n 0.00576464f $X=0.52 $Y=4.28 $X2=0 $Y2=0
cc_1044 N_S[1]_c_1017_n N_VGND_c_6267_n 0.00374526f $X=0.645 $Y=4.705 $X2=0
+ $Y2=0
cc_1045 N_S[1]_c_1036_n N_VGND_c_6267_n 0.0116218f $X=0.58 $Y=4.28 $X2=0 $Y2=0
cc_1046 N_S[1]_c_1020_n N_VGND_c_6269_n 0.00173127f $X=1.065 $Y=4.705 $X2=0
+ $Y2=0
cc_1047 N_S[1]_c_1021_n N_VGND_c_6269_n 0.00525833f $X=1.525 $Y=4.63 $X2=0 $Y2=0
cc_1048 N_S[1]_c_1022_n N_VGND_c_6269_n 0.00862298f $X=1.6 $Y=5.185 $X2=0 $Y2=0
cc_1049 N_S[1]_c_1030_n N_VGND_c_6271_n 0.0028166f $X=3.545 $Y=5.26 $X2=0 $Y2=0
cc_1050 N_S[1]_c_1031_n N_VGND_c_6271_n 5.5039e-19 $X=3.62 $Y=5.185 $X2=0 $Y2=0
cc_1051 N_S[1]_c_1017_n N_VGND_c_6310_n 0.00585385f $X=0.645 $Y=4.705 $X2=0
+ $Y2=0
cc_1052 N_S[1]_c_1018_n N_VGND_c_6310_n 2.16067e-19 $X=0.99 $Y=4.63 $X2=0 $Y2=0
cc_1053 N_S[1]_c_1020_n N_VGND_c_6310_n 0.00542362f $X=1.065 $Y=4.705 $X2=0
+ $Y2=0
cc_1054 N_S[1]_c_1024_n N_VGND_c_6314_n 0.0559651f $X=1.675 $Y=5.26 $X2=0 $Y2=0
cc_1055 N_S[1]_c_1017_n N_VGND_c_6371_n 0.0117149f $X=0.645 $Y=4.705 $X2=0 $Y2=0
cc_1056 N_S[1]_c_1020_n N_VGND_c_6371_n 0.00990284f $X=1.065 $Y=4.705 $X2=0
+ $Y2=0
cc_1057 N_S[1]_c_1023_n N_VGND_c_6371_n 0.0244174f $X=2.285 $Y=5.26 $X2=0 $Y2=0
cc_1058 N_S[1]_c_1024_n N_VGND_c_6371_n 0.0101627f $X=1.675 $Y=5.26 $X2=0 $Y2=0
cc_1059 N_S[1]_c_1026_n N_VGND_c_6371_n 0.00642387f $X=2.705 $Y=5.26 $X2=0 $Y2=0
cc_1060 N_S[1]_c_1028_n N_VGND_c_6371_n 0.0064237f $X=3.125 $Y=5.26 $X2=0 $Y2=0
cc_1061 N_S[1]_c_1030_n N_VGND_c_6371_n 0.0123437f $X=3.545 $Y=5.26 $X2=0 $Y2=0
cc_1062 N_S[1]_c_1033_n N_VGND_c_6371_n 0.00366655f $X=2.36 $Y=5.26 $X2=0 $Y2=0
cc_1063 N_S[1]_c_1034_n N_VGND_c_6371_n 0.00366655f $X=2.78 $Y=5.26 $X2=0 $Y2=0
cc_1064 N_S[1]_c_1035_n N_VGND_c_6371_n 0.00366655f $X=3.2 $Y=5.26 $X2=0 $Y2=0
cc_1065 N_S[1]_c_1021_n N_A_405_918#_c_7010_n 0.00529837f $X=1.525 $Y=4.63 $X2=0
+ $Y2=0
cc_1066 N_S[1]_c_1025_n N_A_405_918#_c_7011_n 0.0112916f $X=2.36 $Y=5.185 $X2=0
+ $Y2=0
cc_1067 N_S[1]_c_1026_n N_A_405_918#_c_7011_n 0.00211351f $X=2.705 $Y=5.26 $X2=0
+ $Y2=0
cc_1068 N_S[1]_c_1027_n N_A_405_918#_c_7011_n 0.0106844f $X=2.78 $Y=5.185 $X2=0
+ $Y2=0
cc_1069 N_S[1]_c_1022_n N_A_405_918#_c_7012_n 0.00189496f $X=1.6 $Y=5.185 $X2=0
+ $Y2=0
cc_1070 N_S[1]_c_1023_n N_A_405_918#_c_7012_n 0.00685838f $X=2.285 $Y=5.26 $X2=0
+ $Y2=0
cc_1071 N_S[1]_c_1029_n N_A_405_918#_c_7013_n 0.0106826f $X=3.2 $Y=5.185 $X2=0
+ $Y2=0
cc_1072 N_S[1]_c_1030_n N_A_405_918#_c_7013_n 0.00211351f $X=3.545 $Y=5.26 $X2=0
+ $Y2=0
cc_1073 N_S[1]_c_1031_n N_A_405_918#_c_7013_n 0.0139014f $X=3.62 $Y=5.185 $X2=0
+ $Y2=0
cc_1074 N_S[1]_c_1031_n N_A_405_918#_c_7016_n 0.00206084f $X=3.62 $Y=5.185 $X2=0
+ $Y2=0
cc_1075 N_S[1]_c_1028_n N_A_405_918#_c_7029_n 0.0034777f $X=3.125 $Y=5.26 $X2=0
+ $Y2=0
cc_1076 N_A_142_325#_c_1141_n N_A_142_599#_c_1253_n 0.0129371f $X=2.135 $Y=1.475
+ $X2=0 $Y2=0
cc_1077 N_A_142_325#_c_1144_n N_A_142_599#_c_1256_n 0.0129371f $X=2.605 $Y=1.475
+ $X2=0 $Y2=0
cc_1078 N_A_142_325#_c_1146_n N_A_142_599#_c_1258_n 0.0129371f $X=3.075 $Y=1.475
+ $X2=0 $Y2=0
cc_1079 N_A_142_325#_c_1148_n N_A_142_599#_c_1260_n 0.0129371f $X=3.545 $Y=1.475
+ $X2=0 $Y2=0
cc_1080 N_A_142_325#_c_1151_n N_VPWR_c_3586_n 0.03379f $X=0.855 $Y=1.77 $X2=0
+ $Y2=0
cc_1081 N_A_142_325#_c_1141_n N_VPWR_c_3588_n 0.00377407f $X=2.135 $Y=1.475
+ $X2=0 $Y2=0
cc_1082 N_A_142_325#_c_1151_n N_VPWR_c_3588_n 0.0302744f $X=0.855 $Y=1.77 $X2=0
+ $Y2=0
cc_1083 N_A_142_325#_c_1137_n N_VPWR_c_3588_n 0.0208071f $X=1.905 $Y=1.23 $X2=0
+ $Y2=0
cc_1084 N_A_142_325#_c_1140_n N_VPWR_c_3588_n 6.4101e-19 $X=1.815 $Y=1.23 $X2=0
+ $Y2=0
cc_1085 N_A_142_325#_c_1148_n N_VPWR_c_3590_n 0.00324472f $X=3.545 $Y=1.475
+ $X2=0 $Y2=0
cc_1086 N_A_142_325#_c_1151_n N_VPWR_c_3626_n 0.0233824f $X=0.855 $Y=1.77 $X2=0
+ $Y2=0
cc_1087 N_A_142_325#_c_1141_n N_VPWR_c_3661_n 0.00473731f $X=2.135 $Y=1.475
+ $X2=0 $Y2=0
cc_1088 N_A_142_325#_c_1144_n N_VPWR_c_3661_n 0.00362156f $X=2.605 $Y=1.475
+ $X2=0 $Y2=0
cc_1089 N_A_142_325#_c_1146_n N_VPWR_c_3661_n 0.00362156f $X=3.075 $Y=1.475
+ $X2=0 $Y2=0
cc_1090 N_A_142_325#_c_1148_n N_VPWR_c_3661_n 0.00473731f $X=3.545 $Y=1.475
+ $X2=0 $Y2=0
cc_1091 N_A_142_325#_c_1151_n N_VPWR_c_3661_n 0.0124581f $X=0.855 $Y=1.77 $X2=0
+ $Y2=0
cc_1092 N_A_142_325#_c_1148_n N_A_355_311#_c_4335_n 0.00151141f $X=3.545
+ $Y=1.475 $X2=0 $Y2=0
cc_1093 N_A_142_325#_c_1141_n N_A_355_311#_c_4343_n 0.00799829f $X=2.135
+ $Y=1.475 $X2=0 $Y2=0
cc_1094 N_A_142_325#_c_1144_n N_A_355_311#_c_4343_n 0.00307958f $X=2.605
+ $Y=1.475 $X2=0 $Y2=0
cc_1095 N_A_142_325#_c_1146_n N_A_355_311#_c_4345_n 0.00307958f $X=3.075
+ $Y=1.475 $X2=0 $Y2=0
cc_1096 N_A_142_325#_c_1148_n N_A_355_311#_c_4345_n 0.00307958f $X=3.545
+ $Y=1.475 $X2=0 $Y2=0
cc_1097 N_A_142_325#_c_1141_n N_A_355_311#_c_4337_n 0.00483827f $X=2.135
+ $Y=1.475 $X2=0 $Y2=0
cc_1098 N_A_142_325#_c_1134_n N_A_355_311#_c_4337_n 0.00561627f $X=2.225 $Y=1.4
+ $X2=0 $Y2=0
cc_1099 N_A_142_325#_c_1137_n N_A_355_311#_c_4337_n 0.0229374f $X=1.905 $Y=1.23
+ $X2=0 $Y2=0
cc_1100 N_A_142_325#_c_1140_n N_A_355_311#_c_4337_n 5.74251e-19 $X=1.815 $Y=1.23
+ $X2=0 $Y2=0
cc_1101 N_A_142_325#_c_1144_n N_A_355_311#_c_4338_n 0.00210632f $X=2.605
+ $Y=1.475 $X2=0 $Y2=0
cc_1102 N_A_142_325#_c_1145_n N_A_355_311#_c_4338_n 0.00251792f $X=2.985 $Y=1.4
+ $X2=0 $Y2=0
cc_1103 N_A_142_325#_c_1146_n N_A_355_311#_c_4338_n 0.00210632f $X=3.075
+ $Y=1.475 $X2=0 $Y2=0
cc_1104 N_A_142_325#_c_1148_n N_A_355_311#_c_4339_n 0.00554566f $X=3.545
+ $Y=1.475 $X2=0 $Y2=0
cc_1105 N_A_142_325#_c_1145_n N_Z_c_4590_n 0.00762343f $X=2.985 $Y=1.4 $X2=0
+ $Y2=0
cc_1106 N_A_142_325#_c_1150_n N_Z_c_4590_n 0.00704092f $X=3.075 $Y=1.4 $X2=0
+ $Y2=0
cc_1107 N_A_142_325#_c_1142_n N_Z_c_4608_n 0.00597584f $X=2.515 $Y=1.4 $X2=0
+ $Y2=0
cc_1108 N_A_142_325#_c_1134_n N_Z_c_4608_n 0.00747617f $X=2.225 $Y=1.4 $X2=0
+ $Y2=0
cc_1109 N_A_142_325#_c_1145_n N_Z_c_4608_n 0.00145542f $X=2.985 $Y=1.4 $X2=0
+ $Y2=0
cc_1110 N_A_142_325#_c_1149_n N_Z_c_4608_n 0.00909323f $X=2.605 $Y=1.4 $X2=0
+ $Y2=0
cc_1111 N_A_142_325#_c_1137_n N_Z_c_4608_n 0.0266078f $X=1.905 $Y=1.23 $X2=0
+ $Y2=0
cc_1112 N_A_142_325#_c_1147_n N_Z_c_4610_n 0.00918337f $X=3.455 $Y=1.4 $X2=0
+ $Y2=0
cc_1113 N_A_142_325#_c_1150_n N_Z_c_4610_n 2.98555e-19 $X=3.075 $Y=1.4 $X2=0
+ $Y2=0
cc_1114 N_A_142_325#_c_1147_n N_Z_c_4612_n 0.00248496f $X=3.455 $Y=1.4 $X2=0
+ $Y2=0
cc_1115 N_A_142_325#_c_1148_n N_Z_c_4644_n 0.00834829f $X=3.545 $Y=1.475 $X2=0
+ $Y2=0
cc_1116 N_A_142_325#_c_1144_n N_Z_c_4693_n 0.00372248f $X=2.605 $Y=1.475 $X2=0
+ $Y2=0
cc_1117 N_A_142_325#_c_1146_n N_Z_c_4693_n 0.00372458f $X=3.075 $Y=1.475 $X2=0
+ $Y2=0
cc_1118 N_A_142_325#_c_1141_n N_Z_c_4650_n 0.0226667f $X=2.135 $Y=1.475 $X2=0
+ $Y2=0
cc_1119 N_A_142_325#_c_1142_n N_Z_c_4650_n 0.00560592f $X=2.515 $Y=1.4 $X2=0
+ $Y2=0
cc_1120 N_A_142_325#_c_1134_n N_Z_c_4650_n 0.00425035f $X=2.225 $Y=1.4 $X2=0
+ $Y2=0
cc_1121 N_A_142_325#_c_1144_n N_Z_c_4650_n 0.0181262f $X=2.605 $Y=1.475 $X2=0
+ $Y2=0
cc_1122 N_A_142_325#_c_1146_n N_Z_c_4650_n 9.74366e-19 $X=3.075 $Y=1.475 $X2=0
+ $Y2=0
cc_1123 N_A_142_325#_c_1149_n N_Z_c_4650_n 0.00181273f $X=2.605 $Y=1.4 $X2=0
+ $Y2=0
cc_1124 N_A_142_325#_c_1137_n N_Z_c_4650_n 0.00240108f $X=1.905 $Y=1.23 $X2=0
+ $Y2=0
cc_1125 N_A_142_325#_c_1144_n N_Z_c_4651_n 9.74366e-19 $X=2.605 $Y=1.475 $X2=0
+ $Y2=0
cc_1126 N_A_142_325#_c_1146_n N_Z_c_4651_n 0.0181262f $X=3.075 $Y=1.475 $X2=0
+ $Y2=0
cc_1127 N_A_142_325#_c_1147_n N_Z_c_4651_n 0.0103509f $X=3.455 $Y=1.4 $X2=0
+ $Y2=0
cc_1128 N_A_142_325#_c_1148_n N_Z_c_4651_n 0.0199111f $X=3.545 $Y=1.475 $X2=0
+ $Y2=0
cc_1129 N_A_142_325#_c_1150_n N_Z_c_4651_n 0.00415268f $X=3.075 $Y=1.4 $X2=0
+ $Y2=0
cc_1130 N_A_142_325#_c_1137_n N_VGND_c_6268_n 0.0123065f $X=1.905 $Y=1.23 $X2=0
+ $Y2=0
cc_1131 N_A_142_325#_c_1140_n N_VGND_c_6268_n 2.04129e-19 $X=1.815 $Y=1.23 $X2=0
+ $Y2=0
cc_1132 N_A_142_325#_c_1135_n N_VGND_c_6308_n 0.0129994f $X=0.855 $Y=0.445 $X2=0
+ $Y2=0
cc_1133 N_A_142_325#_M1043_s N_VGND_c_6370_n 0.00394793f $X=0.72 $Y=0.235 $X2=0
+ $Y2=0
cc_1134 N_A_142_325#_c_1135_n N_VGND_c_6370_n 0.00927134f $X=0.855 $Y=0.445
+ $X2=0 $Y2=0
cc_1135 N_A_142_325#_c_1134_n N_A_405_66#_c_6926_n 0.00600378f $X=2.225 $Y=1.4
+ $X2=0 $Y2=0
cc_1136 N_A_142_325#_c_1137_n N_A_405_66#_c_6926_n 0.0028695f $X=1.905 $Y=1.23
+ $X2=0 $Y2=0
cc_1137 N_A_142_325#_c_1145_n N_A_405_66#_c_6948_n 7.0477e-19 $X=2.985 $Y=1.4
+ $X2=0 $Y2=0
cc_1138 N_A_142_599#_c_1263_n N_VPWR_c_3587_n 0.03379f $X=0.855 $Y=3.14 $X2=0
+ $Y2=0
cc_1139 N_A_142_599#_c_1253_n N_VPWR_c_3589_n 0.00377407f $X=2.135 $Y=3.965
+ $X2=0 $Y2=0
cc_1140 N_A_142_599#_c_1263_n N_VPWR_c_3589_n 0.0302744f $X=0.855 $Y=3.14 $X2=0
+ $Y2=0
cc_1141 N_A_142_599#_c_1249_n N_VPWR_c_3589_n 0.0208071f $X=1.905 $Y=4.21 $X2=0
+ $Y2=0
cc_1142 N_A_142_599#_c_1252_n N_VPWR_c_3589_n 6.4101e-19 $X=1.815 $Y=4.21 $X2=0
+ $Y2=0
cc_1143 N_A_142_599#_c_1260_n N_VPWR_c_3591_n 0.00324472f $X=3.545 $Y=3.965
+ $X2=0 $Y2=0
cc_1144 N_A_142_599#_c_1263_n N_VPWR_c_3626_n 0.0233824f $X=0.855 $Y=3.14 $X2=0
+ $Y2=0
cc_1145 N_A_142_599#_c_1253_n N_VPWR_c_3661_n 0.00473731f $X=2.135 $Y=3.965
+ $X2=0 $Y2=0
cc_1146 N_A_142_599#_c_1256_n N_VPWR_c_3661_n 0.00362156f $X=2.605 $Y=3.965
+ $X2=0 $Y2=0
cc_1147 N_A_142_599#_c_1258_n N_VPWR_c_3661_n 0.00362156f $X=3.075 $Y=3.965
+ $X2=0 $Y2=0
cc_1148 N_A_142_599#_c_1260_n N_VPWR_c_3661_n 0.00473731f $X=3.545 $Y=3.965
+ $X2=0 $Y2=0
cc_1149 N_A_142_599#_c_1263_n N_VPWR_c_3661_n 0.0124581f $X=0.855 $Y=3.14 $X2=0
+ $Y2=0
cc_1150 N_A_142_599#_c_1260_n N_A_355_613#_c_4462_n 0.00151141f $X=3.545
+ $Y=3.965 $X2=0 $Y2=0
cc_1151 N_A_142_599#_c_1253_n N_A_355_613#_c_4470_n 0.00799829f $X=2.135
+ $Y=3.965 $X2=0 $Y2=0
cc_1152 N_A_142_599#_c_1256_n N_A_355_613#_c_4470_n 0.00307958f $X=2.605
+ $Y=3.965 $X2=0 $Y2=0
cc_1153 N_A_142_599#_c_1258_n N_A_355_613#_c_4472_n 0.00307958f $X=3.075
+ $Y=3.965 $X2=0 $Y2=0
cc_1154 N_A_142_599#_c_1260_n N_A_355_613#_c_4472_n 0.00307958f $X=3.545
+ $Y=3.965 $X2=0 $Y2=0
cc_1155 N_A_142_599#_c_1253_n N_A_355_613#_c_4464_n 0.00483827f $X=2.135
+ $Y=3.965 $X2=0 $Y2=0
cc_1156 N_A_142_599#_c_1246_n N_A_355_613#_c_4464_n 0.00561627f $X=2.225 $Y=4.04
+ $X2=0 $Y2=0
cc_1157 N_A_142_599#_c_1249_n N_A_355_613#_c_4464_n 0.0229374f $X=1.905 $Y=4.21
+ $X2=0 $Y2=0
cc_1158 N_A_142_599#_c_1252_n N_A_355_613#_c_4464_n 5.74251e-19 $X=1.815 $Y=4.21
+ $X2=0 $Y2=0
cc_1159 N_A_142_599#_c_1256_n N_A_355_613#_c_4465_n 0.00210632f $X=2.605
+ $Y=3.965 $X2=0 $Y2=0
cc_1160 N_A_142_599#_c_1257_n N_A_355_613#_c_4465_n 0.00251792f $X=2.985 $Y=4.04
+ $X2=0 $Y2=0
cc_1161 N_A_142_599#_c_1258_n N_A_355_613#_c_4465_n 0.00210632f $X=3.075
+ $Y=3.965 $X2=0 $Y2=0
cc_1162 N_A_142_599#_c_1260_n N_A_355_613#_c_4466_n 0.00554566f $X=3.545
+ $Y=3.965 $X2=0 $Y2=0
cc_1163 N_A_142_599#_c_1257_n N_Z_c_4591_n 0.00762343f $X=2.985 $Y=4.04 $X2=0
+ $Y2=0
cc_1164 N_A_142_599#_c_1262_n N_Z_c_4591_n 0.00704092f $X=3.075 $Y=4.04 $X2=0
+ $Y2=0
cc_1165 N_A_142_599#_c_1254_n N_Z_c_4609_n 0.00597584f $X=2.515 $Y=4.04 $X2=0
+ $Y2=0
cc_1166 N_A_142_599#_c_1246_n N_Z_c_4609_n 0.00747617f $X=2.225 $Y=4.04 $X2=0
+ $Y2=0
cc_1167 N_A_142_599#_c_1257_n N_Z_c_4609_n 0.00145542f $X=2.985 $Y=4.04 $X2=0
+ $Y2=0
cc_1168 N_A_142_599#_c_1261_n N_Z_c_4609_n 0.00909323f $X=2.605 $Y=4.04 $X2=0
+ $Y2=0
cc_1169 N_A_142_599#_c_1249_n N_Z_c_4609_n 0.0266078f $X=1.905 $Y=4.21 $X2=0
+ $Y2=0
cc_1170 N_A_142_599#_c_1259_n N_Z_c_4611_n 0.00918337f $X=3.455 $Y=4.04 $X2=0
+ $Y2=0
cc_1171 N_A_142_599#_c_1262_n N_Z_c_4611_n 2.98555e-19 $X=3.075 $Y=4.04 $X2=0
+ $Y2=0
cc_1172 N_A_142_599#_c_1259_n N_Z_c_4613_n 0.00248496f $X=3.455 $Y=4.04 $X2=0
+ $Y2=0
cc_1173 N_A_142_599#_c_1260_n N_Z_c_4645_n 0.00834829f $X=3.545 $Y=3.965 $X2=0
+ $Y2=0
cc_1174 N_A_142_599#_c_1256_n N_Z_c_4718_n 0.00372248f $X=2.605 $Y=3.965 $X2=0
+ $Y2=0
cc_1175 N_A_142_599#_c_1258_n N_Z_c_4718_n 0.00372458f $X=3.075 $Y=3.965 $X2=0
+ $Y2=0
cc_1176 N_A_142_599#_c_1253_n N_Z_c_4650_n 0.0226667f $X=2.135 $Y=3.965 $X2=0
+ $Y2=0
cc_1177 N_A_142_599#_c_1254_n N_Z_c_4650_n 0.00560592f $X=2.515 $Y=4.04 $X2=0
+ $Y2=0
cc_1178 N_A_142_599#_c_1246_n N_Z_c_4650_n 0.00425035f $X=2.225 $Y=4.04 $X2=0
+ $Y2=0
cc_1179 N_A_142_599#_c_1256_n N_Z_c_4650_n 0.0181262f $X=2.605 $Y=3.965 $X2=0
+ $Y2=0
cc_1180 N_A_142_599#_c_1258_n N_Z_c_4650_n 9.74366e-19 $X=3.075 $Y=3.965 $X2=0
+ $Y2=0
cc_1181 N_A_142_599#_c_1261_n N_Z_c_4650_n 0.00181273f $X=2.605 $Y=4.04 $X2=0
+ $Y2=0
cc_1182 N_A_142_599#_c_1249_n N_Z_c_4650_n 0.00240108f $X=1.905 $Y=4.21 $X2=0
+ $Y2=0
cc_1183 N_A_142_599#_c_1256_n N_Z_c_4651_n 9.74366e-19 $X=2.605 $Y=3.965 $X2=0
+ $Y2=0
cc_1184 N_A_142_599#_c_1258_n N_Z_c_4651_n 0.0181262f $X=3.075 $Y=3.965 $X2=0
+ $Y2=0
cc_1185 N_A_142_599#_c_1259_n N_Z_c_4651_n 0.0103509f $X=3.455 $Y=4.04 $X2=0
+ $Y2=0
cc_1186 N_A_142_599#_c_1260_n N_Z_c_4651_n 0.0199111f $X=3.545 $Y=3.965 $X2=0
+ $Y2=0
cc_1187 N_A_142_599#_c_1262_n N_Z_c_4651_n 0.00415268f $X=3.075 $Y=4.04 $X2=0
+ $Y2=0
cc_1188 N_A_142_599#_c_1249_n N_VGND_c_6269_n 0.0123065f $X=1.905 $Y=4.21 $X2=0
+ $Y2=0
cc_1189 N_A_142_599#_c_1252_n N_VGND_c_6269_n 2.04129e-19 $X=1.815 $Y=4.21 $X2=0
+ $Y2=0
cc_1190 N_A_142_599#_c_1248_n N_VGND_c_6310_n 0.0129994f $X=0.855 $Y=4.995 $X2=0
+ $Y2=0
cc_1191 N_A_142_599#_M1084_d N_VGND_c_6371_n 0.00394793f $X=0.72 $Y=4.785 $X2=0
+ $Y2=0
cc_1192 N_A_142_599#_c_1248_n N_VGND_c_6371_n 0.00927134f $X=0.855 $Y=4.995
+ $X2=0 $Y2=0
cc_1193 N_A_142_599#_c_1246_n N_A_405_918#_c_7010_n 0.00600378f $X=2.225 $Y=4.04
+ $X2=0 $Y2=0
cc_1194 N_A_142_599#_c_1249_n N_A_405_918#_c_7010_n 0.0028695f $X=1.905 $Y=4.21
+ $X2=0 $Y2=0
cc_1195 N_A_142_599#_c_1257_n N_A_405_918#_c_7032_n 7.0477e-19 $X=2.985 $Y=4.04
+ $X2=0 $Y2=0
cc_1196 N_D[0]_M1012_g N_D[1]_M1017_g 0.0130744f $X=4.535 $Y=1.985 $X2=0 $Y2=0
cc_1197 N_D[0]_M1049_g N_D[1]_M1055_g 0.0130744f $X=5.005 $Y=1.985 $X2=0 $Y2=0
cc_1198 N_D[0]_M1086_g N_D[1]_M1093_g 0.0130744f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1199 N_D[0]_M1137_g N_D[1]_M1141_g 0.0130744f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1200 N_D[0]_M1137_g N_D[2]_M1071_g 0.0129367f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1201 N_D[0]_M1156_g N_D[2]_M1013_g 0.0210205f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_1202 N_D[0]_c_1374_n N_D[2]_c_1569_n 2.99666e-19 $X=5.84 $Y=1.16 $X2=0 $Y2=0
cc_1203 N_D[0]_c_1375_n N_D[2]_c_1569_n 0.0105491f $X=5.945 $Y=1.16 $X2=0 $Y2=0
cc_1204 N_D[0]_c_1374_n N_D[2]_c_1570_n 0.0135469f $X=5.84 $Y=1.16 $X2=0 $Y2=0
cc_1205 N_D[0]_c_1375_n N_D[2]_c_1570_n 2.99666e-19 $X=5.945 $Y=1.16 $X2=0 $Y2=0
cc_1206 N_D[0]_M1012_g N_VPWR_c_3590_n 0.00389633f $X=4.535 $Y=1.985 $X2=0 $Y2=0
cc_1207 N_D[0]_M1049_g N_VPWR_c_3592_n 0.00208662f $X=5.005 $Y=1.985 $X2=0 $Y2=0
cc_1208 N_D[0]_M1086_g N_VPWR_c_3592_n 0.00208662f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1209 N_D[0]_M1137_g N_VPWR_c_3594_n 0.00207065f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1210 N_D[0]_M1012_g N_VPWR_c_3641_n 0.0035837f $X=4.535 $Y=1.985 $X2=0 $Y2=0
cc_1211 N_D[0]_M1049_g N_VPWR_c_3641_n 0.0035837f $X=5.005 $Y=1.985 $X2=0 $Y2=0
cc_1212 N_D[0]_M1086_g N_VPWR_c_3642_n 0.0035837f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1213 N_D[0]_M1137_g N_VPWR_c_3642_n 0.0035837f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1214 N_D[0]_M1012_g N_VPWR_c_3661_n 0.00573859f $X=4.535 $Y=1.985 $X2=0 $Y2=0
cc_1215 N_D[0]_M1049_g N_VPWR_c_3661_n 0.00445624f $X=5.005 $Y=1.985 $X2=0 $Y2=0
cc_1216 N_D[0]_M1086_g N_VPWR_c_3661_n 0.00445624f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1217 N_D[0]_M1137_g N_VPWR_c_3661_n 0.00579371f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1218 N_D[0]_M1012_g N_A_355_311#_c_4334_n 0.013247f $X=4.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1219 N_D[0]_M1049_g N_A_355_311#_c_4356_n 0.00916655f $X=5.005 $Y=1.985 $X2=0
+ $Y2=0
cc_1220 N_D[0]_M1086_g N_A_355_311#_c_4356_n 0.00916655f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_1221 N_D[0]_c_1372_n N_A_355_311#_c_4356_n 7.15862e-19 $X=5.385 $Y=1.16 $X2=0
+ $Y2=0
cc_1222 N_D[0]_c_1374_n N_A_355_311#_c_4356_n 0.0387168f $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_1223 N_D[0]_M1012_g N_A_355_311#_c_4360_n 8.61029e-19 $X=4.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1224 N_D[0]_M1049_g N_A_355_311#_c_4360_n 5.79575e-19 $X=5.005 $Y=1.985 $X2=0
+ $Y2=0
cc_1225 N_D[0]_c_1373_n N_A_355_311#_c_4360_n 8.03631e-19 $X=5.095 $Y=1.16 $X2=0
+ $Y2=0
cc_1226 N_D[0]_c_1374_n N_A_355_311#_c_4360_n 0.0191156f $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_1227 N_D[0]_M1086_g N_A_355_311#_c_4364_n 5.79575e-19 $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_1228 N_D[0]_M1137_g N_A_355_311#_c_4364_n 0.002088f $X=5.945 $Y=1.985 $X2=0
+ $Y2=0
cc_1229 N_D[0]_c_1374_n N_A_355_311#_c_4364_n 0.0217153f $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_1230 N_D[0]_c_1375_n N_A_355_311#_c_4364_n 8.03631e-19 $X=5.945 $Y=1.16 $X2=0
+ $Y2=0
cc_1231 N_D[0]_M1012_g N_A_355_311#_c_4336_n 0.00232998f $X=4.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1232 N_D[0]_M1049_g N_A_355_311#_c_4369_n 0.00232998f $X=5.005 $Y=1.985 $X2=0
+ $Y2=0
cc_1233 N_D[0]_M1086_g N_A_355_311#_c_4369_n 0.00232998f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_1234 N_D[0]_M1012_g N_A_355_311#_c_4371_n 0.00977623f $X=4.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1235 N_D[0]_M1049_g N_A_355_311#_c_4371_n 0.00911325f $X=5.005 $Y=1.985 $X2=0
+ $Y2=0
cc_1236 N_D[0]_M1086_g N_A_355_311#_c_4371_n 7.05028e-19 $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_1237 N_D[0]_M1049_g N_A_355_311#_c_4374_n 7.05028e-19 $X=5.005 $Y=1.985 $X2=0
+ $Y2=0
cc_1238 N_D[0]_M1086_g N_A_355_311#_c_4374_n 0.00911325f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_1239 N_D[0]_M1137_g N_A_355_311#_c_4374_n 0.00819194f $X=5.945 $Y=1.985 $X2=0
+ $Y2=0
cc_1240 N_D[0]_M1012_g N_A_355_311#_c_4339_n 0.00333758f $X=4.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1241 N_D[0]_M1012_g N_Z_c_4644_n 0.00311896f $X=4.535 $Y=1.985 $X2=0 $Y2=0
cc_1242 N_D[0]_M1049_g N_Z_c_4644_n 0.00306964f $X=5.005 $Y=1.985 $X2=0 $Y2=0
cc_1243 N_D[0]_M1086_g N_Z_c_4644_n 0.00306964f $X=5.475 $Y=1.985 $X2=0 $Y2=0
cc_1244 N_D[0]_M1137_g N_Z_c_4644_n 0.00470782f $X=5.945 $Y=1.985 $X2=0 $Y2=0
cc_1245 N_D[0]_c_1374_n N_Z_c_4644_n 0.00846955f $X=5.84 $Y=1.16 $X2=0 $Y2=0
cc_1246 N_D[0]_M1065_g N_VGND_c_6270_n 0.00321269f $X=4.56 $Y=0.56 $X2=0 $Y2=0
cc_1247 N_D[0]_M1097_g N_VGND_c_6270_n 2.6376e-19 $X=4.98 $Y=0.56 $X2=0 $Y2=0
cc_1248 N_D[0]_M1097_g N_VGND_c_6272_n 0.0019152f $X=4.98 $Y=0.56 $X2=0 $Y2=0
cc_1249 N_D[0]_M1151_g N_VGND_c_6272_n 0.00166854f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_1250 N_D[0]_M1156_g N_VGND_c_6272_n 2.64031e-19 $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_1251 N_D[0]_M1156_g N_VGND_c_6274_n 0.0058918f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_1252 N_D[0]_M1065_g N_VGND_c_6340_n 0.00422241f $X=4.56 $Y=0.56 $X2=0 $Y2=0
cc_1253 N_D[0]_M1097_g N_VGND_c_6340_n 0.00430643f $X=4.98 $Y=0.56 $X2=0 $Y2=0
cc_1254 N_D[0]_M1151_g N_VGND_c_6342_n 0.00422241f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_1255 N_D[0]_M1156_g N_VGND_c_6342_n 0.00551064f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_1256 N_D[0]_M1065_g N_VGND_c_6370_n 0.00702263f $X=4.56 $Y=0.56 $X2=0 $Y2=0
cc_1257 N_D[0]_M1097_g N_VGND_c_6370_n 0.00624811f $X=4.98 $Y=0.56 $X2=0 $Y2=0
cc_1258 N_D[0]_M1151_g N_VGND_c_6370_n 0.00593887f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_1259 N_D[0]_M1156_g N_VGND_c_6370_n 0.0101978f $X=5.92 $Y=0.56 $X2=0 $Y2=0
cc_1260 N_D[0]_M1065_g N_A_405_66#_c_6930_n 0.00261078f $X=4.56 $Y=0.56 $X2=0
+ $Y2=0
cc_1261 N_D[0]_M1065_g N_A_405_66#_c_6931_n 0.0121912f $X=4.56 $Y=0.56 $X2=0
+ $Y2=0
cc_1262 N_D[0]_M1065_g N_A_405_66#_c_6951_n 0.00699463f $X=4.56 $Y=0.56 $X2=0
+ $Y2=0
cc_1263 N_D[0]_M1097_g N_A_405_66#_c_6951_n 0.00661764f $X=4.98 $Y=0.56 $X2=0
+ $Y2=0
cc_1264 N_D[0]_M1151_g N_A_405_66#_c_6951_n 5.22365e-19 $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_1265 N_D[0]_M1097_g N_A_405_66#_c_6933_n 0.00900364f $X=4.98 $Y=0.56 $X2=0
+ $Y2=0
cc_1266 N_D[0]_M1151_g N_A_405_66#_c_6933_n 0.00986515f $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_1267 N_D[0]_M1156_g N_A_405_66#_c_6933_n 0.00222549f $X=5.92 $Y=0.56 $X2=0
+ $Y2=0
cc_1268 N_D[0]_c_1372_n N_A_405_66#_c_6933_n 0.00463549f $X=5.385 $Y=1.16 $X2=0
+ $Y2=0
cc_1269 N_D[0]_c_1374_n N_A_405_66#_c_6933_n 0.0608884f $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_1270 N_D[0]_c_1375_n N_A_405_66#_c_6933_n 0.00208088f $X=5.945 $Y=1.16 $X2=0
+ $Y2=0
cc_1271 N_D[0]_M1097_g N_A_405_66#_c_6960_n 5.22365e-19 $X=4.98 $Y=0.56 $X2=0
+ $Y2=0
cc_1272 N_D[0]_M1151_g N_A_405_66#_c_6960_n 0.00661134f $X=5.5 $Y=0.56 $X2=0
+ $Y2=0
cc_1273 N_D[0]_M1156_g N_A_405_66#_c_6960_n 0.00514241f $X=5.92 $Y=0.56 $X2=0
+ $Y2=0
cc_1274 N_D[0]_M1065_g N_A_405_66#_c_6934_n 0.00128201f $X=4.56 $Y=0.56 $X2=0
+ $Y2=0
cc_1275 N_D[0]_M1097_g N_A_405_66#_c_6934_n 8.68782e-19 $X=4.98 $Y=0.56 $X2=0
+ $Y2=0
cc_1276 N_D[0]_c_1373_n N_A_405_66#_c_6934_n 0.00208088f $X=5.095 $Y=1.16 $X2=0
+ $Y2=0
cc_1277 N_D[0]_c_1374_n N_A_405_66#_c_6934_n 0.018367f $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_1278 N_D[1]_M1141_g N_D[3]_M1000_g 0.0129367f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1279 N_D[1]_M1157_g N_D[3]_M1015_g 0.0210205f $X=5.92 $Y=4.88 $X2=0 $Y2=0
cc_1280 N_D[1]_c_1473_n N_D[3]_c_1670_n 2.99666e-19 $X=5.84 $Y=4.28 $X2=0 $Y2=0
cc_1281 N_D[1]_c_1474_n N_D[3]_c_1670_n 0.0105491f $X=5.945 $Y=4.28 $X2=0 $Y2=0
cc_1282 N_D[1]_c_1473_n N_D[3]_c_1671_n 0.0135469f $X=5.84 $Y=4.28 $X2=0 $Y2=0
cc_1283 N_D[1]_c_1474_n N_D[3]_c_1671_n 2.99666e-19 $X=5.945 $Y=4.28 $X2=0 $Y2=0
cc_1284 N_D[1]_M1017_g N_VPWR_c_3591_n 0.00389633f $X=4.535 $Y=3.455 $X2=0 $Y2=0
cc_1285 N_D[1]_M1055_g N_VPWR_c_3593_n 0.00208662f $X=5.005 $Y=3.455 $X2=0 $Y2=0
cc_1286 N_D[1]_M1093_g N_VPWR_c_3593_n 0.00208662f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1287 N_D[1]_M1141_g N_VPWR_c_3595_n 0.00207065f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1288 N_D[1]_M1017_g N_VPWR_c_3641_n 0.0035837f $X=4.535 $Y=3.455 $X2=0 $Y2=0
cc_1289 N_D[1]_M1055_g N_VPWR_c_3641_n 0.0035837f $X=5.005 $Y=3.455 $X2=0 $Y2=0
cc_1290 N_D[1]_M1093_g N_VPWR_c_3642_n 0.0035837f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1291 N_D[1]_M1141_g N_VPWR_c_3642_n 0.0035837f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1292 N_D[1]_M1017_g N_VPWR_c_3661_n 0.00573859f $X=4.535 $Y=3.455 $X2=0 $Y2=0
cc_1293 N_D[1]_M1055_g N_VPWR_c_3661_n 0.00445624f $X=5.005 $Y=3.455 $X2=0 $Y2=0
cc_1294 N_D[1]_M1093_g N_VPWR_c_3661_n 0.00445624f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1295 N_D[1]_M1141_g N_VPWR_c_3661_n 0.00579371f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1296 N_D[1]_M1017_g N_A_355_613#_c_4461_n 0.013247f $X=4.535 $Y=3.455 $X2=0
+ $Y2=0
cc_1297 N_D[1]_M1055_g N_A_355_613#_c_4483_n 0.00916655f $X=5.005 $Y=3.455 $X2=0
+ $Y2=0
cc_1298 N_D[1]_M1093_g N_A_355_613#_c_4483_n 0.00916655f $X=5.475 $Y=3.455 $X2=0
+ $Y2=0
cc_1299 N_D[1]_c_1471_n N_A_355_613#_c_4483_n 7.15862e-19 $X=5.385 $Y=4.28 $X2=0
+ $Y2=0
cc_1300 N_D[1]_c_1473_n N_A_355_613#_c_4483_n 0.0387168f $X=5.84 $Y=4.28 $X2=0
+ $Y2=0
cc_1301 N_D[1]_M1017_g N_A_355_613#_c_4487_n 8.61029e-19 $X=4.535 $Y=3.455 $X2=0
+ $Y2=0
cc_1302 N_D[1]_M1055_g N_A_355_613#_c_4487_n 5.79575e-19 $X=5.005 $Y=3.455 $X2=0
+ $Y2=0
cc_1303 N_D[1]_c_1472_n N_A_355_613#_c_4487_n 8.03631e-19 $X=5.095 $Y=4.28 $X2=0
+ $Y2=0
cc_1304 N_D[1]_c_1473_n N_A_355_613#_c_4487_n 0.0191156f $X=5.84 $Y=4.28 $X2=0
+ $Y2=0
cc_1305 N_D[1]_M1093_g N_A_355_613#_c_4491_n 5.79575e-19 $X=5.475 $Y=3.455 $X2=0
+ $Y2=0
cc_1306 N_D[1]_M1141_g N_A_355_613#_c_4491_n 0.002088f $X=5.945 $Y=3.455 $X2=0
+ $Y2=0
cc_1307 N_D[1]_c_1473_n N_A_355_613#_c_4491_n 0.0217153f $X=5.84 $Y=4.28 $X2=0
+ $Y2=0
cc_1308 N_D[1]_c_1474_n N_A_355_613#_c_4491_n 8.03631e-19 $X=5.945 $Y=4.28 $X2=0
+ $Y2=0
cc_1309 N_D[1]_M1017_g N_A_355_613#_c_4463_n 0.00232998f $X=4.535 $Y=3.455 $X2=0
+ $Y2=0
cc_1310 N_D[1]_M1055_g N_A_355_613#_c_4496_n 0.00232998f $X=5.005 $Y=3.455 $X2=0
+ $Y2=0
cc_1311 N_D[1]_M1093_g N_A_355_613#_c_4496_n 0.00232998f $X=5.475 $Y=3.455 $X2=0
+ $Y2=0
cc_1312 N_D[1]_M1017_g N_A_355_613#_c_4466_n 0.00333758f $X=4.535 $Y=3.455 $X2=0
+ $Y2=0
cc_1313 N_D[1]_M1017_g N_A_355_613#_c_4499_n 0.00977623f $X=4.535 $Y=3.455 $X2=0
+ $Y2=0
cc_1314 N_D[1]_M1055_g N_A_355_613#_c_4499_n 0.00911325f $X=5.005 $Y=3.455 $X2=0
+ $Y2=0
cc_1315 N_D[1]_M1093_g N_A_355_613#_c_4499_n 7.05028e-19 $X=5.475 $Y=3.455 $X2=0
+ $Y2=0
cc_1316 N_D[1]_M1055_g N_A_355_613#_c_4502_n 7.05028e-19 $X=5.005 $Y=3.455 $X2=0
+ $Y2=0
cc_1317 N_D[1]_M1093_g N_A_355_613#_c_4502_n 0.00911325f $X=5.475 $Y=3.455 $X2=0
+ $Y2=0
cc_1318 N_D[1]_M1141_g N_A_355_613#_c_4502_n 0.00819194f $X=5.945 $Y=3.455 $X2=0
+ $Y2=0
cc_1319 N_D[1]_M1017_g N_Z_c_4645_n 0.00311896f $X=4.535 $Y=3.455 $X2=0 $Y2=0
cc_1320 N_D[1]_M1055_g N_Z_c_4645_n 0.00306964f $X=5.005 $Y=3.455 $X2=0 $Y2=0
cc_1321 N_D[1]_M1093_g N_Z_c_4645_n 0.00306964f $X=5.475 $Y=3.455 $X2=0 $Y2=0
cc_1322 N_D[1]_M1141_g N_Z_c_4645_n 0.00470782f $X=5.945 $Y=3.455 $X2=0 $Y2=0
cc_1323 N_D[1]_c_1473_n N_Z_c_4645_n 0.00846955f $X=5.84 $Y=4.28 $X2=0 $Y2=0
cc_1324 N_D[1]_M1030_g N_VGND_c_6271_n 0.00321269f $X=4.56 $Y=4.88 $X2=0 $Y2=0
cc_1325 N_D[1]_M1059_g N_VGND_c_6271_n 2.6376e-19 $X=4.98 $Y=4.88 $X2=0 $Y2=0
cc_1326 N_D[1]_M1059_g N_VGND_c_6273_n 0.0019152f $X=4.98 $Y=4.88 $X2=0 $Y2=0
cc_1327 N_D[1]_M1068_g N_VGND_c_6273_n 0.00166854f $X=5.5 $Y=4.88 $X2=0 $Y2=0
cc_1328 N_D[1]_M1157_g N_VGND_c_6273_n 2.64031e-19 $X=5.92 $Y=4.88 $X2=0 $Y2=0
cc_1329 N_D[1]_M1157_g N_VGND_c_6275_n 0.0058918f $X=5.92 $Y=4.88 $X2=0 $Y2=0
cc_1330 N_D[1]_M1030_g N_VGND_c_6341_n 0.00422241f $X=4.56 $Y=4.88 $X2=0 $Y2=0
cc_1331 N_D[1]_M1059_g N_VGND_c_6341_n 0.00430643f $X=4.98 $Y=4.88 $X2=0 $Y2=0
cc_1332 N_D[1]_M1068_g N_VGND_c_6343_n 0.00422241f $X=5.5 $Y=4.88 $X2=0 $Y2=0
cc_1333 N_D[1]_M1157_g N_VGND_c_6343_n 0.00551064f $X=5.92 $Y=4.88 $X2=0 $Y2=0
cc_1334 N_D[1]_M1030_g N_VGND_c_6371_n 0.00702263f $X=4.56 $Y=4.88 $X2=0 $Y2=0
cc_1335 N_D[1]_M1059_g N_VGND_c_6371_n 0.00624811f $X=4.98 $Y=4.88 $X2=0 $Y2=0
cc_1336 N_D[1]_M1068_g N_VGND_c_6371_n 0.00593887f $X=5.5 $Y=4.88 $X2=0 $Y2=0
cc_1337 N_D[1]_M1157_g N_VGND_c_6371_n 0.0101978f $X=5.92 $Y=4.88 $X2=0 $Y2=0
cc_1338 N_D[1]_M1030_g N_A_405_918#_c_7014_n 0.00261078f $X=4.56 $Y=4.88 $X2=0
+ $Y2=0
cc_1339 N_D[1]_M1030_g N_A_405_918#_c_7015_n 0.0121912f $X=4.56 $Y=4.88 $X2=0
+ $Y2=0
cc_1340 N_D[1]_M1059_g N_A_405_918#_c_7035_n 0.00900364f $X=4.98 $Y=4.88 $X2=0
+ $Y2=0
cc_1341 N_D[1]_M1068_g N_A_405_918#_c_7035_n 0.00899636f $X=5.5 $Y=4.88 $X2=0
+ $Y2=0
cc_1342 N_D[1]_c_1471_n N_A_405_918#_c_7035_n 0.00463549f $X=5.385 $Y=4.28 $X2=0
+ $Y2=0
cc_1343 N_D[1]_c_1473_n N_A_405_918#_c_7035_n 0.0394855f $X=5.84 $Y=4.28 $X2=0
+ $Y2=0
cc_1344 N_D[1]_M1030_g N_A_405_918#_c_7017_n 0.00827664f $X=4.56 $Y=4.88 $X2=0
+ $Y2=0
cc_1345 N_D[1]_M1059_g N_A_405_918#_c_7017_n 0.00748643f $X=4.98 $Y=4.88 $X2=0
+ $Y2=0
cc_1346 N_D[1]_M1068_g N_A_405_918#_c_7017_n 5.22365e-19 $X=5.5 $Y=4.88 $X2=0
+ $Y2=0
cc_1347 N_D[1]_c_1472_n N_A_405_918#_c_7017_n 0.00208088f $X=5.095 $Y=4.28 $X2=0
+ $Y2=0
cc_1348 N_D[1]_c_1473_n N_A_405_918#_c_7017_n 0.018367f $X=5.84 $Y=4.28 $X2=0
+ $Y2=0
cc_1349 N_D[1]_M1059_g N_A_405_918#_c_7018_n 5.22365e-19 $X=4.98 $Y=4.88 $X2=0
+ $Y2=0
cc_1350 N_D[1]_M1068_g N_A_405_918#_c_7018_n 0.00748012f $X=5.5 $Y=4.88 $X2=0
+ $Y2=0
cc_1351 N_D[1]_M1157_g N_A_405_918#_c_7018_n 0.0073679f $X=5.92 $Y=4.88 $X2=0
+ $Y2=0
cc_1352 N_D[1]_c_1473_n N_A_405_918#_c_7018_n 0.021403f $X=5.84 $Y=4.28 $X2=0
+ $Y2=0
cc_1353 N_D[1]_c_1474_n N_A_405_918#_c_7018_n 0.00208088f $X=5.945 $Y=4.28 $X2=0
+ $Y2=0
cc_1354 N_D[2]_M1071_g N_D[3]_M1000_g 0.0130744f $X=6.475 $Y=1.985 $X2=0 $Y2=0
cc_1355 N_D[2]_M1090_g N_D[3]_M1076_g 0.0130744f $X=6.945 $Y=1.985 $X2=0 $Y2=0
cc_1356 N_D[2]_M1118_g N_D[3]_M1095_g 0.0130744f $X=7.415 $Y=1.985 $X2=0 $Y2=0
cc_1357 N_D[2]_M1158_g N_D[3]_M1120_g 0.0130744f $X=7.885 $Y=1.985 $X2=0 $Y2=0
cc_1358 N_D[2]_M1071_g N_VPWR_c_3594_n 0.00207065f $X=6.475 $Y=1.985 $X2=0 $Y2=0
cc_1359 N_D[2]_M1090_g N_VPWR_c_3596_n 0.00208662f $X=6.945 $Y=1.985 $X2=0 $Y2=0
cc_1360 N_D[2]_M1118_g N_VPWR_c_3596_n 0.00208662f $X=7.415 $Y=1.985 $X2=0 $Y2=0
cc_1361 N_D[2]_M1118_g N_VPWR_c_3598_n 0.0035837f $X=7.415 $Y=1.985 $X2=0 $Y2=0
cc_1362 N_D[2]_M1158_g N_VPWR_c_3598_n 0.0035837f $X=7.885 $Y=1.985 $X2=0 $Y2=0
cc_1363 N_D[2]_M1158_g N_VPWR_c_3599_n 0.00389633f $X=7.885 $Y=1.985 $X2=0 $Y2=0
cc_1364 N_D[2]_M1071_g N_VPWR_c_3643_n 0.0035837f $X=6.475 $Y=1.985 $X2=0 $Y2=0
cc_1365 N_D[2]_M1090_g N_VPWR_c_3643_n 0.0035837f $X=6.945 $Y=1.985 $X2=0 $Y2=0
cc_1366 N_D[2]_M1071_g N_VPWR_c_3661_n 0.00579371f $X=6.475 $Y=1.985 $X2=0 $Y2=0
cc_1367 N_D[2]_M1090_g N_VPWR_c_3661_n 0.00445624f $X=6.945 $Y=1.985 $X2=0 $Y2=0
cc_1368 N_D[2]_M1118_g N_VPWR_c_3661_n 0.00445624f $X=7.415 $Y=1.985 $X2=0 $Y2=0
cc_1369 N_D[2]_M1158_g N_VPWR_c_3661_n 0.00573859f $X=7.885 $Y=1.985 $X2=0 $Y2=0
cc_1370 N_D[2]_M1071_g N_Z_c_4644_n 0.00470782f $X=6.475 $Y=1.985 $X2=0 $Y2=0
cc_1371 N_D[2]_M1090_g N_Z_c_4644_n 0.00306964f $X=6.945 $Y=1.985 $X2=0 $Y2=0
cc_1372 N_D[2]_M1118_g N_Z_c_4644_n 0.00306964f $X=7.415 $Y=1.985 $X2=0 $Y2=0
cc_1373 N_D[2]_M1158_g N_Z_c_4644_n 0.00311896f $X=7.885 $Y=1.985 $X2=0 $Y2=0
cc_1374 N_D[2]_c_1570_n N_Z_c_4644_n 0.00846955f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_1375 N_D[2]_M1090_g N_A_1313_297#_c_5507_n 0.00916655f $X=6.945 $Y=1.985
+ $X2=0 $Y2=0
cc_1376 N_D[2]_M1118_g N_A_1313_297#_c_5507_n 0.00916655f $X=7.415 $Y=1.985
+ $X2=0 $Y2=0
cc_1377 N_D[2]_c_1568_n N_A_1313_297#_c_5507_n 7.15862e-19 $X=7.325 $Y=1.16
+ $X2=0 $Y2=0
cc_1378 N_D[2]_c_1570_n N_A_1313_297#_c_5507_n 0.0387168f $X=7.6 $Y=1.16 $X2=0
+ $Y2=0
cc_1379 N_D[2]_M1158_g N_A_1313_297#_c_5502_n 0.013247f $X=7.885 $Y=1.985 $X2=0
+ $Y2=0
cc_1380 N_D[2]_M1071_g N_A_1313_297#_c_5512_n 0.002088f $X=6.475 $Y=1.985 $X2=0
+ $Y2=0
cc_1381 N_D[2]_M1090_g N_A_1313_297#_c_5512_n 5.79575e-19 $X=6.945 $Y=1.985
+ $X2=0 $Y2=0
cc_1382 N_D[2]_c_1569_n N_A_1313_297#_c_5512_n 8.03631e-19 $X=7.035 $Y=1.16
+ $X2=0 $Y2=0
cc_1383 N_D[2]_c_1570_n N_A_1313_297#_c_5512_n 0.0217153f $X=7.6 $Y=1.16 $X2=0
+ $Y2=0
cc_1384 N_D[2]_M1118_g N_A_1313_297#_c_5516_n 5.79575e-19 $X=7.415 $Y=1.985
+ $X2=0 $Y2=0
cc_1385 N_D[2]_M1158_g N_A_1313_297#_c_5516_n 8.61029e-19 $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_1386 N_D[2]_c_1570_n N_A_1313_297#_c_5516_n 0.0191156f $X=7.6 $Y=1.16 $X2=0
+ $Y2=0
cc_1387 N_D[2]_c_1571_n N_A_1313_297#_c_5516_n 8.03631e-19 $X=7.885 $Y=1.16
+ $X2=0 $Y2=0
cc_1388 N_D[2]_M1090_g N_A_1313_297#_c_5520_n 0.00232998f $X=6.945 $Y=1.985
+ $X2=0 $Y2=0
cc_1389 N_D[2]_M1118_g N_A_1313_297#_c_5520_n 0.00232998f $X=7.415 $Y=1.985
+ $X2=0 $Y2=0
cc_1390 N_D[2]_M1158_g N_A_1313_297#_c_5503_n 0.00232998f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_1391 N_D[2]_M1071_g N_A_1313_297#_c_5523_n 0.00819194f $X=6.475 $Y=1.985
+ $X2=0 $Y2=0
cc_1392 N_D[2]_M1090_g N_A_1313_297#_c_5523_n 0.00911325f $X=6.945 $Y=1.985
+ $X2=0 $Y2=0
cc_1393 N_D[2]_M1118_g N_A_1313_297#_c_5523_n 7.05028e-19 $X=7.415 $Y=1.985
+ $X2=0 $Y2=0
cc_1394 N_D[2]_M1090_g N_A_1313_297#_c_5526_n 7.05028e-19 $X=6.945 $Y=1.985
+ $X2=0 $Y2=0
cc_1395 N_D[2]_M1118_g N_A_1313_297#_c_5526_n 0.00911325f $X=7.415 $Y=1.985
+ $X2=0 $Y2=0
cc_1396 N_D[2]_M1158_g N_A_1313_297#_c_5526_n 0.00977623f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_1397 N_D[2]_M1158_g N_A_1313_297#_c_5504_n 0.00333758f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_1398 N_D[2]_M1013_g N_VGND_c_6274_n 0.0058918f $X=6.5 $Y=0.56 $X2=0 $Y2=0
cc_1399 N_D[2]_M1013_g N_VGND_c_6276_n 2.64031e-19 $X=6.5 $Y=0.56 $X2=0 $Y2=0
cc_1400 N_D[2]_M1037_g N_VGND_c_6276_n 0.00166854f $X=6.92 $Y=0.56 $X2=0 $Y2=0
cc_1401 N_D[2]_M1069_g N_VGND_c_6276_n 0.0019152f $X=7.44 $Y=0.56 $X2=0 $Y2=0
cc_1402 N_D[2]_M1069_g N_VGND_c_6278_n 0.00430643f $X=7.44 $Y=0.56 $X2=0 $Y2=0
cc_1403 N_D[2]_M1150_g N_VGND_c_6278_n 0.00422241f $X=7.86 $Y=0.56 $X2=0 $Y2=0
cc_1404 N_D[2]_M1069_g N_VGND_c_6280_n 2.6376e-19 $X=7.44 $Y=0.56 $X2=0 $Y2=0
cc_1405 N_D[2]_M1150_g N_VGND_c_6280_n 0.00321269f $X=7.86 $Y=0.56 $X2=0 $Y2=0
cc_1406 N_D[2]_M1013_g N_VGND_c_6344_n 0.00551064f $X=6.5 $Y=0.56 $X2=0 $Y2=0
cc_1407 N_D[2]_M1037_g N_VGND_c_6344_n 0.00422241f $X=6.92 $Y=0.56 $X2=0 $Y2=0
cc_1408 N_D[2]_M1013_g N_VGND_c_6370_n 0.0101978f $X=6.5 $Y=0.56 $X2=0 $Y2=0
cc_1409 N_D[2]_M1037_g N_VGND_c_6370_n 0.00593887f $X=6.92 $Y=0.56 $X2=0 $Y2=0
cc_1410 N_D[2]_M1069_g N_VGND_c_6370_n 0.00624811f $X=7.44 $Y=0.56 $X2=0 $Y2=0
cc_1411 N_D[2]_M1150_g N_VGND_c_6370_n 0.00702263f $X=7.86 $Y=0.56 $X2=0 $Y2=0
cc_1412 N_D[2]_M1013_g N_A_1315_47#_c_7100_n 0.00514241f $X=6.5 $Y=0.56 $X2=0
+ $Y2=0
cc_1413 N_D[2]_M1037_g N_A_1315_47#_c_7100_n 0.00661134f $X=6.92 $Y=0.56 $X2=0
+ $Y2=0
cc_1414 N_D[2]_M1069_g N_A_1315_47#_c_7100_n 5.22365e-19 $X=7.44 $Y=0.56 $X2=0
+ $Y2=0
cc_1415 N_D[2]_M1037_g N_A_1315_47#_c_7103_n 0.00899636f $X=6.92 $Y=0.56 $X2=0
+ $Y2=0
cc_1416 N_D[2]_M1069_g N_A_1315_47#_c_7103_n 0.00900364f $X=7.44 $Y=0.56 $X2=0
+ $Y2=0
cc_1417 N_D[2]_c_1568_n N_A_1315_47#_c_7103_n 0.00463549f $X=7.325 $Y=1.16 $X2=0
+ $Y2=0
cc_1418 N_D[2]_c_1570_n N_A_1315_47#_c_7103_n 0.0394855f $X=7.6 $Y=1.16 $X2=0
+ $Y2=0
cc_1419 N_D[2]_M1013_g N_A_1315_47#_c_7092_n 0.00222549f $X=6.5 $Y=0.56 $X2=0
+ $Y2=0
cc_1420 N_D[2]_M1037_g N_A_1315_47#_c_7092_n 8.68782e-19 $X=6.92 $Y=0.56 $X2=0
+ $Y2=0
cc_1421 N_D[2]_c_1569_n N_A_1315_47#_c_7092_n 0.00208088f $X=7.035 $Y=1.16 $X2=0
+ $Y2=0
cc_1422 N_D[2]_c_1570_n N_A_1315_47#_c_7092_n 0.021403f $X=7.6 $Y=1.16 $X2=0
+ $Y2=0
cc_1423 N_D[2]_M1037_g N_A_1315_47#_c_7111_n 5.22365e-19 $X=6.92 $Y=0.56 $X2=0
+ $Y2=0
cc_1424 N_D[2]_M1069_g N_A_1315_47#_c_7111_n 0.00661764f $X=7.44 $Y=0.56 $X2=0
+ $Y2=0
cc_1425 N_D[2]_M1150_g N_A_1315_47#_c_7111_n 0.00699463f $X=7.86 $Y=0.56 $X2=0
+ $Y2=0
cc_1426 N_D[2]_M1150_g N_A_1315_47#_c_7093_n 0.0121912f $X=7.86 $Y=0.56 $X2=0
+ $Y2=0
cc_1427 N_D[2]_M1150_g N_A_1315_47#_c_7094_n 0.00261078f $X=7.86 $Y=0.56 $X2=0
+ $Y2=0
cc_1428 N_D[2]_M1069_g N_A_1315_47#_c_7099_n 8.68782e-19 $X=7.44 $Y=0.56 $X2=0
+ $Y2=0
cc_1429 N_D[2]_M1150_g N_A_1315_47#_c_7099_n 0.00128201f $X=7.86 $Y=0.56 $X2=0
+ $Y2=0
cc_1430 N_D[2]_c_1570_n N_A_1315_47#_c_7099_n 0.018367f $X=7.6 $Y=1.16 $X2=0
+ $Y2=0
cc_1431 N_D[2]_c_1571_n N_A_1315_47#_c_7099_n 0.00208088f $X=7.885 $Y=1.16 $X2=0
+ $Y2=0
cc_1432 N_D[3]_M1000_g N_VPWR_c_3595_n 0.00207065f $X=6.475 $Y=3.455 $X2=0 $Y2=0
cc_1433 N_D[3]_M1076_g N_VPWR_c_3597_n 0.00208662f $X=6.945 $Y=3.455 $X2=0 $Y2=0
cc_1434 N_D[3]_M1095_g N_VPWR_c_3597_n 0.00208662f $X=7.415 $Y=3.455 $X2=0 $Y2=0
cc_1435 N_D[3]_M1095_g N_VPWR_c_3598_n 0.0035837f $X=7.415 $Y=3.455 $X2=0 $Y2=0
cc_1436 N_D[3]_M1120_g N_VPWR_c_3598_n 0.0035837f $X=7.885 $Y=3.455 $X2=0 $Y2=0
cc_1437 N_D[3]_M1120_g N_VPWR_c_3600_n 0.00389633f $X=7.885 $Y=3.455 $X2=0 $Y2=0
cc_1438 N_D[3]_M1000_g N_VPWR_c_3643_n 0.0035837f $X=6.475 $Y=3.455 $X2=0 $Y2=0
cc_1439 N_D[3]_M1076_g N_VPWR_c_3643_n 0.0035837f $X=6.945 $Y=3.455 $X2=0 $Y2=0
cc_1440 N_D[3]_M1000_g N_VPWR_c_3661_n 0.00579371f $X=6.475 $Y=3.455 $X2=0 $Y2=0
cc_1441 N_D[3]_M1076_g N_VPWR_c_3661_n 0.00445624f $X=6.945 $Y=3.455 $X2=0 $Y2=0
cc_1442 N_D[3]_M1095_g N_VPWR_c_3661_n 0.00445624f $X=7.415 $Y=3.455 $X2=0 $Y2=0
cc_1443 N_D[3]_M1120_g N_VPWR_c_3661_n 0.00573859f $X=7.885 $Y=3.455 $X2=0 $Y2=0
cc_1444 N_D[3]_M1000_g N_Z_c_4645_n 0.00470782f $X=6.475 $Y=3.455 $X2=0 $Y2=0
cc_1445 N_D[3]_M1076_g N_Z_c_4645_n 0.00306964f $X=6.945 $Y=3.455 $X2=0 $Y2=0
cc_1446 N_D[3]_M1095_g N_Z_c_4645_n 0.00306964f $X=7.415 $Y=3.455 $X2=0 $Y2=0
cc_1447 N_D[3]_M1120_g N_Z_c_4645_n 0.00311896f $X=7.885 $Y=3.455 $X2=0 $Y2=0
cc_1448 N_D[3]_c_1671_n N_Z_c_4645_n 0.00846955f $X=7.6 $Y=4.28 $X2=0 $Y2=0
cc_1449 N_D[3]_M1076_g N_A_1313_591#_c_5635_n 0.00916655f $X=6.945 $Y=3.455
+ $X2=0 $Y2=0
cc_1450 N_D[3]_M1095_g N_A_1313_591#_c_5635_n 0.00916655f $X=7.415 $Y=3.455
+ $X2=0 $Y2=0
cc_1451 N_D[3]_c_1669_n N_A_1313_591#_c_5635_n 7.15862e-19 $X=7.325 $Y=4.28
+ $X2=0 $Y2=0
cc_1452 N_D[3]_c_1671_n N_A_1313_591#_c_5635_n 0.0387168f $X=7.6 $Y=4.28 $X2=0
+ $Y2=0
cc_1453 N_D[3]_M1120_g N_A_1313_591#_c_5630_n 0.013247f $X=7.885 $Y=3.455 $X2=0
+ $Y2=0
cc_1454 N_D[3]_M1000_g N_A_1313_591#_c_5640_n 0.002088f $X=6.475 $Y=3.455 $X2=0
+ $Y2=0
cc_1455 N_D[3]_M1076_g N_A_1313_591#_c_5640_n 5.79575e-19 $X=6.945 $Y=3.455
+ $X2=0 $Y2=0
cc_1456 N_D[3]_c_1670_n N_A_1313_591#_c_5640_n 8.03631e-19 $X=7.035 $Y=4.28
+ $X2=0 $Y2=0
cc_1457 N_D[3]_c_1671_n N_A_1313_591#_c_5640_n 0.0217153f $X=7.6 $Y=4.28 $X2=0
+ $Y2=0
cc_1458 N_D[3]_M1095_g N_A_1313_591#_c_5644_n 5.79575e-19 $X=7.415 $Y=3.455
+ $X2=0 $Y2=0
cc_1459 N_D[3]_M1120_g N_A_1313_591#_c_5644_n 8.61029e-19 $X=7.885 $Y=3.455
+ $X2=0 $Y2=0
cc_1460 N_D[3]_c_1671_n N_A_1313_591#_c_5644_n 0.0191156f $X=7.6 $Y=4.28 $X2=0
+ $Y2=0
cc_1461 N_D[3]_c_1672_n N_A_1313_591#_c_5644_n 8.03631e-19 $X=7.885 $Y=4.28
+ $X2=0 $Y2=0
cc_1462 N_D[3]_M1076_g N_A_1313_591#_c_5648_n 0.00232998f $X=6.945 $Y=3.455
+ $X2=0 $Y2=0
cc_1463 N_D[3]_M1095_g N_A_1313_591#_c_5648_n 0.00232998f $X=7.415 $Y=3.455
+ $X2=0 $Y2=0
cc_1464 N_D[3]_M1120_g N_A_1313_591#_c_5631_n 0.00232998f $X=7.885 $Y=3.455
+ $X2=0 $Y2=0
cc_1465 N_D[3]_M1000_g N_A_1313_591#_c_5651_n 0.00819194f $X=6.475 $Y=3.455
+ $X2=0 $Y2=0
cc_1466 N_D[3]_M1076_g N_A_1313_591#_c_5651_n 0.00911325f $X=6.945 $Y=3.455
+ $X2=0 $Y2=0
cc_1467 N_D[3]_M1095_g N_A_1313_591#_c_5651_n 7.05028e-19 $X=7.415 $Y=3.455
+ $X2=0 $Y2=0
cc_1468 N_D[3]_M1076_g N_A_1313_591#_c_5654_n 7.05028e-19 $X=6.945 $Y=3.455
+ $X2=0 $Y2=0
cc_1469 N_D[3]_M1095_g N_A_1313_591#_c_5654_n 0.00911325f $X=7.415 $Y=3.455
+ $X2=0 $Y2=0
cc_1470 N_D[3]_M1120_g N_A_1313_591#_c_5654_n 0.00977623f $X=7.885 $Y=3.455
+ $X2=0 $Y2=0
cc_1471 N_D[3]_M1120_g N_A_1313_591#_c_5632_n 0.00333758f $X=7.885 $Y=3.455
+ $X2=0 $Y2=0
cc_1472 N_D[3]_M1015_g N_VGND_c_6275_n 0.0058918f $X=6.5 $Y=4.88 $X2=0 $Y2=0
cc_1473 N_D[3]_M1015_g N_VGND_c_6277_n 2.64031e-19 $X=6.5 $Y=4.88 $X2=0 $Y2=0
cc_1474 N_D[3]_M1047_g N_VGND_c_6277_n 0.00166854f $X=6.92 $Y=4.88 $X2=0 $Y2=0
cc_1475 N_D[3]_M1104_g N_VGND_c_6277_n 0.0019152f $X=7.44 $Y=4.88 $X2=0 $Y2=0
cc_1476 N_D[3]_M1104_g N_VGND_c_6279_n 0.00430643f $X=7.44 $Y=4.88 $X2=0 $Y2=0
cc_1477 N_D[3]_M1136_g N_VGND_c_6279_n 0.00422241f $X=7.86 $Y=4.88 $X2=0 $Y2=0
cc_1478 N_D[3]_M1104_g N_VGND_c_6281_n 2.6376e-19 $X=7.44 $Y=4.88 $X2=0 $Y2=0
cc_1479 N_D[3]_M1136_g N_VGND_c_6281_n 0.00321269f $X=7.86 $Y=4.88 $X2=0 $Y2=0
cc_1480 N_D[3]_M1015_g N_VGND_c_6345_n 0.00551064f $X=6.5 $Y=4.88 $X2=0 $Y2=0
cc_1481 N_D[3]_M1047_g N_VGND_c_6345_n 0.00422241f $X=6.92 $Y=4.88 $X2=0 $Y2=0
cc_1482 N_D[3]_M1015_g N_VGND_c_6371_n 0.0101978f $X=6.5 $Y=4.88 $X2=0 $Y2=0
cc_1483 N_D[3]_M1047_g N_VGND_c_6371_n 0.00593887f $X=6.92 $Y=4.88 $X2=0 $Y2=0
cc_1484 N_D[3]_M1104_g N_VGND_c_6371_n 0.00624811f $X=7.44 $Y=4.88 $X2=0 $Y2=0
cc_1485 N_D[3]_M1136_g N_VGND_c_6371_n 0.00702263f $X=7.86 $Y=4.88 $X2=0 $Y2=0
cc_1486 N_D[3]_M1047_g N_A_1315_911#_c_7183_n 0.00899636f $X=6.92 $Y=4.88 $X2=0
+ $Y2=0
cc_1487 N_D[3]_M1104_g N_A_1315_911#_c_7183_n 0.00900364f $X=7.44 $Y=4.88 $X2=0
+ $Y2=0
cc_1488 N_D[3]_c_1669_n N_A_1315_911#_c_7183_n 0.00463549f $X=7.325 $Y=4.28
+ $X2=0 $Y2=0
cc_1489 N_D[3]_c_1671_n N_A_1315_911#_c_7183_n 0.0394855f $X=7.6 $Y=4.28 $X2=0
+ $Y2=0
cc_1490 N_D[3]_M1136_g N_A_1315_911#_c_7175_n 0.0121912f $X=7.86 $Y=4.88 $X2=0
+ $Y2=0
cc_1491 N_D[3]_M1136_g N_A_1315_911#_c_7176_n 0.00261078f $X=7.86 $Y=4.88 $X2=0
+ $Y2=0
cc_1492 N_D[3]_M1015_g N_A_1315_911#_c_7181_n 0.0073679f $X=6.5 $Y=4.88 $X2=0
+ $Y2=0
cc_1493 N_D[3]_M1047_g N_A_1315_911#_c_7181_n 0.00748012f $X=6.92 $Y=4.88 $X2=0
+ $Y2=0
cc_1494 N_D[3]_M1104_g N_A_1315_911#_c_7181_n 5.22365e-19 $X=7.44 $Y=4.88 $X2=0
+ $Y2=0
cc_1495 N_D[3]_c_1670_n N_A_1315_911#_c_7181_n 0.00208088f $X=7.035 $Y=4.28
+ $X2=0 $Y2=0
cc_1496 N_D[3]_c_1671_n N_A_1315_911#_c_7181_n 0.021403f $X=7.6 $Y=4.28 $X2=0
+ $Y2=0
cc_1497 N_D[3]_M1047_g N_A_1315_911#_c_7182_n 5.22365e-19 $X=6.92 $Y=4.88 $X2=0
+ $Y2=0
cc_1498 N_D[3]_M1104_g N_A_1315_911#_c_7182_n 0.00748643f $X=7.44 $Y=4.88 $X2=0
+ $Y2=0
cc_1499 N_D[3]_M1136_g N_A_1315_911#_c_7182_n 0.00827664f $X=7.86 $Y=4.88 $X2=0
+ $Y2=0
cc_1500 N_D[3]_c_1671_n N_A_1315_911#_c_7182_n 0.018367f $X=7.6 $Y=4.28 $X2=0
+ $Y2=0
cc_1501 N_D[3]_c_1672_n N_A_1315_911#_c_7182_n 0.00208088f $X=7.885 $Y=4.28
+ $X2=0 $Y2=0
cc_1502 N_A_1755_265#_c_1765_n N_A_1755_793#_c_1884_n 0.0129371f $X=8.875
+ $Y=1.475 $X2=0 $Y2=0
cc_1503 N_A_1755_265#_c_1768_n N_A_1755_793#_c_1887_n 0.0129371f $X=9.345
+ $Y=1.475 $X2=0 $Y2=0
cc_1504 N_A_1755_265#_c_1770_n N_A_1755_793#_c_1889_n 0.0129371f $X=9.815
+ $Y=1.475 $X2=0 $Y2=0
cc_1505 N_A_1755_265#_c_1772_n N_A_1755_793#_c_1891_n 0.0129371f $X=10.285
+ $Y=1.475 $X2=0 $Y2=0
cc_1506 N_A_1755_265#_c_1767_n N_S[2]_c_2002_n 0.00507426f $X=8.965 $Y=1.4
+ $X2=-0.19 $Y2=-0.24
cc_1507 N_A_1755_265#_c_1766_n N_S[2]_c_2005_n 0.00509391f $X=9.255 $Y=1.4 $X2=0
+ $Y2=0
cc_1508 N_A_1755_265#_c_1769_n N_S[2]_c_2007_n 0.00509204f $X=9.725 $Y=1.4 $X2=0
+ $Y2=0
cc_1509 N_A_1755_265#_c_1771_n N_S[2]_c_2009_n 0.00507688f $X=10.195 $Y=1.4
+ $X2=0 $Y2=0
cc_1510 N_A_1755_265#_c_1760_n N_S[2]_c_2011_n 6.53442e-19 $X=11.565 $Y=0.445
+ $X2=0 $Y2=0
cc_1511 N_A_1755_265#_c_1758_n N_S[2]_c_2013_n 0.0103812f $X=11.4 $Y=1.23 $X2=0
+ $Y2=0
cc_1512 N_A_1755_265#_c_1759_n N_S[2]_c_2013_n 0.0179529f $X=10.855 $Y=1.23
+ $X2=0 $Y2=0
cc_1513 N_A_1755_265#_c_1758_n N_S[2]_c_2014_n 0.0206368f $X=11.4 $Y=1.23 $X2=0
+ $Y2=0
cc_1514 N_A_1755_265#_c_1759_n N_S[2]_c_2014_n 0.0175393f $X=10.855 $Y=1.23
+ $X2=0 $Y2=0
cc_1515 N_A_1755_265#_c_1761_n N_S[2]_c_2014_n 0.0085951f $X=11.485 $Y=1.065
+ $X2=0 $Y2=0
cc_1516 N_A_1755_265#_c_1763_n N_S[2]_c_2014_n 0.00322131f $X=11.485 $Y=1.23
+ $X2=0 $Y2=0
cc_1517 N_A_1755_265#_c_1779_n N_S[2]_c_2014_n 0.00255921f $X=11.565 $Y=1.605
+ $X2=0 $Y2=0
cc_1518 N_A_1755_265#_c_1764_n N_S[2]_c_2014_n 0.00262132f $X=10.605 $Y=1.23
+ $X2=0 $Y2=0
cc_1519 N_A_1755_265#_c_1777_n N_S[2]_c_2025_n 0.0118698f $X=11.565 $Y=1.77
+ $X2=0 $Y2=0
cc_1520 N_A_1755_265#_c_1779_n N_S[2]_c_2025_n 0.00762115f $X=11.565 $Y=1.605
+ $X2=0 $Y2=0
cc_1521 N_A_1755_265#_c_1760_n N_S[2]_c_2015_n 0.00603996f $X=11.565 $Y=0.445
+ $X2=0 $Y2=0
cc_1522 N_A_1755_265#_c_1762_n N_S[2]_c_2015_n 9.67113e-19 $X=11.525 $Y=0.825
+ $X2=0 $Y2=0
cc_1523 N_A_1755_265#_c_1761_n N_S[2]_c_2016_n 0.00429801f $X=11.485 $Y=1.065
+ $X2=0 $Y2=0
cc_1524 N_A_1755_265#_c_1762_n N_S[2]_c_2016_n 0.0111895f $X=11.525 $Y=0.825
+ $X2=0 $Y2=0
cc_1525 N_A_1755_265#_c_1760_n N_S[2]_c_2017_n 0.00207203f $X=11.565 $Y=0.445
+ $X2=0 $Y2=0
cc_1526 N_A_1755_265#_c_1761_n N_S[2]_c_2018_n 0.00289358f $X=11.485 $Y=1.065
+ $X2=0 $Y2=0
cc_1527 N_A_1755_265#_c_1777_n N_S[2]_c_2018_n 0.0128834f $X=11.565 $Y=1.77
+ $X2=0 $Y2=0
cc_1528 N_A_1755_265#_c_1763_n N_S[2]_c_2018_n 0.00416423f $X=11.485 $Y=1.23
+ $X2=0 $Y2=0
cc_1529 N_A_1755_265#_c_1779_n N_S[2]_c_2018_n 0.00454075f $X=11.565 $Y=1.605
+ $X2=0 $Y2=0
cc_1530 N_A_1755_265#_c_1761_n N_S[2]_c_2022_n 0.00268644f $X=11.485 $Y=1.065
+ $X2=0 $Y2=0
cc_1531 N_A_1755_265#_c_1762_n N_S[2]_c_2022_n 0.00426435f $X=11.525 $Y=0.825
+ $X2=0 $Y2=0
cc_1532 N_A_1755_265#_c_1761_n S[2] 0.00541767f $X=11.485 $Y=1.065 $X2=0 $Y2=0
cc_1533 N_A_1755_265#_c_1763_n S[2] 0.0228692f $X=11.485 $Y=1.23 $X2=0 $Y2=0
cc_1534 N_A_1755_265#_c_1765_n N_VPWR_c_3599_n 0.00324472f $X=8.875 $Y=1.475
+ $X2=0 $Y2=0
cc_1535 N_A_1755_265#_c_1772_n N_VPWR_c_3601_n 0.00367058f $X=10.285 $Y=1.475
+ $X2=0 $Y2=0
cc_1536 N_A_1755_265#_c_1758_n N_VPWR_c_3601_n 0.0193185f $X=11.4 $Y=1.23 $X2=0
+ $Y2=0
cc_1537 N_A_1755_265#_c_1759_n N_VPWR_c_3601_n 6.4101e-19 $X=10.855 $Y=1.23
+ $X2=0 $Y2=0
cc_1538 N_A_1755_265#_c_1777_n N_VPWR_c_3601_n 0.0316788f $X=11.565 $Y=1.77
+ $X2=0 $Y2=0
cc_1539 N_A_1755_265#_c_1777_n N_VPWR_c_3603_n 0.0356181f $X=11.565 $Y=1.77
+ $X2=0 $Y2=0
cc_1540 N_A_1755_265#_c_1777_n N_VPWR_c_3632_n 0.0233824f $X=11.565 $Y=1.77
+ $X2=0 $Y2=0
cc_1541 N_A_1755_265#_c_1765_n N_VPWR_c_3661_n 0.00473731f $X=8.875 $Y=1.475
+ $X2=0 $Y2=0
cc_1542 N_A_1755_265#_c_1768_n N_VPWR_c_3661_n 0.00362156f $X=9.345 $Y=1.475
+ $X2=0 $Y2=0
cc_1543 N_A_1755_265#_c_1770_n N_VPWR_c_3661_n 0.00362156f $X=9.815 $Y=1.475
+ $X2=0 $Y2=0
cc_1544 N_A_1755_265#_c_1772_n N_VPWR_c_3661_n 0.00473731f $X=10.285 $Y=1.475
+ $X2=0 $Y2=0
cc_1545 N_A_1755_265#_c_1777_n N_VPWR_c_3661_n 0.00593513f $X=11.565 $Y=1.77
+ $X2=0 $Y2=0
cc_1546 N_A_1755_265#_c_1769_n N_Z_c_4594_n 0.00762343f $X=9.725 $Y=1.4 $X2=0
+ $Y2=0
cc_1547 N_A_1755_265#_c_1773_n N_Z_c_4594_n 0.00704092f $X=9.345 $Y=1.4 $X2=0
+ $Y2=0
cc_1548 N_A_1755_265#_c_1767_n N_Z_c_4615_n 0.00248496f $X=8.965 $Y=1.4 $X2=0
+ $Y2=0
cc_1549 N_A_1755_265#_c_1766_n N_Z_c_4618_n 0.00678861f $X=9.255 $Y=1.4 $X2=0
+ $Y2=0
cc_1550 N_A_1755_265#_c_1767_n N_Z_c_4618_n 0.00239476f $X=8.965 $Y=1.4 $X2=0
+ $Y2=0
cc_1551 N_A_1755_265#_c_1773_n N_Z_c_4618_n 2.98555e-19 $X=9.345 $Y=1.4 $X2=0
+ $Y2=0
cc_1552 N_A_1755_265#_c_1769_n N_Z_c_4620_n 0.00145542f $X=9.725 $Y=1.4 $X2=0
+ $Y2=0
cc_1553 N_A_1755_265#_c_1771_n N_Z_c_4620_n 0.00597584f $X=10.195 $Y=1.4 $X2=0
+ $Y2=0
cc_1554 N_A_1755_265#_c_1774_n N_Z_c_4620_n 0.00909323f $X=9.815 $Y=1.4 $X2=0
+ $Y2=0
cc_1555 N_A_1755_265#_c_1758_n N_Z_c_4620_n 0.0266078f $X=11.4 $Y=1.23 $X2=0
+ $Y2=0
cc_1556 N_A_1755_265#_c_1764_n N_Z_c_4620_n 0.00747617f $X=10.605 $Y=1.23 $X2=0
+ $Y2=0
cc_1557 N_A_1755_265#_c_1765_n N_Z_c_4644_n 0.00834829f $X=8.875 $Y=1.475 $X2=0
+ $Y2=0
cc_1558 N_A_1755_265#_c_1772_n N_Z_c_4646_n 0.00795576f $X=10.285 $Y=1.475 $X2=0
+ $Y2=0
cc_1559 N_A_1755_265#_c_1758_n N_Z_c_4646_n 0.0186685f $X=11.4 $Y=1.23 $X2=0
+ $Y2=0
cc_1560 N_A_1755_265#_c_1777_n N_Z_c_4646_n 0.0329704f $X=11.565 $Y=1.77 $X2=0
+ $Y2=0
cc_1561 N_A_1755_265#_c_1764_n N_Z_c_4646_n 2.19754e-19 $X=10.605 $Y=1.23 $X2=0
+ $Y2=0
cc_1562 N_A_1755_265#_c_1768_n Z 0.00372458f $X=9.345 $Y=1.475 $X2=0 $Y2=0
cc_1563 N_A_1755_265#_c_1770_n Z 0.00372248f $X=9.815 $Y=1.475 $X2=0 $Y2=0
cc_1564 N_A_1755_265#_c_1765_n N_Z_c_4652_n 0.0199111f $X=8.875 $Y=1.475 $X2=0
+ $Y2=0
cc_1565 N_A_1755_265#_c_1766_n N_Z_c_4652_n 0.00560592f $X=9.255 $Y=1.4 $X2=0
+ $Y2=0
cc_1566 N_A_1755_265#_c_1767_n N_Z_c_4652_n 0.00474497f $X=8.965 $Y=1.4 $X2=0
+ $Y2=0
cc_1567 N_A_1755_265#_c_1768_n N_Z_c_4652_n 0.0181262f $X=9.345 $Y=1.475 $X2=0
+ $Y2=0
cc_1568 N_A_1755_265#_c_1770_n N_Z_c_4652_n 9.74366e-19 $X=9.815 $Y=1.475 $X2=0
+ $Y2=0
cc_1569 N_A_1755_265#_c_1773_n N_Z_c_4652_n 0.00415268f $X=9.345 $Y=1.4 $X2=0
+ $Y2=0
cc_1570 N_A_1755_265#_c_1768_n N_Z_c_4653_n 9.74366e-19 $X=9.345 $Y=1.475 $X2=0
+ $Y2=0
cc_1571 N_A_1755_265#_c_1770_n N_Z_c_4653_n 0.0181262f $X=9.815 $Y=1.475 $X2=0
+ $Y2=0
cc_1572 N_A_1755_265#_c_1771_n N_Z_c_4653_n 0.00560592f $X=10.195 $Y=1.4 $X2=0
+ $Y2=0
cc_1573 N_A_1755_265#_c_1772_n N_Z_c_4653_n 0.0221748f $X=10.285 $Y=1.475 $X2=0
+ $Y2=0
cc_1574 N_A_1755_265#_c_1774_n N_Z_c_4653_n 0.00181273f $X=9.815 $Y=1.4 $X2=0
+ $Y2=0
cc_1575 N_A_1755_265#_c_1758_n N_Z_c_4653_n 0.00240108f $X=11.4 $Y=1.23 $X2=0
+ $Y2=0
cc_1576 N_A_1755_265#_c_1764_n N_Z_c_4653_n 0.00425035f $X=10.605 $Y=1.23 $X2=0
+ $Y2=0
cc_1577 N_A_1755_265#_c_1765_n N_A_1313_297#_c_5502_n 0.00151141f $X=8.875
+ $Y=1.475 $X2=0 $Y2=0
cc_1578 N_A_1755_265#_c_1765_n N_A_1313_297#_c_5531_n 0.00307958f $X=8.875
+ $Y=1.475 $X2=0 $Y2=0
cc_1579 N_A_1755_265#_c_1768_n N_A_1313_297#_c_5531_n 0.00307958f $X=9.345
+ $Y=1.475 $X2=0 $Y2=0
cc_1580 N_A_1755_265#_c_1770_n N_A_1313_297#_c_5533_n 0.00307958f $X=9.815
+ $Y=1.475 $X2=0 $Y2=0
cc_1581 N_A_1755_265#_c_1772_n N_A_1313_297#_c_5533_n 0.00307958f $X=10.285
+ $Y=1.475 $X2=0 $Y2=0
cc_1582 N_A_1755_265#_c_1765_n N_A_1313_297#_c_5504_n 0.00554566f $X=8.875
+ $Y=1.475 $X2=0 $Y2=0
cc_1583 N_A_1755_265#_c_1768_n N_A_1313_297#_c_5505_n 0.00210632f $X=9.345
+ $Y=1.475 $X2=0 $Y2=0
cc_1584 N_A_1755_265#_c_1769_n N_A_1313_297#_c_5505_n 0.00251792f $X=9.725
+ $Y=1.4 $X2=0 $Y2=0
cc_1585 N_A_1755_265#_c_1770_n N_A_1313_297#_c_5505_n 0.00210632f $X=9.815
+ $Y=1.475 $X2=0 $Y2=0
cc_1586 N_A_1755_265#_c_1772_n N_A_1313_297#_c_5506_n 0.00499839f $X=10.285
+ $Y=1.475 $X2=0 $Y2=0
cc_1587 N_A_1755_265#_c_1758_n N_A_1313_297#_c_5506_n 0.0218124f $X=11.4 $Y=1.23
+ $X2=0 $Y2=0
cc_1588 N_A_1755_265#_c_1759_n N_A_1313_297#_c_5506_n 5.74251e-19 $X=10.855
+ $Y=1.23 $X2=0 $Y2=0
cc_1589 N_A_1755_265#_c_1764_n N_A_1313_297#_c_5506_n 0.00561627f $X=10.605
+ $Y=1.23 $X2=0 $Y2=0
cc_1590 N_A_1755_265#_c_1758_n N_VGND_c_6282_n 0.0123065f $X=11.4 $Y=1.23 $X2=0
+ $Y2=0
cc_1591 N_A_1755_265#_c_1759_n N_VGND_c_6282_n 2.04129e-19 $X=10.855 $Y=1.23
+ $X2=0 $Y2=0
cc_1592 N_A_1755_265#_c_1760_n N_VGND_c_6320_n 0.0129994f $X=11.565 $Y=0.445
+ $X2=0 $Y2=0
cc_1593 N_A_1755_265#_M1094_s N_VGND_c_6370_n 0.00394793f $X=11.43 $Y=0.235
+ $X2=0 $Y2=0
cc_1594 N_A_1755_265#_c_1760_n N_VGND_c_6370_n 0.00927134f $X=11.565 $Y=0.445
+ $X2=0 $Y2=0
cc_1595 N_A_1755_265#_c_1773_n N_A_1315_47#_c_7120_n 7.0477e-19 $X=9.345 $Y=1.4
+ $X2=0 $Y2=0
cc_1596 N_A_1755_265#_c_1758_n N_A_1315_47#_c_7098_n 0.0028695f $X=11.4 $Y=1.23
+ $X2=0 $Y2=0
cc_1597 N_A_1755_265#_c_1764_n N_A_1315_47#_c_7098_n 0.00589316f $X=10.605
+ $Y=1.23 $X2=0 $Y2=0
cc_1598 N_A_1755_793#_c_1886_n N_S[3]_c_2119_n 0.00507426f $X=8.965 $Y=4.04
+ $X2=-0.19 $Y2=-0.24
cc_1599 N_A_1755_793#_c_1885_n N_S[3]_c_2122_n 0.00509391f $X=9.255 $Y=4.04
+ $X2=0 $Y2=0
cc_1600 N_A_1755_793#_c_1888_n N_S[3]_c_2124_n 0.00509204f $X=9.725 $Y=4.04
+ $X2=0 $Y2=0
cc_1601 N_A_1755_793#_c_1890_n N_S[3]_c_2126_n 0.00507688f $X=10.195 $Y=4.04
+ $X2=0 $Y2=0
cc_1602 N_A_1755_793#_c_1879_n N_S[3]_c_2128_n 6.53442e-19 $X=11.525 $Y=4.74
+ $X2=0 $Y2=0
cc_1603 N_A_1755_793#_c_1877_n N_S[3]_c_2130_n 0.0103812f $X=11.4 $Y=4.21 $X2=0
+ $Y2=0
cc_1604 N_A_1755_793#_c_1878_n N_S[3]_c_2130_n 0.0179529f $X=10.855 $Y=4.21
+ $X2=0 $Y2=0
cc_1605 N_A_1755_793#_c_1897_n N_S[3]_c_2140_n 0.00508008f $X=11.485 $Y=4.045
+ $X2=0 $Y2=0
cc_1606 N_A_1755_793#_c_1883_n N_S[3]_c_2140_n 0.00262132f $X=10.605 $Y=4.21
+ $X2=0 $Y2=0
cc_1607 N_A_1755_793#_c_1877_n N_S[3]_c_2131_n 0.0206368f $X=11.4 $Y=4.21 $X2=0
+ $Y2=0
cc_1608 N_A_1755_793#_c_1878_n N_S[3]_c_2131_n 0.0175393f $X=10.855 $Y=4.21
+ $X2=0 $Y2=0
cc_1609 N_A_1755_793#_c_1897_n N_S[3]_c_2131_n 0.00255921f $X=11.485 $Y=4.045
+ $X2=0 $Y2=0
cc_1610 N_A_1755_793#_c_1881_n N_S[3]_c_2131_n 0.00322131f $X=11.485 $Y=4.21
+ $X2=0 $Y2=0
cc_1611 N_A_1755_793#_c_1882_n N_S[3]_c_2131_n 0.0085951f $X=11.525 $Y=4.615
+ $X2=0 $Y2=0
cc_1612 N_A_1755_793#_c_1896_n N_S[3]_c_2142_n 0.00970559f $X=11.565 $Y=3.14
+ $X2=0 $Y2=0
cc_1613 N_A_1755_793#_c_1897_n N_S[3]_c_2142_n 0.00254107f $X=11.485 $Y=4.045
+ $X2=0 $Y2=0
cc_1614 N_A_1755_793#_c_1898_n N_S[3]_c_2142_n 0.00216424f $X=11.565 $Y=3.835
+ $X2=0 $Y2=0
cc_1615 N_A_1755_793#_c_1879_n N_S[3]_c_2132_n 9.67113e-19 $X=11.525 $Y=4.74
+ $X2=0 $Y2=0
cc_1616 N_A_1755_793#_c_1880_n N_S[3]_c_2132_n 0.00603996f $X=11.565 $Y=4.995
+ $X2=0 $Y2=0
cc_1617 N_A_1755_793#_c_1879_n N_S[3]_c_2133_n 0.0111895f $X=11.525 $Y=4.74
+ $X2=0 $Y2=0
cc_1618 N_A_1755_793#_c_1882_n N_S[3]_c_2133_n 0.00429801f $X=11.525 $Y=4.615
+ $X2=0 $Y2=0
cc_1619 N_A_1755_793#_c_1897_n N_S[3]_c_2134_n 0.00336772f $X=11.485 $Y=4.045
+ $X2=0 $Y2=0
cc_1620 N_A_1755_793#_c_1879_n N_S[3]_c_2134_n 0.00207203f $X=11.525 $Y=4.74
+ $X2=0 $Y2=0
cc_1621 N_A_1755_793#_c_1898_n N_S[3]_c_2134_n 5.48523e-19 $X=11.565 $Y=3.835
+ $X2=0 $Y2=0
cc_1622 N_A_1755_793#_c_1881_n N_S[3]_c_2134_n 0.00416423f $X=11.485 $Y=4.21
+ $X2=0 $Y2=0
cc_1623 N_A_1755_793#_c_1882_n N_S[3]_c_2134_n 0.00289358f $X=11.525 $Y=4.615
+ $X2=0 $Y2=0
cc_1624 N_A_1755_793#_c_1896_n N_S[3]_c_2144_n 0.00929139f $X=11.565 $Y=3.14
+ $X2=0 $Y2=0
cc_1625 N_A_1755_793#_c_1897_n N_S[3]_c_2144_n 0.00117303f $X=11.485 $Y=4.045
+ $X2=0 $Y2=0
cc_1626 N_A_1755_793#_c_1898_n N_S[3]_c_2144_n 0.00304348f $X=11.565 $Y=3.835
+ $X2=0 $Y2=0
cc_1627 N_A_1755_793#_c_1879_n N_S[3]_c_2138_n 0.00426435f $X=11.525 $Y=4.74
+ $X2=0 $Y2=0
cc_1628 N_A_1755_793#_c_1882_n N_S[3]_c_2138_n 0.00268644f $X=11.525 $Y=4.615
+ $X2=0 $Y2=0
cc_1629 N_A_1755_793#_c_1881_n S[3] 0.0228692f $X=11.485 $Y=4.21 $X2=0 $Y2=0
cc_1630 N_A_1755_793#_c_1882_n S[3] 0.00541767f $X=11.525 $Y=4.615 $X2=0 $Y2=0
cc_1631 N_A_1755_793#_c_1884_n N_VPWR_c_3600_n 0.00324472f $X=8.875 $Y=3.965
+ $X2=0 $Y2=0
cc_1632 N_A_1755_793#_c_1891_n N_VPWR_c_3602_n 0.00367058f $X=10.285 $Y=3.965
+ $X2=0 $Y2=0
cc_1633 N_A_1755_793#_c_1877_n N_VPWR_c_3602_n 0.0193185f $X=11.4 $Y=4.21 $X2=0
+ $Y2=0
cc_1634 N_A_1755_793#_c_1878_n N_VPWR_c_3602_n 6.4101e-19 $X=10.855 $Y=4.21
+ $X2=0 $Y2=0
cc_1635 N_A_1755_793#_c_1896_n N_VPWR_c_3602_n 0.0316788f $X=11.565 $Y=3.14
+ $X2=0 $Y2=0
cc_1636 N_A_1755_793#_c_1896_n N_VPWR_c_3604_n 0.0356181f $X=11.565 $Y=3.14
+ $X2=0 $Y2=0
cc_1637 N_A_1755_793#_c_1896_n N_VPWR_c_3632_n 0.0233824f $X=11.565 $Y=3.14
+ $X2=0 $Y2=0
cc_1638 N_A_1755_793#_c_1884_n N_VPWR_c_3661_n 0.00473731f $X=8.875 $Y=3.965
+ $X2=0 $Y2=0
cc_1639 N_A_1755_793#_c_1887_n N_VPWR_c_3661_n 0.00362156f $X=9.345 $Y=3.965
+ $X2=0 $Y2=0
cc_1640 N_A_1755_793#_c_1889_n N_VPWR_c_3661_n 0.00362156f $X=9.815 $Y=3.965
+ $X2=0 $Y2=0
cc_1641 N_A_1755_793#_c_1891_n N_VPWR_c_3661_n 0.00473731f $X=10.285 $Y=3.965
+ $X2=0 $Y2=0
cc_1642 N_A_1755_793#_c_1896_n N_VPWR_c_3661_n 0.00593513f $X=11.565 $Y=3.14
+ $X2=0 $Y2=0
cc_1643 N_A_1755_793#_c_1888_n N_Z_c_4595_n 0.00762343f $X=9.725 $Y=4.04 $X2=0
+ $Y2=0
cc_1644 N_A_1755_793#_c_1892_n N_Z_c_4595_n 0.00704092f $X=9.345 $Y=4.04 $X2=0
+ $Y2=0
cc_1645 N_A_1755_793#_c_1886_n N_Z_c_4616_n 0.00248496f $X=8.965 $Y=4.04 $X2=0
+ $Y2=0
cc_1646 N_A_1755_793#_c_1885_n N_Z_c_4619_n 0.00678861f $X=9.255 $Y=4.04 $X2=0
+ $Y2=0
cc_1647 N_A_1755_793#_c_1886_n N_Z_c_4619_n 0.00239476f $X=8.965 $Y=4.04 $X2=0
+ $Y2=0
cc_1648 N_A_1755_793#_c_1892_n N_Z_c_4619_n 2.98555e-19 $X=9.345 $Y=4.04 $X2=0
+ $Y2=0
cc_1649 N_A_1755_793#_c_1888_n N_Z_c_4621_n 0.00145542f $X=9.725 $Y=4.04 $X2=0
+ $Y2=0
cc_1650 N_A_1755_793#_c_1890_n N_Z_c_4621_n 0.00597584f $X=10.195 $Y=4.04 $X2=0
+ $Y2=0
cc_1651 N_A_1755_793#_c_1893_n N_Z_c_4621_n 0.00909323f $X=9.815 $Y=4.04 $X2=0
+ $Y2=0
cc_1652 N_A_1755_793#_c_1877_n N_Z_c_4621_n 0.0266078f $X=11.4 $Y=4.21 $X2=0
+ $Y2=0
cc_1653 N_A_1755_793#_c_1883_n N_Z_c_4621_n 0.00747617f $X=10.605 $Y=4.21 $X2=0
+ $Y2=0
cc_1654 N_A_1755_793#_c_1884_n N_Z_c_4645_n 0.00834829f $X=8.875 $Y=3.965 $X2=0
+ $Y2=0
cc_1655 N_A_1755_793#_c_1891_n N_Z_c_4647_n 0.00795576f $X=10.285 $Y=3.965 $X2=0
+ $Y2=0
cc_1656 N_A_1755_793#_c_1877_n N_Z_c_4647_n 0.0186685f $X=11.4 $Y=4.21 $X2=0
+ $Y2=0
cc_1657 N_A_1755_793#_c_1896_n N_Z_c_4647_n 0.0329704f $X=11.565 $Y=3.14 $X2=0
+ $Y2=0
cc_1658 N_A_1755_793#_c_1883_n N_Z_c_4647_n 2.19754e-19 $X=10.605 $Y=4.21 $X2=0
+ $Y2=0
cc_1659 N_A_1755_793#_c_1887_n Z 0.00372458f $X=9.345 $Y=3.965 $X2=0 $Y2=0
cc_1660 N_A_1755_793#_c_1889_n Z 0.00372248f $X=9.815 $Y=3.965 $X2=0 $Y2=0
cc_1661 N_A_1755_793#_c_1884_n N_Z_c_4652_n 0.0199111f $X=8.875 $Y=3.965 $X2=0
+ $Y2=0
cc_1662 N_A_1755_793#_c_1885_n N_Z_c_4652_n 0.00560592f $X=9.255 $Y=4.04 $X2=0
+ $Y2=0
cc_1663 N_A_1755_793#_c_1886_n N_Z_c_4652_n 0.00474497f $X=8.965 $Y=4.04 $X2=0
+ $Y2=0
cc_1664 N_A_1755_793#_c_1887_n N_Z_c_4652_n 0.0181262f $X=9.345 $Y=3.965 $X2=0
+ $Y2=0
cc_1665 N_A_1755_793#_c_1889_n N_Z_c_4652_n 9.74366e-19 $X=9.815 $Y=3.965 $X2=0
+ $Y2=0
cc_1666 N_A_1755_793#_c_1892_n N_Z_c_4652_n 0.00415268f $X=9.345 $Y=4.04 $X2=0
+ $Y2=0
cc_1667 N_A_1755_793#_c_1887_n N_Z_c_4653_n 9.74366e-19 $X=9.345 $Y=3.965 $X2=0
+ $Y2=0
cc_1668 N_A_1755_793#_c_1889_n N_Z_c_4653_n 0.0181262f $X=9.815 $Y=3.965 $X2=0
+ $Y2=0
cc_1669 N_A_1755_793#_c_1890_n N_Z_c_4653_n 0.00560592f $X=10.195 $Y=4.04 $X2=0
+ $Y2=0
cc_1670 N_A_1755_793#_c_1891_n N_Z_c_4653_n 0.0221748f $X=10.285 $Y=3.965 $X2=0
+ $Y2=0
cc_1671 N_A_1755_793#_c_1893_n N_Z_c_4653_n 0.00181273f $X=9.815 $Y=4.04 $X2=0
+ $Y2=0
cc_1672 N_A_1755_793#_c_1877_n N_Z_c_4653_n 0.00240108f $X=11.4 $Y=4.21 $X2=0
+ $Y2=0
cc_1673 N_A_1755_793#_c_1883_n N_Z_c_4653_n 0.00425035f $X=10.605 $Y=4.21 $X2=0
+ $Y2=0
cc_1674 N_A_1755_793#_c_1884_n N_A_1313_591#_c_5630_n 0.00151141f $X=8.875
+ $Y=3.965 $X2=0 $Y2=0
cc_1675 N_A_1755_793#_c_1884_n N_A_1313_591#_c_5659_n 0.00307958f $X=8.875
+ $Y=3.965 $X2=0 $Y2=0
cc_1676 N_A_1755_793#_c_1887_n N_A_1313_591#_c_5659_n 0.00307958f $X=9.345
+ $Y=3.965 $X2=0 $Y2=0
cc_1677 N_A_1755_793#_c_1889_n N_A_1313_591#_c_5661_n 0.00307958f $X=9.815
+ $Y=3.965 $X2=0 $Y2=0
cc_1678 N_A_1755_793#_c_1891_n N_A_1313_591#_c_5661_n 0.00307958f $X=10.285
+ $Y=3.965 $X2=0 $Y2=0
cc_1679 N_A_1755_793#_c_1884_n N_A_1313_591#_c_5632_n 0.00554566f $X=8.875
+ $Y=3.965 $X2=0 $Y2=0
cc_1680 N_A_1755_793#_c_1887_n N_A_1313_591#_c_5633_n 0.00210632f $X=9.345
+ $Y=3.965 $X2=0 $Y2=0
cc_1681 N_A_1755_793#_c_1888_n N_A_1313_591#_c_5633_n 0.00251792f $X=9.725
+ $Y=4.04 $X2=0 $Y2=0
cc_1682 N_A_1755_793#_c_1889_n N_A_1313_591#_c_5633_n 0.00210632f $X=9.815
+ $Y=3.965 $X2=0 $Y2=0
cc_1683 N_A_1755_793#_c_1891_n N_A_1313_591#_c_5634_n 0.00499839f $X=10.285
+ $Y=3.965 $X2=0 $Y2=0
cc_1684 N_A_1755_793#_c_1877_n N_A_1313_591#_c_5634_n 0.0218124f $X=11.4 $Y=4.21
+ $X2=0 $Y2=0
cc_1685 N_A_1755_793#_c_1878_n N_A_1313_591#_c_5634_n 5.74251e-19 $X=10.855
+ $Y=4.21 $X2=0 $Y2=0
cc_1686 N_A_1755_793#_c_1883_n N_A_1313_591#_c_5634_n 0.00561627f $X=10.605
+ $Y=4.21 $X2=0 $Y2=0
cc_1687 N_A_1755_793#_c_1877_n N_VGND_c_6283_n 0.0123065f $X=11.4 $Y=4.21 $X2=0
+ $Y2=0
cc_1688 N_A_1755_793#_c_1878_n N_VGND_c_6283_n 2.04129e-19 $X=10.855 $Y=4.21
+ $X2=0 $Y2=0
cc_1689 N_A_1755_793#_c_1880_n N_VGND_c_6322_n 0.0129994f $X=11.565 $Y=4.995
+ $X2=0 $Y2=0
cc_1690 N_A_1755_793#_M1060_s N_VGND_c_6371_n 0.00394793f $X=11.43 $Y=4.785
+ $X2=0 $Y2=0
cc_1691 N_A_1755_793#_c_1880_n N_VGND_c_6371_n 0.00927134f $X=11.565 $Y=4.995
+ $X2=0 $Y2=0
cc_1692 N_A_1755_793#_c_1892_n N_A_1315_911#_c_7199_n 7.0477e-19 $X=9.345
+ $Y=4.04 $X2=0 $Y2=0
cc_1693 N_A_1755_793#_c_1877_n N_A_1315_911#_c_7180_n 0.0028695f $X=11.4 $Y=4.21
+ $X2=0 $Y2=0
cc_1694 N_A_1755_793#_c_1883_n N_A_1315_911#_c_7180_n 0.00589316f $X=10.605
+ $Y=4.21 $X2=0 $Y2=0
cc_1695 N_S[2]_c_2025_n N_S[3]_c_2142_n 0.0130744f $X=11.33 $Y=1.55 $X2=0 $Y2=0
cc_1696 N_S[2]_c_2018_n N_S[3]_c_2144_n 0.0130744f $X=11.8 $Y=1.55 $X2=0 $Y2=0
cc_1697 N_S[2]_c_2018_n N_S[4]_c_2244_n 0.0215827f $X=11.8 $Y=1.55 $X2=-0.19
+ $Y2=-0.24
cc_1698 S[2] N_S[4]_c_2244_n 0.00113563f $X=12.105 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_1699 N_S[2]_c_2018_n N_S[4]_c_2265_n 0.00113563f $X=11.8 $Y=1.55 $X2=0 $Y2=0
cc_1700 S[2] N_S[4]_c_2265_n 0.0301108f $X=12.105 $Y=1.105 $X2=0 $Y2=0
cc_1701 N_S[2]_c_2025_n N_VPWR_c_3601_n 0.00950399f $X=11.33 $Y=1.55 $X2=0 $Y2=0
cc_1702 N_S[2]_c_2018_n N_VPWR_c_3603_n 0.016386f $X=11.8 $Y=1.55 $X2=0 $Y2=0
cc_1703 S[2] N_VPWR_c_3603_n 0.0157609f $X=12.105 $Y=1.105 $X2=0 $Y2=0
cc_1704 N_S[2]_c_2025_n N_VPWR_c_3632_n 0.0035837f $X=11.33 $Y=1.55 $X2=0 $Y2=0
cc_1705 N_S[2]_c_2018_n N_VPWR_c_3632_n 0.0035837f $X=11.8 $Y=1.55 $X2=0 $Y2=0
cc_1706 N_S[2]_c_2025_n N_VPWR_c_3661_n 0.00711603f $X=11.33 $Y=1.55 $X2=0 $Y2=0
cc_1707 N_S[2]_c_2018_n N_VPWR_c_3661_n 0.0070533f $X=11.8 $Y=1.55 $X2=0 $Y2=0
cc_1708 N_S[2]_c_2002_n N_Z_c_4593_n 0.002324f $X=8.8 $Y=0.255 $X2=0 $Y2=0
cc_1709 N_S[2]_c_2005_n N_Z_c_4593_n 0.00283489f $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_1710 N_S[2]_c_2005_n N_Z_c_4594_n 3.10191e-19 $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_1711 N_S[2]_c_2007_n N_Z_c_4594_n 0.00190704f $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_1712 N_S[2]_c_2005_n N_Z_c_4596_n 6.35774e-19 $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_1713 N_S[2]_c_2007_n N_Z_c_4596_n 0.0077801f $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_1714 N_S[2]_c_2009_n N_Z_c_4596_n 0.0134253f $X=10.06 $Y=0.255 $X2=0 $Y2=0
cc_1715 N_S[2]_c_2002_n N_Z_c_4615_n 0.00443615f $X=8.8 $Y=0.255 $X2=0 $Y2=0
cc_1716 N_S[2]_c_2005_n N_Z_c_4615_n 0.00462308f $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_1717 N_S[2]_c_2007_n N_Z_c_4615_n 6.35664e-19 $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_1718 N_S[2]_c_2005_n N_Z_c_4618_n 0.00180363f $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_1719 N_S[2]_c_2009_n N_Z_c_4620_n 0.00216436f $X=10.06 $Y=0.255 $X2=0 $Y2=0
cc_1720 N_S[2]_c_2025_n N_Z_c_4646_n 0.00478771f $X=11.33 $Y=1.55 $X2=0 $Y2=0
cc_1721 N_S[2]_c_2018_n N_Z_c_4646_n 0.00760321f $X=11.8 $Y=1.55 $X2=0 $Y2=0
cc_1722 S[2] N_Z_c_4646_n 0.010609f $X=12.105 $Y=1.105 $X2=0 $Y2=0
cc_1723 N_S[2]_c_2002_n N_A_1313_297#_c_5502_n 0.00168571f $X=8.8 $Y=0.255 $X2=0
+ $Y2=0
cc_1724 N_S[2]_c_2025_n N_A_1313_297#_c_5506_n 0.00239129f $X=11.33 $Y=1.55
+ $X2=0 $Y2=0
cc_1725 N_S[2]_c_2002_n N_VGND_c_6280_n 5.5039e-19 $X=8.8 $Y=0.255 $X2=0 $Y2=0
cc_1726 N_S[2]_c_2004_n N_VGND_c_6280_n 0.0028166f $X=8.875 $Y=0.18 $X2=0 $Y2=0
cc_1727 N_S[2]_c_2010_n N_VGND_c_6282_n 0.00862298f $X=10.745 $Y=0.18 $X2=0
+ $Y2=0
cc_1728 N_S[2]_c_2012_n N_VGND_c_6282_n 0.00525833f $X=11.23 $Y=0.81 $X2=0 $Y2=0
cc_1729 N_S[2]_c_2015_n N_VGND_c_6282_n 0.00173127f $X=11.355 $Y=0.735 $X2=0
+ $Y2=0
cc_1730 N_S[2]_c_2017_n N_VGND_c_6284_n 0.00374526f $X=11.775 $Y=0.735 $X2=0
+ $Y2=0
cc_1731 N_S[2]_c_2018_n N_VGND_c_6284_n 0.00578076f $X=11.8 $Y=1.55 $X2=0 $Y2=0
cc_1732 S[2] N_VGND_c_6284_n 0.0116413f $X=12.105 $Y=1.105 $X2=0 $Y2=0
cc_1733 N_S[2]_c_2004_n N_VGND_c_6316_n 0.0559651f $X=8.875 $Y=0.18 $X2=0 $Y2=0
cc_1734 N_S[2]_c_2015_n N_VGND_c_6320_n 0.00542362f $X=11.355 $Y=0.735 $X2=0
+ $Y2=0
cc_1735 N_S[2]_c_2016_n N_VGND_c_6320_n 2.16067e-19 $X=11.7 $Y=0.81 $X2=0 $Y2=0
cc_1736 N_S[2]_c_2017_n N_VGND_c_6320_n 0.00585385f $X=11.775 $Y=0.735 $X2=0
+ $Y2=0
cc_1737 N_S[2]_c_2003_n N_VGND_c_6370_n 0.00642387f $X=9.145 $Y=0.18 $X2=0 $Y2=0
cc_1738 N_S[2]_c_2004_n N_VGND_c_6370_n 0.00591981f $X=8.875 $Y=0.18 $X2=0 $Y2=0
cc_1739 N_S[2]_c_2006_n N_VGND_c_6370_n 0.0064237f $X=9.565 $Y=0.18 $X2=0 $Y2=0
cc_1740 N_S[2]_c_2008_n N_VGND_c_6370_n 0.00642387f $X=9.985 $Y=0.18 $X2=0 $Y2=0
cc_1741 N_S[2]_c_2010_n N_VGND_c_6370_n 0.0345801f $X=10.745 $Y=0.18 $X2=0 $Y2=0
cc_1742 N_S[2]_c_2015_n N_VGND_c_6370_n 0.00990284f $X=11.355 $Y=0.735 $X2=0
+ $Y2=0
cc_1743 N_S[2]_c_2017_n N_VGND_c_6370_n 0.0119653f $X=11.775 $Y=0.735 $X2=0
+ $Y2=0
cc_1744 N_S[2]_c_2019_n N_VGND_c_6370_n 0.00366655f $X=9.22 $Y=0.18 $X2=0 $Y2=0
cc_1745 N_S[2]_c_2020_n N_VGND_c_6370_n 0.00366655f $X=9.64 $Y=0.18 $X2=0 $Y2=0
cc_1746 N_S[2]_c_2021_n N_VGND_c_6370_n 0.00366655f $X=10.06 $Y=0.18 $X2=0 $Y2=0
cc_1747 N_S[2]_c_2002_n N_A_1315_47#_c_7093_n 0.00206084f $X=8.8 $Y=0.255 $X2=0
+ $Y2=0
cc_1748 N_S[2]_c_2002_n N_A_1315_47#_c_7095_n 0.0139014f $X=8.8 $Y=0.255 $X2=0
+ $Y2=0
cc_1749 N_S[2]_c_2003_n N_A_1315_47#_c_7095_n 0.00211351f $X=9.145 $Y=0.18 $X2=0
+ $Y2=0
cc_1750 N_S[2]_c_2005_n N_A_1315_47#_c_7095_n 0.0106826f $X=9.22 $Y=0.255 $X2=0
+ $Y2=0
cc_1751 N_S[2]_c_2007_n N_A_1315_47#_c_7097_n 0.0106844f $X=9.64 $Y=0.255 $X2=0
+ $Y2=0
cc_1752 N_S[2]_c_2008_n N_A_1315_47#_c_7097_n 0.00211351f $X=9.985 $Y=0.18 $X2=0
+ $Y2=0
cc_1753 N_S[2]_c_2009_n N_A_1315_47#_c_7097_n 0.0112916f $X=10.06 $Y=0.255 $X2=0
+ $Y2=0
cc_1754 N_S[2]_c_2010_n N_A_1315_47#_c_7097_n 0.00685838f $X=10.745 $Y=0.18
+ $X2=0 $Y2=0
cc_1755 N_S[2]_c_2011_n N_A_1315_47#_c_7097_n 0.00189496f $X=10.82 $Y=0.735
+ $X2=0 $Y2=0
cc_1756 N_S[2]_c_2011_n N_A_1315_47#_c_7098_n 0.00529837f $X=10.82 $Y=0.735
+ $X2=0 $Y2=0
cc_1757 N_S[2]_c_2006_n N_A_1315_47#_c_7133_n 0.0034777f $X=9.565 $Y=0.18 $X2=0
+ $Y2=0
cc_1758 N_S[3]_c_2134_n N_S[5]_c_2364_n 0.0215827f $X=11.775 $Y=4.705 $X2=-0.19
+ $Y2=-0.24
cc_1759 S[3] N_S[5]_c_2364_n 0.00113563f $X=12.105 $Y=4.165 $X2=-0.19 $Y2=-0.24
cc_1760 N_S[3]_c_2134_n N_S[5]_c_2384_n 0.00113563f $X=11.775 $Y=4.705 $X2=0
+ $Y2=0
cc_1761 S[3] N_S[5]_c_2384_n 0.0301108f $X=12.105 $Y=4.165 $X2=0 $Y2=0
cc_1762 N_S[3]_c_2142_n N_VPWR_c_3602_n 0.00950399f $X=11.33 $Y=3.89 $X2=0 $Y2=0
cc_1763 N_S[3]_c_2134_n N_VPWR_c_3604_n 0.00652399f $X=11.775 $Y=4.705 $X2=0
+ $Y2=0
cc_1764 N_S[3]_c_2144_n N_VPWR_c_3604_n 0.00986205f $X=11.8 $Y=3.89 $X2=0 $Y2=0
cc_1765 S[3] N_VPWR_c_3604_n 0.0157609f $X=12.105 $Y=4.165 $X2=0 $Y2=0
cc_1766 N_S[3]_c_2142_n N_VPWR_c_3632_n 0.0035837f $X=11.33 $Y=3.89 $X2=0 $Y2=0
cc_1767 N_S[3]_c_2144_n N_VPWR_c_3632_n 0.0035837f $X=11.8 $Y=3.89 $X2=0 $Y2=0
cc_1768 N_S[3]_c_2142_n N_VPWR_c_3661_n 0.00711603f $X=11.33 $Y=3.89 $X2=0 $Y2=0
cc_1769 N_S[3]_c_2144_n N_VPWR_c_3661_n 0.0070533f $X=11.8 $Y=3.89 $X2=0 $Y2=0
cc_1770 N_S[3]_c_2122_n N_Z_c_4595_n 3.10191e-19 $X=9.22 $Y=5.185 $X2=0 $Y2=0
cc_1771 N_S[3]_c_2124_n N_Z_c_4595_n 0.00190704f $X=9.64 $Y=5.185 $X2=0 $Y2=0
cc_1772 N_S[3]_c_2122_n N_Z_c_4597_n 6.35774e-19 $X=9.22 $Y=5.185 $X2=0 $Y2=0
cc_1773 N_S[3]_c_2124_n N_Z_c_4597_n 0.0077801f $X=9.64 $Y=5.185 $X2=0 $Y2=0
cc_1774 N_S[3]_c_2126_n N_Z_c_4597_n 0.0134253f $X=10.06 $Y=5.185 $X2=0 $Y2=0
cc_1775 N_S[3]_c_2119_n N_Z_c_4616_n 0.00443615f $X=8.8 $Y=5.185 $X2=0 $Y2=0
cc_1776 N_S[3]_c_2122_n N_Z_c_4616_n 0.00462308f $X=9.22 $Y=5.185 $X2=0 $Y2=0
cc_1777 N_S[3]_c_2119_n N_Z_c_4617_n 0.002324f $X=8.8 $Y=5.185 $X2=0 $Y2=0
cc_1778 N_S[3]_c_2122_n N_Z_c_4617_n 0.00283489f $X=9.22 $Y=5.185 $X2=0 $Y2=0
cc_1779 N_S[3]_c_2124_n N_Z_c_4617_n 6.35664e-19 $X=9.64 $Y=5.185 $X2=0 $Y2=0
cc_1780 N_S[3]_c_2122_n N_Z_c_4619_n 0.00180363f $X=9.22 $Y=5.185 $X2=0 $Y2=0
cc_1781 N_S[3]_c_2126_n N_Z_c_4621_n 0.00216436f $X=10.06 $Y=5.185 $X2=0 $Y2=0
cc_1782 N_S[3]_c_2140_n N_Z_c_4647_n 2.55735e-19 $X=11.33 $Y=3.99 $X2=0 $Y2=0
cc_1783 N_S[3]_c_2142_n N_Z_c_4647_n 0.00453198f $X=11.33 $Y=3.89 $X2=0 $Y2=0
cc_1784 N_S[3]_c_2134_n N_Z_c_4647_n 0.00258545f $X=11.775 $Y=4.705 $X2=0 $Y2=0
cc_1785 N_S[3]_c_2144_n N_Z_c_4647_n 0.00501777f $X=11.8 $Y=3.89 $X2=0 $Y2=0
cc_1786 S[3] N_Z_c_4647_n 0.010609f $X=12.105 $Y=4.165 $X2=0 $Y2=0
cc_1787 N_S[3]_c_2119_n N_A_1313_591#_c_5630_n 0.00168571f $X=8.8 $Y=5.185 $X2=0
+ $Y2=0
cc_1788 N_S[3]_c_2142_n N_A_1313_591#_c_5634_n 0.00239129f $X=11.33 $Y=3.89
+ $X2=0 $Y2=0
cc_1789 N_S[3]_c_2119_n N_VGND_c_6281_n 5.5039e-19 $X=8.8 $Y=5.185 $X2=0 $Y2=0
cc_1790 N_S[3]_c_2121_n N_VGND_c_6281_n 0.0028166f $X=8.875 $Y=5.26 $X2=0 $Y2=0
cc_1791 N_S[3]_c_2128_n N_VGND_c_6283_n 0.00862298f $X=10.82 $Y=5.185 $X2=0
+ $Y2=0
cc_1792 N_S[3]_c_2129_n N_VGND_c_6283_n 0.00525833f $X=11.23 $Y=4.63 $X2=0 $Y2=0
cc_1793 N_S[3]_c_2132_n N_VGND_c_6283_n 0.00173127f $X=11.355 $Y=4.705 $X2=0
+ $Y2=0
cc_1794 N_S[3]_c_2134_n N_VGND_c_6285_n 0.00952602f $X=11.775 $Y=4.705 $X2=0
+ $Y2=0
cc_1795 S[3] N_VGND_c_6285_n 0.0116413f $X=12.105 $Y=4.165 $X2=0 $Y2=0
cc_1796 N_S[3]_c_2121_n N_VGND_c_6318_n 0.0559651f $X=8.875 $Y=5.26 $X2=0 $Y2=0
cc_1797 N_S[3]_c_2132_n N_VGND_c_6322_n 0.00542362f $X=11.355 $Y=4.705 $X2=0
+ $Y2=0
cc_1798 N_S[3]_c_2133_n N_VGND_c_6322_n 2.16067e-19 $X=11.7 $Y=4.63 $X2=0 $Y2=0
cc_1799 N_S[3]_c_2134_n N_VGND_c_6322_n 0.00585385f $X=11.775 $Y=4.705 $X2=0
+ $Y2=0
cc_1800 N_S[3]_c_2120_n N_VGND_c_6371_n 0.00642387f $X=9.145 $Y=5.26 $X2=0 $Y2=0
cc_1801 N_S[3]_c_2121_n N_VGND_c_6371_n 0.00591981f $X=8.875 $Y=5.26 $X2=0 $Y2=0
cc_1802 N_S[3]_c_2123_n N_VGND_c_6371_n 0.0064237f $X=9.565 $Y=5.26 $X2=0 $Y2=0
cc_1803 N_S[3]_c_2125_n N_VGND_c_6371_n 0.00642387f $X=9.985 $Y=5.26 $X2=0 $Y2=0
cc_1804 N_S[3]_c_2127_n N_VGND_c_6371_n 0.0345801f $X=10.745 $Y=5.26 $X2=0 $Y2=0
cc_1805 N_S[3]_c_2132_n N_VGND_c_6371_n 0.00990284f $X=11.355 $Y=4.705 $X2=0
+ $Y2=0
cc_1806 N_S[3]_c_2134_n N_VGND_c_6371_n 0.0119653f $X=11.775 $Y=4.705 $X2=0
+ $Y2=0
cc_1807 N_S[3]_c_2135_n N_VGND_c_6371_n 0.00366655f $X=9.22 $Y=5.26 $X2=0 $Y2=0
cc_1808 N_S[3]_c_2136_n N_VGND_c_6371_n 0.00366655f $X=9.64 $Y=5.26 $X2=0 $Y2=0
cc_1809 N_S[3]_c_2137_n N_VGND_c_6371_n 0.00366655f $X=10.06 $Y=5.26 $X2=0 $Y2=0
cc_1810 N_S[3]_c_2119_n N_A_1315_911#_c_7175_n 0.00206084f $X=8.8 $Y=5.185 $X2=0
+ $Y2=0
cc_1811 N_S[3]_c_2119_n N_A_1315_911#_c_7177_n 0.0139014f $X=8.8 $Y=5.185 $X2=0
+ $Y2=0
cc_1812 N_S[3]_c_2120_n N_A_1315_911#_c_7177_n 0.00211351f $X=9.145 $Y=5.26
+ $X2=0 $Y2=0
cc_1813 N_S[3]_c_2122_n N_A_1315_911#_c_7177_n 0.0106826f $X=9.22 $Y=5.185 $X2=0
+ $Y2=0
cc_1814 N_S[3]_c_2124_n N_A_1315_911#_c_7179_n 0.0106844f $X=9.64 $Y=5.185 $X2=0
+ $Y2=0
cc_1815 N_S[3]_c_2125_n N_A_1315_911#_c_7179_n 0.00211351f $X=9.985 $Y=5.26
+ $X2=0 $Y2=0
cc_1816 N_S[3]_c_2126_n N_A_1315_911#_c_7179_n 0.0112916f $X=10.06 $Y=5.185
+ $X2=0 $Y2=0
cc_1817 N_S[3]_c_2127_n N_A_1315_911#_c_7179_n 0.00685838f $X=10.745 $Y=5.26
+ $X2=0 $Y2=0
cc_1818 N_S[3]_c_2128_n N_A_1315_911#_c_7179_n 0.00189496f $X=10.82 $Y=5.185
+ $X2=0 $Y2=0
cc_1819 N_S[3]_c_2130_n N_A_1315_911#_c_7180_n 0.00529837f $X=10.895 $Y=4.63
+ $X2=0 $Y2=0
cc_1820 N_S[3]_c_2123_n N_A_1315_911#_c_7212_n 0.0034777f $X=9.565 $Y=5.26 $X2=0
+ $Y2=0
cc_1821 N_S[4]_c_2245_n N_S[5]_c_2386_n 0.0130744f $X=13.04 $Y=1.55 $X2=0 $Y2=0
cc_1822 N_S[4]_c_2269_n N_S[5]_c_2390_n 0.0130744f $X=13.51 $Y=1.55 $X2=0 $Y2=0
cc_1823 N_S[4]_c_2254_n N_A_2626_325#_c_2500_n 0.00507688f $X=14.78 $Y=0.255
+ $X2=0 $Y2=0
cc_1824 N_S[4]_c_2249_n N_A_2626_325#_c_2492_n 0.00262132f $X=13.51 $Y=1.45
+ $X2=0 $Y2=0
cc_1825 N_S[4]_c_2256_n N_A_2626_325#_c_2503_n 0.00509204f $X=15.2 $Y=0.255
+ $X2=0 $Y2=0
cc_1826 N_S[4]_c_2260_n N_A_2626_325#_c_2505_n 0.00507426f $X=16.04 $Y=0.255
+ $X2=0 $Y2=0
cc_1827 N_S[4]_c_2258_n N_A_2626_325#_c_2508_n 0.00509391f $X=15.62 $Y=0.255
+ $X2=0 $Y2=0
cc_1828 N_S[4]_c_2245_n N_A_2626_325#_c_2509_n 0.0128834f $X=13.04 $Y=1.55 $X2=0
+ $Y2=0
cc_1829 N_S[4]_c_2269_n N_A_2626_325#_c_2509_n 0.0118698f $X=13.51 $Y=1.55 $X2=0
+ $Y2=0
cc_1830 N_S[4]_c_2246_n N_A_2626_325#_c_2493_n 0.00207203f $X=13.065 $Y=0.735
+ $X2=0 $Y2=0
cc_1831 N_S[4]_c_2248_n N_A_2626_325#_c_2493_n 0.00603996f $X=13.485 $Y=0.735
+ $X2=0 $Y2=0
cc_1832 N_S[4]_c_2251_n N_A_2626_325#_c_2493_n 6.53442e-19 $X=14.02 $Y=0.735
+ $X2=0 $Y2=0
cc_1833 N_S[4]_c_2245_n N_A_2626_325#_c_2494_n 0.00289358f $X=13.04 $Y=1.55
+ $X2=0 $Y2=0
cc_1834 N_S[4]_c_2247_n N_A_2626_325#_c_2494_n 0.00429801f $X=13.41 $Y=0.81
+ $X2=0 $Y2=0
cc_1835 N_S[4]_c_2249_n N_A_2626_325#_c_2494_n 0.0085951f $X=13.51 $Y=1.45 $X2=0
+ $Y2=0
cc_1836 N_S[4]_c_2261_n N_A_2626_325#_c_2494_n 0.00268644f $X=13.51 $Y=0.81
+ $X2=0 $Y2=0
cc_1837 N_S[4]_c_2265_n N_A_2626_325#_c_2494_n 0.00541767f $X=13 $Y=1.16 $X2=0
+ $Y2=0
cc_1838 N_S[4]_c_2249_n N_A_2626_325#_c_2495_n 0.0206368f $X=13.51 $Y=1.45 $X2=0
+ $Y2=0
cc_1839 N_S[4]_c_2250_n N_A_2626_325#_c_2495_n 0.0103812f $X=13.945 $Y=0.81
+ $X2=0 $Y2=0
cc_1840 N_S[4]_c_2245_n N_A_2626_325#_c_2511_n 0.00454075f $X=13.04 $Y=1.55
+ $X2=0 $Y2=0
cc_1841 N_S[4]_c_2249_n N_A_2626_325#_c_2511_n 0.00255921f $X=13.51 $Y=1.45
+ $X2=0 $Y2=0
cc_1842 N_S[4]_c_2269_n N_A_2626_325#_c_2511_n 0.00762115f $X=13.51 $Y=1.55
+ $X2=0 $Y2=0
cc_1843 N_S[4]_c_2247_n N_A_2626_325#_c_2496_n 0.0111895f $X=13.41 $Y=0.81 $X2=0
+ $Y2=0
cc_1844 N_S[4]_c_2248_n N_A_2626_325#_c_2496_n 9.67113e-19 $X=13.485 $Y=0.735
+ $X2=0 $Y2=0
cc_1845 N_S[4]_c_2261_n N_A_2626_325#_c_2496_n 0.00426435f $X=13.51 $Y=0.81
+ $X2=0 $Y2=0
cc_1846 N_S[4]_c_2245_n N_A_2626_325#_c_2497_n 0.00416423f $X=13.04 $Y=1.55
+ $X2=0 $Y2=0
cc_1847 N_S[4]_c_2249_n N_A_2626_325#_c_2497_n 0.00322131f $X=13.51 $Y=1.45
+ $X2=0 $Y2=0
cc_1848 N_S[4]_c_2265_n N_A_2626_325#_c_2497_n 0.0228692f $X=13 $Y=1.16 $X2=0
+ $Y2=0
cc_1849 N_S[4]_c_2249_n N_A_2626_325#_c_2498_n 0.0175393f $X=13.51 $Y=1.45 $X2=0
+ $Y2=0
cc_1850 N_S[4]_c_2250_n N_A_2626_325#_c_2498_n 0.0179529f $X=13.945 $Y=0.81
+ $X2=0 $Y2=0
cc_1851 N_S[4]_c_2244_n N_VPWR_c_3606_n 0.00652399f $X=12.94 $Y=1.16 $X2=0 $Y2=0
cc_1852 N_S[4]_c_2245_n N_VPWR_c_3606_n 0.00986205f $X=13.04 $Y=1.55 $X2=0 $Y2=0
cc_1853 N_S[4]_c_2265_n N_VPWR_c_3606_n 0.0157609f $X=13 $Y=1.16 $X2=0 $Y2=0
cc_1854 N_S[4]_c_2269_n N_VPWR_c_3608_n 0.00950399f $X=13.51 $Y=1.55 $X2=0 $Y2=0
cc_1855 N_S[4]_c_2245_n N_VPWR_c_3635_n 0.0035837f $X=13.04 $Y=1.55 $X2=0 $Y2=0
cc_1856 N_S[4]_c_2269_n N_VPWR_c_3635_n 0.0035837f $X=13.51 $Y=1.55 $X2=0 $Y2=0
cc_1857 N_S[4]_c_2245_n N_VPWR_c_3661_n 0.0070533f $X=13.04 $Y=1.55 $X2=0 $Y2=0
cc_1858 N_S[4]_c_2269_n N_VPWR_c_3661_n 0.00711603f $X=13.51 $Y=1.55 $X2=0 $Y2=0
cc_1859 N_S[4]_c_2254_n N_Z_c_4598_n 0.0134253f $X=14.78 $Y=0.255 $X2=0 $Y2=0
cc_1860 N_S[4]_c_2256_n N_Z_c_4598_n 0.0077801f $X=15.2 $Y=0.255 $X2=0 $Y2=0
cc_1861 N_S[4]_c_2258_n N_Z_c_4598_n 6.35774e-19 $X=15.62 $Y=0.255 $X2=0 $Y2=0
cc_1862 N_S[4]_c_2256_n N_Z_c_4600_n 0.00190704f $X=15.2 $Y=0.255 $X2=0 $Y2=0
cc_1863 N_S[4]_c_2258_n N_Z_c_4600_n 3.10191e-19 $X=15.62 $Y=0.255 $X2=0 $Y2=0
cc_1864 N_S[4]_c_2258_n N_Z_c_4602_n 0.00283489f $X=15.62 $Y=0.255 $X2=0 $Y2=0
cc_1865 N_S[4]_c_2260_n N_Z_c_4602_n 0.002324f $X=16.04 $Y=0.255 $X2=0 $Y2=0
cc_1866 N_S[4]_c_2254_n N_Z_c_4622_n 0.00216436f $X=14.78 $Y=0.255 $X2=0 $Y2=0
cc_1867 N_S[4]_c_2258_n N_Z_c_4624_n 0.00180363f $X=15.62 $Y=0.255 $X2=0 $Y2=0
cc_1868 N_S[4]_c_2256_n N_Z_c_4626_n 6.35664e-19 $X=15.2 $Y=0.255 $X2=0 $Y2=0
cc_1869 N_S[4]_c_2258_n N_Z_c_4626_n 0.00462308f $X=15.62 $Y=0.255 $X2=0 $Y2=0
cc_1870 N_S[4]_c_2260_n N_Z_c_4626_n 0.00443615f $X=16.04 $Y=0.255 $X2=0 $Y2=0
cc_1871 N_S[4]_c_2244_n N_Z_c_4646_n 0.00234109f $X=12.94 $Y=1.16 $X2=0 $Y2=0
cc_1872 N_S[4]_c_2245_n N_Z_c_4646_n 0.0052507f $X=13.04 $Y=1.55 $X2=0 $Y2=0
cc_1873 N_S[4]_c_2269_n N_Z_c_4646_n 0.00478771f $X=13.51 $Y=1.55 $X2=0 $Y2=0
cc_1874 N_S[4]_c_2265_n N_Z_c_4646_n 0.0105931f $X=13 $Y=1.16 $X2=0 $Y2=0
cc_1875 N_S[4]_c_2260_n N_A_2839_311#_c_5759_n 0.00168571f $X=16.04 $Y=0.255
+ $X2=0 $Y2=0
cc_1876 N_S[4]_c_2269_n N_A_2839_311#_c_5761_n 0.00239129f $X=13.51 $Y=1.55
+ $X2=0 $Y2=0
cc_1877 N_S[4]_c_2244_n N_VGND_c_6286_n 0.00576464f $X=12.94 $Y=1.16 $X2=0 $Y2=0
cc_1878 N_S[4]_c_2246_n N_VGND_c_6286_n 0.00374526f $X=13.065 $Y=0.735 $X2=0
+ $Y2=0
cc_1879 N_S[4]_c_2265_n N_VGND_c_6286_n 0.0116218f $X=13 $Y=1.16 $X2=0 $Y2=0
cc_1880 N_S[4]_c_2248_n N_VGND_c_6288_n 0.00173127f $X=13.485 $Y=0.735 $X2=0
+ $Y2=0
cc_1881 N_S[4]_c_2250_n N_VGND_c_6288_n 0.00525833f $X=13.945 $Y=0.81 $X2=0
+ $Y2=0
cc_1882 N_S[4]_c_2253_n N_VGND_c_6288_n 0.00862298f $X=14.095 $Y=0.18 $X2=0
+ $Y2=0
cc_1883 N_S[4]_c_2259_n N_VGND_c_6290_n 0.0028166f $X=15.965 $Y=0.18 $X2=0 $Y2=0
cc_1884 N_S[4]_c_2260_n N_VGND_c_6290_n 5.5039e-19 $X=16.04 $Y=0.255 $X2=0 $Y2=0
cc_1885 N_S[4]_c_2246_n N_VGND_c_6328_n 0.00585385f $X=13.065 $Y=0.735 $X2=0
+ $Y2=0
cc_1886 N_S[4]_c_2247_n N_VGND_c_6328_n 2.16067e-19 $X=13.41 $Y=0.81 $X2=0 $Y2=0
cc_1887 N_S[4]_c_2248_n N_VGND_c_6328_n 0.00542362f $X=13.485 $Y=0.735 $X2=0
+ $Y2=0
cc_1888 N_S[4]_c_2253_n N_VGND_c_6332_n 0.0559651f $X=14.095 $Y=0.18 $X2=0 $Y2=0
cc_1889 N_S[4]_c_2246_n N_VGND_c_6370_n 0.0119653f $X=13.065 $Y=0.735 $X2=0
+ $Y2=0
cc_1890 N_S[4]_c_2248_n N_VGND_c_6370_n 0.00990284f $X=13.485 $Y=0.735 $X2=0
+ $Y2=0
cc_1891 N_S[4]_c_2252_n N_VGND_c_6370_n 0.0244174f $X=14.705 $Y=0.18 $X2=0 $Y2=0
cc_1892 N_S[4]_c_2253_n N_VGND_c_6370_n 0.0101627f $X=14.095 $Y=0.18 $X2=0 $Y2=0
cc_1893 N_S[4]_c_2255_n N_VGND_c_6370_n 0.00642387f $X=15.125 $Y=0.18 $X2=0
+ $Y2=0
cc_1894 N_S[4]_c_2257_n N_VGND_c_6370_n 0.0064237f $X=15.545 $Y=0.18 $X2=0 $Y2=0
cc_1895 N_S[4]_c_2259_n N_VGND_c_6370_n 0.0123437f $X=15.965 $Y=0.18 $X2=0 $Y2=0
cc_1896 N_S[4]_c_2262_n N_VGND_c_6370_n 0.00366655f $X=14.78 $Y=0.18 $X2=0 $Y2=0
cc_1897 N_S[4]_c_2263_n N_VGND_c_6370_n 0.00366655f $X=15.2 $Y=0.18 $X2=0 $Y2=0
cc_1898 N_S[4]_c_2264_n N_VGND_c_6370_n 0.00366655f $X=15.62 $Y=0.18 $X2=0 $Y2=0
cc_1899 N_S[4]_c_2251_n N_A_2889_66#_c_7254_n 0.00529837f $X=14.02 $Y=0.735
+ $X2=0 $Y2=0
cc_1900 N_S[4]_c_2254_n N_A_2889_66#_c_7255_n 0.0112916f $X=14.78 $Y=0.255 $X2=0
+ $Y2=0
cc_1901 N_S[4]_c_2255_n N_A_2889_66#_c_7255_n 0.00211351f $X=15.125 $Y=0.18
+ $X2=0 $Y2=0
cc_1902 N_S[4]_c_2256_n N_A_2889_66#_c_7255_n 0.0106844f $X=15.2 $Y=0.255 $X2=0
+ $Y2=0
cc_1903 N_S[4]_c_2251_n N_A_2889_66#_c_7256_n 0.00189496f $X=14.02 $Y=0.735
+ $X2=0 $Y2=0
cc_1904 N_S[4]_c_2252_n N_A_2889_66#_c_7256_n 0.00685838f $X=14.705 $Y=0.18
+ $X2=0 $Y2=0
cc_1905 N_S[4]_c_2258_n N_A_2889_66#_c_7257_n 0.0106826f $X=15.62 $Y=0.255 $X2=0
+ $Y2=0
cc_1906 N_S[4]_c_2259_n N_A_2889_66#_c_7257_n 0.00211351f $X=15.965 $Y=0.18
+ $X2=0 $Y2=0
cc_1907 N_S[4]_c_2260_n N_A_2889_66#_c_7257_n 0.0139014f $X=16.04 $Y=0.255 $X2=0
+ $Y2=0
cc_1908 N_S[4]_c_2260_n N_A_2889_66#_c_7260_n 0.00206084f $X=16.04 $Y=0.255
+ $X2=0 $Y2=0
cc_1909 N_S[4]_c_2257_n N_A_2889_66#_c_7273_n 0.0034777f $X=15.545 $Y=0.18 $X2=0
+ $Y2=0
cc_1910 N_S[5]_c_2373_n N_A_2626_599#_c_2616_n 0.00507688f $X=14.78 $Y=5.185
+ $X2=0 $Y2=0
cc_1911 N_S[5]_c_2388_n N_A_2626_599#_c_2608_n 0.00262132f $X=13.51 $Y=3.99
+ $X2=0 $Y2=0
cc_1912 N_S[5]_c_2375_n N_A_2626_599#_c_2619_n 0.00509204f $X=15.2 $Y=5.185
+ $X2=0 $Y2=0
cc_1913 N_S[5]_c_2379_n N_A_2626_599#_c_2621_n 0.00507426f $X=16.04 $Y=5.185
+ $X2=0 $Y2=0
cc_1914 N_S[5]_c_2377_n N_A_2626_599#_c_2624_n 0.00509391f $X=15.62 $Y=5.185
+ $X2=0 $Y2=0
cc_1915 N_S[5]_c_2386_n N_A_2626_599#_c_2625_n 0.00929139f $X=13.04 $Y=3.89
+ $X2=0 $Y2=0
cc_1916 N_S[5]_c_2390_n N_A_2626_599#_c_2625_n 0.00970559f $X=13.51 $Y=3.89
+ $X2=0 $Y2=0
cc_1917 N_S[5]_c_2365_n N_A_2626_599#_c_2609_n 0.00207203f $X=13.065 $Y=4.705
+ $X2=0 $Y2=0
cc_1918 N_S[5]_c_2366_n N_A_2626_599#_c_2609_n 0.0111895f $X=13.41 $Y=4.63 $X2=0
+ $Y2=0
cc_1919 N_S[5]_c_2368_n N_A_2626_599#_c_2609_n 9.67113e-19 $X=13.485 $Y=4.705
+ $X2=0 $Y2=0
cc_1920 N_S[5]_c_2370_n N_A_2626_599#_c_2609_n 6.53442e-19 $X=14.02 $Y=5.185
+ $X2=0 $Y2=0
cc_1921 N_S[5]_c_2380_n N_A_2626_599#_c_2609_n 0.00426435f $X=13.51 $Y=4.63
+ $X2=0 $Y2=0
cc_1922 N_S[5]_c_2368_n N_A_2626_599#_c_2610_n 0.00603996f $X=13.485 $Y=4.705
+ $X2=0 $Y2=0
cc_1923 N_S[5]_c_2386_n N_A_2626_599#_c_2626_n 0.00117303f $X=13.04 $Y=3.89
+ $X2=0 $Y2=0
cc_1924 N_S[5]_c_2365_n N_A_2626_599#_c_2626_n 0.00336772f $X=13.065 $Y=4.705
+ $X2=0 $Y2=0
cc_1925 N_S[5]_c_2388_n N_A_2626_599#_c_2626_n 0.00508008f $X=13.51 $Y=3.99
+ $X2=0 $Y2=0
cc_1926 N_S[5]_c_2367_n N_A_2626_599#_c_2626_n 0.00255921f $X=13.51 $Y=4.555
+ $X2=0 $Y2=0
cc_1927 N_S[5]_c_2390_n N_A_2626_599#_c_2626_n 0.00254107f $X=13.51 $Y=3.89
+ $X2=0 $Y2=0
cc_1928 N_S[5]_c_2367_n N_A_2626_599#_c_2611_n 0.0206368f $X=13.51 $Y=4.555
+ $X2=0 $Y2=0
cc_1929 N_S[5]_c_2369_n N_A_2626_599#_c_2611_n 0.0103812f $X=13.945 $Y=4.63
+ $X2=0 $Y2=0
cc_1930 N_S[5]_c_2386_n N_A_2626_599#_c_2628_n 0.00304348f $X=13.04 $Y=3.89
+ $X2=0 $Y2=0
cc_1931 N_S[5]_c_2365_n N_A_2626_599#_c_2628_n 5.48523e-19 $X=13.065 $Y=4.705
+ $X2=0 $Y2=0
cc_1932 N_S[5]_c_2390_n N_A_2626_599#_c_2628_n 0.00216424f $X=13.51 $Y=3.89
+ $X2=0 $Y2=0
cc_1933 N_S[5]_c_2365_n N_A_2626_599#_c_2612_n 0.00289358f $X=13.065 $Y=4.705
+ $X2=0 $Y2=0
cc_1934 N_S[5]_c_2366_n N_A_2626_599#_c_2612_n 0.00429801f $X=13.41 $Y=4.63
+ $X2=0 $Y2=0
cc_1935 N_S[5]_c_2367_n N_A_2626_599#_c_2612_n 0.0085951f $X=13.51 $Y=4.555
+ $X2=0 $Y2=0
cc_1936 N_S[5]_c_2380_n N_A_2626_599#_c_2612_n 0.00268644f $X=13.51 $Y=4.63
+ $X2=0 $Y2=0
cc_1937 N_S[5]_c_2384_n N_A_2626_599#_c_2612_n 0.00541767f $X=13 $Y=4.28 $X2=0
+ $Y2=0
cc_1938 N_S[5]_c_2365_n N_A_2626_599#_c_2613_n 0.00416423f $X=13.065 $Y=4.705
+ $X2=0 $Y2=0
cc_1939 N_S[5]_c_2367_n N_A_2626_599#_c_2613_n 0.00322131f $X=13.51 $Y=4.555
+ $X2=0 $Y2=0
cc_1940 N_S[5]_c_2384_n N_A_2626_599#_c_2613_n 0.0228692f $X=13 $Y=4.28 $X2=0
+ $Y2=0
cc_1941 N_S[5]_c_2367_n N_A_2626_599#_c_2614_n 0.0175393f $X=13.51 $Y=4.555
+ $X2=0 $Y2=0
cc_1942 N_S[5]_c_2369_n N_A_2626_599#_c_2614_n 0.0179529f $X=13.945 $Y=4.63
+ $X2=0 $Y2=0
cc_1943 N_S[5]_c_2364_n N_VPWR_c_3607_n 0.00652399f $X=12.94 $Y=4.28 $X2=0 $Y2=0
cc_1944 N_S[5]_c_2386_n N_VPWR_c_3607_n 0.00986205f $X=13.04 $Y=3.89 $X2=0 $Y2=0
cc_1945 N_S[5]_c_2384_n N_VPWR_c_3607_n 0.0157609f $X=13 $Y=4.28 $X2=0 $Y2=0
cc_1946 N_S[5]_c_2390_n N_VPWR_c_3609_n 0.00950399f $X=13.51 $Y=3.89 $X2=0 $Y2=0
cc_1947 N_S[5]_c_2386_n N_VPWR_c_3635_n 0.0035837f $X=13.04 $Y=3.89 $X2=0 $Y2=0
cc_1948 N_S[5]_c_2390_n N_VPWR_c_3635_n 0.0035837f $X=13.51 $Y=3.89 $X2=0 $Y2=0
cc_1949 N_S[5]_c_2386_n N_VPWR_c_3661_n 0.0070533f $X=13.04 $Y=3.89 $X2=0 $Y2=0
cc_1950 N_S[5]_c_2390_n N_VPWR_c_3661_n 0.00711603f $X=13.51 $Y=3.89 $X2=0 $Y2=0
cc_1951 N_S[5]_c_2373_n N_Z_c_4599_n 0.0134253f $X=14.78 $Y=5.185 $X2=0 $Y2=0
cc_1952 N_S[5]_c_2375_n N_Z_c_4599_n 0.0077801f $X=15.2 $Y=5.185 $X2=0 $Y2=0
cc_1953 N_S[5]_c_2377_n N_Z_c_4599_n 6.35774e-19 $X=15.62 $Y=5.185 $X2=0 $Y2=0
cc_1954 N_S[5]_c_2375_n N_Z_c_4601_n 0.00190704f $X=15.2 $Y=5.185 $X2=0 $Y2=0
cc_1955 N_S[5]_c_2377_n N_Z_c_4601_n 3.10191e-19 $X=15.62 $Y=5.185 $X2=0 $Y2=0
cc_1956 N_S[5]_c_2373_n N_Z_c_4623_n 0.00216436f $X=14.78 $Y=5.185 $X2=0 $Y2=0
cc_1957 N_S[5]_c_2377_n N_Z_c_4625_n 0.00180363f $X=15.62 $Y=5.185 $X2=0 $Y2=0
cc_1958 N_S[5]_c_2377_n N_Z_c_4627_n 0.00462308f $X=15.62 $Y=5.185 $X2=0 $Y2=0
cc_1959 N_S[5]_c_2379_n N_Z_c_4627_n 0.00443615f $X=16.04 $Y=5.185 $X2=0 $Y2=0
cc_1960 N_S[5]_c_2375_n N_Z_c_4628_n 6.35664e-19 $X=15.2 $Y=5.185 $X2=0 $Y2=0
cc_1961 N_S[5]_c_2377_n N_Z_c_4628_n 0.00283489f $X=15.62 $Y=5.185 $X2=0 $Y2=0
cc_1962 N_S[5]_c_2379_n N_Z_c_4628_n 0.002324f $X=16.04 $Y=5.185 $X2=0 $Y2=0
cc_1963 N_S[5]_c_2364_n N_Z_c_4647_n 0.00234109f $X=12.94 $Y=4.28 $X2=0 $Y2=0
cc_1964 N_S[5]_c_2386_n N_Z_c_4647_n 0.00501777f $X=13.04 $Y=3.89 $X2=0 $Y2=0
cc_1965 N_S[5]_c_2365_n N_Z_c_4647_n 2.32936e-19 $X=13.065 $Y=4.705 $X2=0 $Y2=0
cc_1966 N_S[5]_c_2388_n N_Z_c_4647_n 2.55735e-19 $X=13.51 $Y=3.99 $X2=0 $Y2=0
cc_1967 N_S[5]_c_2390_n N_Z_c_4647_n 0.00453198f $X=13.51 $Y=3.89 $X2=0 $Y2=0
cc_1968 N_S[5]_c_2384_n N_Z_c_4647_n 0.0105931f $X=13 $Y=4.28 $X2=0 $Y2=0
cc_1969 N_S[5]_c_2379_n N_A_2839_613#_c_5890_n 0.00168571f $X=16.04 $Y=5.185
+ $X2=0 $Y2=0
cc_1970 N_S[5]_c_2390_n N_A_2839_613#_c_5892_n 0.00239129f $X=13.51 $Y=3.89
+ $X2=0 $Y2=0
cc_1971 N_S[5]_c_2364_n N_VGND_c_6287_n 0.00576464f $X=12.94 $Y=4.28 $X2=0 $Y2=0
cc_1972 N_S[5]_c_2365_n N_VGND_c_6287_n 0.00374526f $X=13.065 $Y=4.705 $X2=0
+ $Y2=0
cc_1973 N_S[5]_c_2384_n N_VGND_c_6287_n 0.0116218f $X=13 $Y=4.28 $X2=0 $Y2=0
cc_1974 N_S[5]_c_2368_n N_VGND_c_6289_n 0.00173127f $X=13.485 $Y=4.705 $X2=0
+ $Y2=0
cc_1975 N_S[5]_c_2369_n N_VGND_c_6289_n 0.00525833f $X=13.945 $Y=4.63 $X2=0
+ $Y2=0
cc_1976 N_S[5]_c_2370_n N_VGND_c_6289_n 0.00862298f $X=14.02 $Y=5.185 $X2=0
+ $Y2=0
cc_1977 N_S[5]_c_2378_n N_VGND_c_6291_n 0.0028166f $X=15.965 $Y=5.26 $X2=0 $Y2=0
cc_1978 N_S[5]_c_2379_n N_VGND_c_6291_n 5.5039e-19 $X=16.04 $Y=5.185 $X2=0 $Y2=0
cc_1979 N_S[5]_c_2365_n N_VGND_c_6330_n 0.00585385f $X=13.065 $Y=4.705 $X2=0
+ $Y2=0
cc_1980 N_S[5]_c_2366_n N_VGND_c_6330_n 2.16067e-19 $X=13.41 $Y=4.63 $X2=0 $Y2=0
cc_1981 N_S[5]_c_2368_n N_VGND_c_6330_n 0.00542362f $X=13.485 $Y=4.705 $X2=0
+ $Y2=0
cc_1982 N_S[5]_c_2372_n N_VGND_c_6334_n 0.0559651f $X=14.095 $Y=5.26 $X2=0 $Y2=0
cc_1983 N_S[5]_c_2365_n N_VGND_c_6371_n 0.0119653f $X=13.065 $Y=4.705 $X2=0
+ $Y2=0
cc_1984 N_S[5]_c_2368_n N_VGND_c_6371_n 0.00990284f $X=13.485 $Y=4.705 $X2=0
+ $Y2=0
cc_1985 N_S[5]_c_2371_n N_VGND_c_6371_n 0.0244174f $X=14.705 $Y=5.26 $X2=0 $Y2=0
cc_1986 N_S[5]_c_2372_n N_VGND_c_6371_n 0.0101627f $X=14.095 $Y=5.26 $X2=0 $Y2=0
cc_1987 N_S[5]_c_2374_n N_VGND_c_6371_n 0.00642387f $X=15.125 $Y=5.26 $X2=0
+ $Y2=0
cc_1988 N_S[5]_c_2376_n N_VGND_c_6371_n 0.0064237f $X=15.545 $Y=5.26 $X2=0 $Y2=0
cc_1989 N_S[5]_c_2378_n N_VGND_c_6371_n 0.0123437f $X=15.965 $Y=5.26 $X2=0 $Y2=0
cc_1990 N_S[5]_c_2381_n N_VGND_c_6371_n 0.00366655f $X=14.78 $Y=5.26 $X2=0 $Y2=0
cc_1991 N_S[5]_c_2382_n N_VGND_c_6371_n 0.00366655f $X=15.2 $Y=5.26 $X2=0 $Y2=0
cc_1992 N_S[5]_c_2383_n N_VGND_c_6371_n 0.00366655f $X=15.62 $Y=5.26 $X2=0 $Y2=0
cc_1993 N_S[5]_c_2369_n N_A_2889_918#_c_7338_n 0.00529837f $X=13.945 $Y=4.63
+ $X2=0 $Y2=0
cc_1994 N_S[5]_c_2373_n N_A_2889_918#_c_7339_n 0.0112916f $X=14.78 $Y=5.185
+ $X2=0 $Y2=0
cc_1995 N_S[5]_c_2374_n N_A_2889_918#_c_7339_n 0.00211351f $X=15.125 $Y=5.26
+ $X2=0 $Y2=0
cc_1996 N_S[5]_c_2375_n N_A_2889_918#_c_7339_n 0.0106844f $X=15.2 $Y=5.185 $X2=0
+ $Y2=0
cc_1997 N_S[5]_c_2370_n N_A_2889_918#_c_7340_n 0.00189496f $X=14.02 $Y=5.185
+ $X2=0 $Y2=0
cc_1998 N_S[5]_c_2371_n N_A_2889_918#_c_7340_n 0.00685838f $X=14.705 $Y=5.26
+ $X2=0 $Y2=0
cc_1999 N_S[5]_c_2377_n N_A_2889_918#_c_7341_n 0.0106826f $X=15.62 $Y=5.185
+ $X2=0 $Y2=0
cc_2000 N_S[5]_c_2378_n N_A_2889_918#_c_7341_n 0.00211351f $X=15.965 $Y=5.26
+ $X2=0 $Y2=0
cc_2001 N_S[5]_c_2379_n N_A_2889_918#_c_7341_n 0.0139014f $X=16.04 $Y=5.185
+ $X2=0 $Y2=0
cc_2002 N_S[5]_c_2379_n N_A_2889_918#_c_7344_n 0.00206084f $X=16.04 $Y=5.185
+ $X2=0 $Y2=0
cc_2003 N_S[5]_c_2376_n N_A_2889_918#_c_7357_n 0.0034777f $X=15.545 $Y=5.26
+ $X2=0 $Y2=0
cc_2004 N_A_2626_325#_c_2499_n N_A_2626_599#_c_2615_n 0.0129371f $X=14.555
+ $Y=1.475 $X2=0 $Y2=0
cc_2005 N_A_2626_325#_c_2502_n N_A_2626_599#_c_2618_n 0.0129371f $X=15.025
+ $Y=1.475 $X2=0 $Y2=0
cc_2006 N_A_2626_325#_c_2504_n N_A_2626_599#_c_2620_n 0.0129371f $X=15.495
+ $Y=1.475 $X2=0 $Y2=0
cc_2007 N_A_2626_325#_c_2506_n N_A_2626_599#_c_2622_n 0.0129371f $X=15.965
+ $Y=1.475 $X2=0 $Y2=0
cc_2008 N_A_2626_325#_c_2509_n N_VPWR_c_3606_n 0.0356181f $X=13.275 $Y=1.77
+ $X2=0 $Y2=0
cc_2009 N_A_2626_325#_c_2499_n N_VPWR_c_3608_n 0.00367058f $X=14.555 $Y=1.475
+ $X2=0 $Y2=0
cc_2010 N_A_2626_325#_c_2509_n N_VPWR_c_3608_n 0.0316788f $X=13.275 $Y=1.77
+ $X2=0 $Y2=0
cc_2011 N_A_2626_325#_c_2495_n N_VPWR_c_3608_n 0.0193185f $X=14.325 $Y=1.23
+ $X2=0 $Y2=0
cc_2012 N_A_2626_325#_c_2498_n N_VPWR_c_3608_n 6.4101e-19 $X=14.235 $Y=1.23
+ $X2=0 $Y2=0
cc_2013 N_A_2626_325#_c_2506_n N_VPWR_c_3610_n 0.00324472f $X=15.965 $Y=1.475
+ $X2=0 $Y2=0
cc_2014 N_A_2626_325#_c_2509_n N_VPWR_c_3635_n 0.0233824f $X=13.275 $Y=1.77
+ $X2=0 $Y2=0
cc_2015 N_A_2626_325#_c_2499_n N_VPWR_c_3661_n 0.00473731f $X=14.555 $Y=1.475
+ $X2=0 $Y2=0
cc_2016 N_A_2626_325#_c_2502_n N_VPWR_c_3661_n 0.00362156f $X=15.025 $Y=1.475
+ $X2=0 $Y2=0
cc_2017 N_A_2626_325#_c_2504_n N_VPWR_c_3661_n 0.00362156f $X=15.495 $Y=1.475
+ $X2=0 $Y2=0
cc_2018 N_A_2626_325#_c_2506_n N_VPWR_c_3661_n 0.00473731f $X=15.965 $Y=1.475
+ $X2=0 $Y2=0
cc_2019 N_A_2626_325#_c_2509_n N_VPWR_c_3661_n 0.00593513f $X=13.275 $Y=1.77
+ $X2=0 $Y2=0
cc_2020 N_A_2626_325#_c_2503_n N_Z_c_4600_n 0.00762343f $X=15.405 $Y=1.4 $X2=0
+ $Y2=0
cc_2021 N_A_2626_325#_c_2508_n N_Z_c_4600_n 0.00704092f $X=15.495 $Y=1.4 $X2=0
+ $Y2=0
cc_2022 N_A_2626_325#_c_2500_n N_Z_c_4622_n 0.00597584f $X=14.935 $Y=1.4 $X2=0
+ $Y2=0
cc_2023 N_A_2626_325#_c_2492_n N_Z_c_4622_n 0.00747617f $X=14.645 $Y=1.4 $X2=0
+ $Y2=0
cc_2024 N_A_2626_325#_c_2503_n N_Z_c_4622_n 0.00145542f $X=15.405 $Y=1.4 $X2=0
+ $Y2=0
cc_2025 N_A_2626_325#_c_2507_n N_Z_c_4622_n 0.00909323f $X=15.025 $Y=1.4 $X2=0
+ $Y2=0
cc_2026 N_A_2626_325#_c_2495_n N_Z_c_4622_n 0.0266078f $X=14.325 $Y=1.23 $X2=0
+ $Y2=0
cc_2027 N_A_2626_325#_c_2505_n N_Z_c_4624_n 0.00918337f $X=15.875 $Y=1.4 $X2=0
+ $Y2=0
cc_2028 N_A_2626_325#_c_2508_n N_Z_c_4624_n 2.98555e-19 $X=15.495 $Y=1.4 $X2=0
+ $Y2=0
cc_2029 N_A_2626_325#_c_2505_n N_Z_c_4626_n 0.00248496f $X=15.875 $Y=1.4 $X2=0
+ $Y2=0
cc_2030 N_A_2626_325#_c_2499_n N_Z_c_4646_n 0.00795576f $X=14.555 $Y=1.475 $X2=0
+ $Y2=0
cc_2031 N_A_2626_325#_c_2492_n N_Z_c_4646_n 2.19754e-19 $X=14.645 $Y=1.4 $X2=0
+ $Y2=0
cc_2032 N_A_2626_325#_c_2509_n N_Z_c_4646_n 0.0329704f $X=13.275 $Y=1.77 $X2=0
+ $Y2=0
cc_2033 N_A_2626_325#_c_2495_n N_Z_c_4646_n 0.0186685f $X=14.325 $Y=1.23 $X2=0
+ $Y2=0
cc_2034 N_A_2626_325#_c_2506_n N_Z_c_4648_n 0.00834829f $X=15.965 $Y=1.475 $X2=0
+ $Y2=0
cc_2035 N_A_2626_325#_c_2502_n N_Z_c_4895_n 0.00372248f $X=15.025 $Y=1.475 $X2=0
+ $Y2=0
cc_2036 N_A_2626_325#_c_2504_n N_Z_c_4895_n 0.00372458f $X=15.495 $Y=1.475 $X2=0
+ $Y2=0
cc_2037 N_A_2626_325#_c_2499_n N_Z_c_4654_n 0.0221748f $X=14.555 $Y=1.475 $X2=0
+ $Y2=0
cc_2038 N_A_2626_325#_c_2500_n N_Z_c_4654_n 0.00560592f $X=14.935 $Y=1.4 $X2=0
+ $Y2=0
cc_2039 N_A_2626_325#_c_2492_n N_Z_c_4654_n 0.00425035f $X=14.645 $Y=1.4 $X2=0
+ $Y2=0
cc_2040 N_A_2626_325#_c_2502_n N_Z_c_4654_n 0.0181262f $X=15.025 $Y=1.475 $X2=0
+ $Y2=0
cc_2041 N_A_2626_325#_c_2504_n N_Z_c_4654_n 9.74366e-19 $X=15.495 $Y=1.475 $X2=0
+ $Y2=0
cc_2042 N_A_2626_325#_c_2507_n N_Z_c_4654_n 0.00181273f $X=15.025 $Y=1.4 $X2=0
+ $Y2=0
cc_2043 N_A_2626_325#_c_2495_n N_Z_c_4654_n 0.00240108f $X=14.325 $Y=1.23 $X2=0
+ $Y2=0
cc_2044 N_A_2626_325#_c_2502_n N_Z_c_4655_n 9.74366e-19 $X=15.025 $Y=1.475 $X2=0
+ $Y2=0
cc_2045 N_A_2626_325#_c_2504_n N_Z_c_4655_n 0.0181262f $X=15.495 $Y=1.475 $X2=0
+ $Y2=0
cc_2046 N_A_2626_325#_c_2505_n N_Z_c_4655_n 0.0103509f $X=15.875 $Y=1.4 $X2=0
+ $Y2=0
cc_2047 N_A_2626_325#_c_2506_n N_Z_c_4655_n 0.0199111f $X=15.965 $Y=1.475 $X2=0
+ $Y2=0
cc_2048 N_A_2626_325#_c_2508_n N_Z_c_4655_n 0.00415268f $X=15.495 $Y=1.4 $X2=0
+ $Y2=0
cc_2049 N_A_2626_325#_c_2506_n N_A_2839_311#_c_5759_n 0.00151141f $X=15.965
+ $Y=1.475 $X2=0 $Y2=0
cc_2050 N_A_2626_325#_c_2499_n N_A_2839_311#_c_5767_n 0.00307958f $X=14.555
+ $Y=1.475 $X2=0 $Y2=0
cc_2051 N_A_2626_325#_c_2502_n N_A_2839_311#_c_5767_n 0.00307958f $X=15.025
+ $Y=1.475 $X2=0 $Y2=0
cc_2052 N_A_2626_325#_c_2504_n N_A_2839_311#_c_5769_n 0.00307958f $X=15.495
+ $Y=1.475 $X2=0 $Y2=0
cc_2053 N_A_2626_325#_c_2506_n N_A_2839_311#_c_5769_n 0.00307958f $X=15.965
+ $Y=1.475 $X2=0 $Y2=0
cc_2054 N_A_2626_325#_c_2499_n N_A_2839_311#_c_5761_n 0.00499839f $X=14.555
+ $Y=1.475 $X2=0 $Y2=0
cc_2055 N_A_2626_325#_c_2492_n N_A_2839_311#_c_5761_n 0.00561627f $X=14.645
+ $Y=1.4 $X2=0 $Y2=0
cc_2056 N_A_2626_325#_c_2495_n N_A_2839_311#_c_5761_n 0.0218124f $X=14.325
+ $Y=1.23 $X2=0 $Y2=0
cc_2057 N_A_2626_325#_c_2498_n N_A_2839_311#_c_5761_n 5.74251e-19 $X=14.235
+ $Y=1.23 $X2=0 $Y2=0
cc_2058 N_A_2626_325#_c_2502_n N_A_2839_311#_c_5762_n 0.00210632f $X=15.025
+ $Y=1.475 $X2=0 $Y2=0
cc_2059 N_A_2626_325#_c_2503_n N_A_2839_311#_c_5762_n 0.00251792f $X=15.405
+ $Y=1.4 $X2=0 $Y2=0
cc_2060 N_A_2626_325#_c_2504_n N_A_2839_311#_c_5762_n 0.00210632f $X=15.495
+ $Y=1.475 $X2=0 $Y2=0
cc_2061 N_A_2626_325#_c_2506_n N_A_2839_311#_c_5763_n 0.00554566f $X=15.965
+ $Y=1.475 $X2=0 $Y2=0
cc_2062 N_A_2626_325#_c_2495_n N_VGND_c_6288_n 0.0123065f $X=14.325 $Y=1.23
+ $X2=0 $Y2=0
cc_2063 N_A_2626_325#_c_2498_n N_VGND_c_6288_n 2.04129e-19 $X=14.235 $Y=1.23
+ $X2=0 $Y2=0
cc_2064 N_A_2626_325#_c_2493_n N_VGND_c_6328_n 0.0129994f $X=13.275 $Y=0.445
+ $X2=0 $Y2=0
cc_2065 N_A_2626_325#_M1121_s N_VGND_c_6370_n 0.00394793f $X=13.14 $Y=0.235
+ $X2=0 $Y2=0
cc_2066 N_A_2626_325#_c_2493_n N_VGND_c_6370_n 0.00927134f $X=13.275 $Y=0.445
+ $X2=0 $Y2=0
cc_2067 N_A_2626_325#_c_2492_n N_A_2889_66#_c_7254_n 0.00600378f $X=14.645
+ $Y=1.4 $X2=0 $Y2=0
cc_2068 N_A_2626_325#_c_2495_n N_A_2889_66#_c_7254_n 0.0028695f $X=14.325
+ $Y=1.23 $X2=0 $Y2=0
cc_2069 N_A_2626_325#_c_2503_n N_A_2889_66#_c_7276_n 7.0477e-19 $X=15.405 $Y=1.4
+ $X2=0 $Y2=0
cc_2070 N_A_2626_599#_c_2625_n N_VPWR_c_3607_n 0.0356181f $X=13.275 $Y=3.14
+ $X2=0 $Y2=0
cc_2071 N_A_2626_599#_c_2615_n N_VPWR_c_3609_n 0.00367058f $X=14.555 $Y=3.965
+ $X2=0 $Y2=0
cc_2072 N_A_2626_599#_c_2625_n N_VPWR_c_3609_n 0.0316788f $X=13.275 $Y=3.14
+ $X2=0 $Y2=0
cc_2073 N_A_2626_599#_c_2611_n N_VPWR_c_3609_n 0.0193185f $X=14.325 $Y=4.21
+ $X2=0 $Y2=0
cc_2074 N_A_2626_599#_c_2614_n N_VPWR_c_3609_n 6.4101e-19 $X=14.235 $Y=4.21
+ $X2=0 $Y2=0
cc_2075 N_A_2626_599#_c_2622_n N_VPWR_c_3611_n 0.00324472f $X=15.965 $Y=3.965
+ $X2=0 $Y2=0
cc_2076 N_A_2626_599#_c_2625_n N_VPWR_c_3635_n 0.0233824f $X=13.275 $Y=3.14
+ $X2=0 $Y2=0
cc_2077 N_A_2626_599#_c_2615_n N_VPWR_c_3661_n 0.00473731f $X=14.555 $Y=3.965
+ $X2=0 $Y2=0
cc_2078 N_A_2626_599#_c_2618_n N_VPWR_c_3661_n 0.00362156f $X=15.025 $Y=3.965
+ $X2=0 $Y2=0
cc_2079 N_A_2626_599#_c_2620_n N_VPWR_c_3661_n 0.00362156f $X=15.495 $Y=3.965
+ $X2=0 $Y2=0
cc_2080 N_A_2626_599#_c_2622_n N_VPWR_c_3661_n 0.00473731f $X=15.965 $Y=3.965
+ $X2=0 $Y2=0
cc_2081 N_A_2626_599#_c_2625_n N_VPWR_c_3661_n 0.00593513f $X=13.275 $Y=3.14
+ $X2=0 $Y2=0
cc_2082 N_A_2626_599#_c_2619_n N_Z_c_4601_n 0.00762343f $X=15.405 $Y=4.04 $X2=0
+ $Y2=0
cc_2083 N_A_2626_599#_c_2624_n N_Z_c_4601_n 0.00704092f $X=15.495 $Y=4.04 $X2=0
+ $Y2=0
cc_2084 N_A_2626_599#_c_2616_n N_Z_c_4623_n 0.00597584f $X=14.935 $Y=4.04 $X2=0
+ $Y2=0
cc_2085 N_A_2626_599#_c_2608_n N_Z_c_4623_n 0.00747617f $X=14.645 $Y=4.04 $X2=0
+ $Y2=0
cc_2086 N_A_2626_599#_c_2619_n N_Z_c_4623_n 0.00145542f $X=15.405 $Y=4.04 $X2=0
+ $Y2=0
cc_2087 N_A_2626_599#_c_2623_n N_Z_c_4623_n 0.00909323f $X=15.025 $Y=4.04 $X2=0
+ $Y2=0
cc_2088 N_A_2626_599#_c_2611_n N_Z_c_4623_n 0.0266078f $X=14.325 $Y=4.21 $X2=0
+ $Y2=0
cc_2089 N_A_2626_599#_c_2621_n N_Z_c_4625_n 0.00918337f $X=15.875 $Y=4.04 $X2=0
+ $Y2=0
cc_2090 N_A_2626_599#_c_2624_n N_Z_c_4625_n 2.98555e-19 $X=15.495 $Y=4.04 $X2=0
+ $Y2=0
cc_2091 N_A_2626_599#_c_2621_n N_Z_c_4627_n 0.00248496f $X=15.875 $Y=4.04 $X2=0
+ $Y2=0
cc_2092 N_A_2626_599#_c_2615_n N_Z_c_4647_n 0.00795576f $X=14.555 $Y=3.965 $X2=0
+ $Y2=0
cc_2093 N_A_2626_599#_c_2608_n N_Z_c_4647_n 2.19754e-19 $X=14.645 $Y=4.04 $X2=0
+ $Y2=0
cc_2094 N_A_2626_599#_c_2625_n N_Z_c_4647_n 0.0329704f $X=13.275 $Y=3.14 $X2=0
+ $Y2=0
cc_2095 N_A_2626_599#_c_2611_n N_Z_c_4647_n 0.0186685f $X=14.325 $Y=4.21 $X2=0
+ $Y2=0
cc_2096 N_A_2626_599#_c_2622_n N_Z_c_4649_n 0.00834829f $X=15.965 $Y=3.965 $X2=0
+ $Y2=0
cc_2097 N_A_2626_599#_c_2618_n N_Z_c_4924_n 0.00372248f $X=15.025 $Y=3.965 $X2=0
+ $Y2=0
cc_2098 N_A_2626_599#_c_2620_n N_Z_c_4924_n 0.00372458f $X=15.495 $Y=3.965 $X2=0
+ $Y2=0
cc_2099 N_A_2626_599#_c_2615_n N_Z_c_4654_n 0.0221748f $X=14.555 $Y=3.965 $X2=0
+ $Y2=0
cc_2100 N_A_2626_599#_c_2616_n N_Z_c_4654_n 0.00560592f $X=14.935 $Y=4.04 $X2=0
+ $Y2=0
cc_2101 N_A_2626_599#_c_2608_n N_Z_c_4654_n 0.00425035f $X=14.645 $Y=4.04 $X2=0
+ $Y2=0
cc_2102 N_A_2626_599#_c_2618_n N_Z_c_4654_n 0.0181262f $X=15.025 $Y=3.965 $X2=0
+ $Y2=0
cc_2103 N_A_2626_599#_c_2620_n N_Z_c_4654_n 9.74366e-19 $X=15.495 $Y=3.965 $X2=0
+ $Y2=0
cc_2104 N_A_2626_599#_c_2623_n N_Z_c_4654_n 0.00181273f $X=15.025 $Y=4.04 $X2=0
+ $Y2=0
cc_2105 N_A_2626_599#_c_2611_n N_Z_c_4654_n 0.00240108f $X=14.325 $Y=4.21 $X2=0
+ $Y2=0
cc_2106 N_A_2626_599#_c_2618_n N_Z_c_4655_n 9.74366e-19 $X=15.025 $Y=3.965 $X2=0
+ $Y2=0
cc_2107 N_A_2626_599#_c_2620_n N_Z_c_4655_n 0.0181262f $X=15.495 $Y=3.965 $X2=0
+ $Y2=0
cc_2108 N_A_2626_599#_c_2621_n N_Z_c_4655_n 0.0103509f $X=15.875 $Y=4.04 $X2=0
+ $Y2=0
cc_2109 N_A_2626_599#_c_2622_n N_Z_c_4655_n 0.0199111f $X=15.965 $Y=3.965 $X2=0
+ $Y2=0
cc_2110 N_A_2626_599#_c_2624_n N_Z_c_4655_n 0.00415268f $X=15.495 $Y=4.04 $X2=0
+ $Y2=0
cc_2111 N_A_2626_599#_c_2622_n N_A_2839_613#_c_5890_n 0.00151141f $X=15.965
+ $Y=3.965 $X2=0 $Y2=0
cc_2112 N_A_2626_599#_c_2615_n N_A_2839_613#_c_5898_n 0.00307958f $X=14.555
+ $Y=3.965 $X2=0 $Y2=0
cc_2113 N_A_2626_599#_c_2618_n N_A_2839_613#_c_5898_n 0.00307958f $X=15.025
+ $Y=3.965 $X2=0 $Y2=0
cc_2114 N_A_2626_599#_c_2620_n N_A_2839_613#_c_5900_n 0.00307958f $X=15.495
+ $Y=3.965 $X2=0 $Y2=0
cc_2115 N_A_2626_599#_c_2622_n N_A_2839_613#_c_5900_n 0.00307958f $X=15.965
+ $Y=3.965 $X2=0 $Y2=0
cc_2116 N_A_2626_599#_c_2615_n N_A_2839_613#_c_5892_n 0.00499839f $X=14.555
+ $Y=3.965 $X2=0 $Y2=0
cc_2117 N_A_2626_599#_c_2608_n N_A_2839_613#_c_5892_n 0.00561627f $X=14.645
+ $Y=4.04 $X2=0 $Y2=0
cc_2118 N_A_2626_599#_c_2611_n N_A_2839_613#_c_5892_n 0.0218124f $X=14.325
+ $Y=4.21 $X2=0 $Y2=0
cc_2119 N_A_2626_599#_c_2614_n N_A_2839_613#_c_5892_n 5.74251e-19 $X=14.235
+ $Y=4.21 $X2=0 $Y2=0
cc_2120 N_A_2626_599#_c_2618_n N_A_2839_613#_c_5893_n 0.00210632f $X=15.025
+ $Y=3.965 $X2=0 $Y2=0
cc_2121 N_A_2626_599#_c_2619_n N_A_2839_613#_c_5893_n 0.00251792f $X=15.405
+ $Y=4.04 $X2=0 $Y2=0
cc_2122 N_A_2626_599#_c_2620_n N_A_2839_613#_c_5893_n 0.00210632f $X=15.495
+ $Y=3.965 $X2=0 $Y2=0
cc_2123 N_A_2626_599#_c_2622_n N_A_2839_613#_c_5894_n 0.00554566f $X=15.965
+ $Y=3.965 $X2=0 $Y2=0
cc_2124 N_A_2626_599#_c_2611_n N_VGND_c_6289_n 0.0123065f $X=14.325 $Y=4.21
+ $X2=0 $Y2=0
cc_2125 N_A_2626_599#_c_2614_n N_VGND_c_6289_n 2.04129e-19 $X=14.235 $Y=4.21
+ $X2=0 $Y2=0
cc_2126 N_A_2626_599#_c_2610_n N_VGND_c_6330_n 0.0129994f $X=13.275 $Y=4.995
+ $X2=0 $Y2=0
cc_2127 N_A_2626_599#_M1074_s N_VGND_c_6371_n 0.00394793f $X=13.14 $Y=4.785
+ $X2=0 $Y2=0
cc_2128 N_A_2626_599#_c_2610_n N_VGND_c_6371_n 0.00927134f $X=13.275 $Y=4.995
+ $X2=0 $Y2=0
cc_2129 N_A_2626_599#_c_2608_n N_A_2889_918#_c_7338_n 0.00600378f $X=14.645
+ $Y=4.04 $X2=0 $Y2=0
cc_2130 N_A_2626_599#_c_2611_n N_A_2889_918#_c_7338_n 0.0028695f $X=14.325
+ $Y=4.21 $X2=0 $Y2=0
cc_2131 N_A_2626_599#_c_2619_n N_A_2889_918#_c_7360_n 7.0477e-19 $X=15.405
+ $Y=4.04 $X2=0 $Y2=0
cc_2132 N_D[4]_M1042_g N_D[5]_M1046_g 0.0130744f $X=16.955 $Y=1.985 $X2=0 $Y2=0
cc_2133 N_D[4]_M1062_g N_D[5]_M1070_g 0.0130744f $X=17.425 $Y=1.985 $X2=0 $Y2=0
cc_2134 N_D[4]_M1105_g N_D[5]_M1113_g 0.0130744f $X=17.895 $Y=1.985 $X2=0 $Y2=0
cc_2135 N_D[4]_M1127_g N_D[5]_M1134_g 0.0130744f $X=18.365 $Y=1.985 $X2=0 $Y2=0
cc_2136 N_D[4]_M1127_g N_D[6]_M1082_g 0.0129367f $X=18.365 $Y=1.985 $X2=0 $Y2=0
cc_2137 N_D[4]_M1079_g N_D[6]_M1005_g 0.0210205f $X=18.34 $Y=0.56 $X2=0 $Y2=0
cc_2138 N_D[4]_c_2740_n N_D[6]_c_2935_n 2.99666e-19 $X=18.26 $Y=1.16 $X2=0 $Y2=0
cc_2139 N_D[4]_c_2741_n N_D[6]_c_2935_n 0.0105491f $X=18.365 $Y=1.16 $X2=0 $Y2=0
cc_2140 N_D[4]_c_2740_n N_D[6]_c_2936_n 0.0135469f $X=18.26 $Y=1.16 $X2=0 $Y2=0
cc_2141 N_D[4]_c_2741_n N_D[6]_c_2936_n 2.99666e-19 $X=18.365 $Y=1.16 $X2=0
+ $Y2=0
cc_2142 N_D[4]_M1042_g N_VPWR_c_3610_n 0.00389633f $X=16.955 $Y=1.985 $X2=0
+ $Y2=0
cc_2143 N_D[4]_M1062_g N_VPWR_c_3612_n 0.00208662f $X=17.425 $Y=1.985 $X2=0
+ $Y2=0
cc_2144 N_D[4]_M1105_g N_VPWR_c_3612_n 0.00208662f $X=17.895 $Y=1.985 $X2=0
+ $Y2=0
cc_2145 N_D[4]_M1127_g N_VPWR_c_3614_n 0.00207065f $X=18.365 $Y=1.985 $X2=0
+ $Y2=0
cc_2146 N_D[4]_M1042_g N_VPWR_c_3645_n 0.0035837f $X=16.955 $Y=1.985 $X2=0 $Y2=0
cc_2147 N_D[4]_M1062_g N_VPWR_c_3645_n 0.0035837f $X=17.425 $Y=1.985 $X2=0 $Y2=0
cc_2148 N_D[4]_M1105_g N_VPWR_c_3646_n 0.0035837f $X=17.895 $Y=1.985 $X2=0 $Y2=0
cc_2149 N_D[4]_M1127_g N_VPWR_c_3646_n 0.0035837f $X=18.365 $Y=1.985 $X2=0 $Y2=0
cc_2150 N_D[4]_M1042_g N_VPWR_c_3661_n 0.00573859f $X=16.955 $Y=1.985 $X2=0
+ $Y2=0
cc_2151 N_D[4]_M1062_g N_VPWR_c_3661_n 0.00445624f $X=17.425 $Y=1.985 $X2=0
+ $Y2=0
cc_2152 N_D[4]_M1105_g N_VPWR_c_3661_n 0.00445624f $X=17.895 $Y=1.985 $X2=0
+ $Y2=0
cc_2153 N_D[4]_M1127_g N_VPWR_c_3661_n 0.00579371f $X=18.365 $Y=1.985 $X2=0
+ $Y2=0
cc_2154 N_D[4]_M1042_g N_Z_c_4648_n 0.00311896f $X=16.955 $Y=1.985 $X2=0 $Y2=0
cc_2155 N_D[4]_M1062_g N_Z_c_4648_n 0.00306964f $X=17.425 $Y=1.985 $X2=0 $Y2=0
cc_2156 N_D[4]_M1105_g N_Z_c_4648_n 0.00306964f $X=17.895 $Y=1.985 $X2=0 $Y2=0
cc_2157 N_D[4]_M1127_g N_Z_c_4648_n 0.00470782f $X=18.365 $Y=1.985 $X2=0 $Y2=0
cc_2158 N_D[4]_c_2740_n N_Z_c_4648_n 0.00846955f $X=18.26 $Y=1.16 $X2=0 $Y2=0
cc_2159 N_D[4]_M1042_g N_A_2839_311#_c_5758_n 0.013247f $X=16.955 $Y=1.985 $X2=0
+ $Y2=0
cc_2160 N_D[4]_M1062_g N_A_2839_311#_c_5780_n 0.00916655f $X=17.425 $Y=1.985
+ $X2=0 $Y2=0
cc_2161 N_D[4]_M1105_g N_A_2839_311#_c_5780_n 0.00916655f $X=17.895 $Y=1.985
+ $X2=0 $Y2=0
cc_2162 N_D[4]_c_2738_n N_A_2839_311#_c_5780_n 7.15862e-19 $X=17.805 $Y=1.16
+ $X2=0 $Y2=0
cc_2163 N_D[4]_c_2740_n N_A_2839_311#_c_5780_n 0.0387168f $X=18.26 $Y=1.16 $X2=0
+ $Y2=0
cc_2164 N_D[4]_M1042_g N_A_2839_311#_c_5784_n 8.61029e-19 $X=16.955 $Y=1.985
+ $X2=0 $Y2=0
cc_2165 N_D[4]_M1062_g N_A_2839_311#_c_5784_n 5.79575e-19 $X=17.425 $Y=1.985
+ $X2=0 $Y2=0
cc_2166 N_D[4]_c_2739_n N_A_2839_311#_c_5784_n 8.03631e-19 $X=17.515 $Y=1.16
+ $X2=0 $Y2=0
cc_2167 N_D[4]_c_2740_n N_A_2839_311#_c_5784_n 0.0191156f $X=18.26 $Y=1.16 $X2=0
+ $Y2=0
cc_2168 N_D[4]_M1105_g N_A_2839_311#_c_5788_n 5.79575e-19 $X=17.895 $Y=1.985
+ $X2=0 $Y2=0
cc_2169 N_D[4]_M1127_g N_A_2839_311#_c_5788_n 0.002088f $X=18.365 $Y=1.985 $X2=0
+ $Y2=0
cc_2170 N_D[4]_c_2740_n N_A_2839_311#_c_5788_n 0.0217153f $X=18.26 $Y=1.16 $X2=0
+ $Y2=0
cc_2171 N_D[4]_c_2741_n N_A_2839_311#_c_5788_n 8.03631e-19 $X=18.365 $Y=1.16
+ $X2=0 $Y2=0
cc_2172 N_D[4]_M1042_g N_A_2839_311#_c_5760_n 0.00232998f $X=16.955 $Y=1.985
+ $X2=0 $Y2=0
cc_2173 N_D[4]_M1062_g N_A_2839_311#_c_5793_n 0.00232998f $X=17.425 $Y=1.985
+ $X2=0 $Y2=0
cc_2174 N_D[4]_M1105_g N_A_2839_311#_c_5793_n 0.00232998f $X=17.895 $Y=1.985
+ $X2=0 $Y2=0
cc_2175 N_D[4]_M1042_g N_A_2839_311#_c_5795_n 0.00977623f $X=16.955 $Y=1.985
+ $X2=0 $Y2=0
cc_2176 N_D[4]_M1062_g N_A_2839_311#_c_5795_n 0.00911325f $X=17.425 $Y=1.985
+ $X2=0 $Y2=0
cc_2177 N_D[4]_M1105_g N_A_2839_311#_c_5795_n 7.05028e-19 $X=17.895 $Y=1.985
+ $X2=0 $Y2=0
cc_2178 N_D[4]_M1062_g N_A_2839_311#_c_5798_n 7.05028e-19 $X=17.425 $Y=1.985
+ $X2=0 $Y2=0
cc_2179 N_D[4]_M1105_g N_A_2839_311#_c_5798_n 0.00911325f $X=17.895 $Y=1.985
+ $X2=0 $Y2=0
cc_2180 N_D[4]_M1127_g N_A_2839_311#_c_5798_n 0.00819194f $X=18.365 $Y=1.985
+ $X2=0 $Y2=0
cc_2181 N_D[4]_M1042_g N_A_2839_311#_c_5763_n 0.00333758f $X=16.955 $Y=1.985
+ $X2=0 $Y2=0
cc_2182 N_D[4]_M1027_g N_VGND_c_6290_n 0.00321269f $X=16.98 $Y=0.56 $X2=0 $Y2=0
cc_2183 N_D[4]_M1034_g N_VGND_c_6290_n 2.6376e-19 $X=17.4 $Y=0.56 $X2=0 $Y2=0
cc_2184 N_D[4]_M1034_g N_VGND_c_6292_n 0.0019152f $X=17.4 $Y=0.56 $X2=0 $Y2=0
cc_2185 N_D[4]_M1045_g N_VGND_c_6292_n 0.00166854f $X=17.92 $Y=0.56 $X2=0 $Y2=0
cc_2186 N_D[4]_M1079_g N_VGND_c_6292_n 2.64031e-19 $X=18.34 $Y=0.56 $X2=0 $Y2=0
cc_2187 N_D[4]_M1079_g N_VGND_c_6294_n 0.0058918f $X=18.34 $Y=0.56 $X2=0 $Y2=0
cc_2188 N_D[4]_M1027_g N_VGND_c_6346_n 0.00422241f $X=16.98 $Y=0.56 $X2=0 $Y2=0
cc_2189 N_D[4]_M1034_g N_VGND_c_6346_n 0.00430643f $X=17.4 $Y=0.56 $X2=0 $Y2=0
cc_2190 N_D[4]_M1045_g N_VGND_c_6348_n 0.00422241f $X=17.92 $Y=0.56 $X2=0 $Y2=0
cc_2191 N_D[4]_M1079_g N_VGND_c_6348_n 0.00551064f $X=18.34 $Y=0.56 $X2=0 $Y2=0
cc_2192 N_D[4]_M1027_g N_VGND_c_6370_n 0.00702263f $X=16.98 $Y=0.56 $X2=0 $Y2=0
cc_2193 N_D[4]_M1034_g N_VGND_c_6370_n 0.00624811f $X=17.4 $Y=0.56 $X2=0 $Y2=0
cc_2194 N_D[4]_M1045_g N_VGND_c_6370_n 0.00593887f $X=17.92 $Y=0.56 $X2=0 $Y2=0
cc_2195 N_D[4]_M1079_g N_VGND_c_6370_n 0.0101978f $X=18.34 $Y=0.56 $X2=0 $Y2=0
cc_2196 N_D[4]_M1027_g N_A_2889_66#_c_7258_n 0.00261078f $X=16.98 $Y=0.56 $X2=0
+ $Y2=0
cc_2197 N_D[4]_M1027_g N_A_2889_66#_c_7259_n 0.0121912f $X=16.98 $Y=0.56 $X2=0
+ $Y2=0
cc_2198 N_D[4]_M1027_g N_A_2889_66#_c_7279_n 0.00699463f $X=16.98 $Y=0.56 $X2=0
+ $Y2=0
cc_2199 N_D[4]_M1034_g N_A_2889_66#_c_7279_n 0.00661764f $X=17.4 $Y=0.56 $X2=0
+ $Y2=0
cc_2200 N_D[4]_M1045_g N_A_2889_66#_c_7279_n 5.22365e-19 $X=17.92 $Y=0.56 $X2=0
+ $Y2=0
cc_2201 N_D[4]_M1034_g N_A_2889_66#_c_7261_n 0.00900364f $X=17.4 $Y=0.56 $X2=0
+ $Y2=0
cc_2202 N_D[4]_M1045_g N_A_2889_66#_c_7261_n 0.00986515f $X=17.92 $Y=0.56 $X2=0
+ $Y2=0
cc_2203 N_D[4]_M1079_g N_A_2889_66#_c_7261_n 0.00222549f $X=18.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2204 N_D[4]_c_2738_n N_A_2889_66#_c_7261_n 0.00463549f $X=17.805 $Y=1.16
+ $X2=0 $Y2=0
cc_2205 N_D[4]_c_2740_n N_A_2889_66#_c_7261_n 0.0608884f $X=18.26 $Y=1.16 $X2=0
+ $Y2=0
cc_2206 N_D[4]_c_2741_n N_A_2889_66#_c_7261_n 0.00208088f $X=18.365 $Y=1.16
+ $X2=0 $Y2=0
cc_2207 N_D[4]_M1034_g N_A_2889_66#_c_7288_n 5.22365e-19 $X=17.4 $Y=0.56 $X2=0
+ $Y2=0
cc_2208 N_D[4]_M1045_g N_A_2889_66#_c_7288_n 0.00661134f $X=17.92 $Y=0.56 $X2=0
+ $Y2=0
cc_2209 N_D[4]_M1079_g N_A_2889_66#_c_7288_n 0.00514241f $X=18.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2210 N_D[4]_M1027_g N_A_2889_66#_c_7262_n 0.00128201f $X=16.98 $Y=0.56 $X2=0
+ $Y2=0
cc_2211 N_D[4]_M1034_g N_A_2889_66#_c_7262_n 8.68782e-19 $X=17.4 $Y=0.56 $X2=0
+ $Y2=0
cc_2212 N_D[4]_c_2739_n N_A_2889_66#_c_7262_n 0.00208088f $X=17.515 $Y=1.16
+ $X2=0 $Y2=0
cc_2213 N_D[4]_c_2740_n N_A_2889_66#_c_7262_n 0.018367f $X=18.26 $Y=1.16 $X2=0
+ $Y2=0
cc_2214 N_D[5]_M1134_g N_D[7]_M1087_g 0.0129367f $X=18.365 $Y=3.455 $X2=0 $Y2=0
cc_2215 N_D[5]_M1107_g N_D[7]_M1014_g 0.0210205f $X=18.34 $Y=4.88 $X2=0 $Y2=0
cc_2216 N_D[5]_c_2839_n N_D[7]_c_3036_n 2.99666e-19 $X=18.26 $Y=4.28 $X2=0 $Y2=0
cc_2217 N_D[5]_c_2840_n N_D[7]_c_3036_n 0.0105491f $X=18.365 $Y=4.28 $X2=0 $Y2=0
cc_2218 N_D[5]_c_2839_n N_D[7]_c_3037_n 0.0135469f $X=18.26 $Y=4.28 $X2=0 $Y2=0
cc_2219 N_D[5]_c_2840_n N_D[7]_c_3037_n 2.99666e-19 $X=18.365 $Y=4.28 $X2=0
+ $Y2=0
cc_2220 N_D[5]_M1046_g N_VPWR_c_3611_n 0.00389633f $X=16.955 $Y=3.455 $X2=0
+ $Y2=0
cc_2221 N_D[5]_M1070_g N_VPWR_c_3613_n 0.00208662f $X=17.425 $Y=3.455 $X2=0
+ $Y2=0
cc_2222 N_D[5]_M1113_g N_VPWR_c_3613_n 0.00208662f $X=17.895 $Y=3.455 $X2=0
+ $Y2=0
cc_2223 N_D[5]_M1134_g N_VPWR_c_3615_n 0.00207065f $X=18.365 $Y=3.455 $X2=0
+ $Y2=0
cc_2224 N_D[5]_M1046_g N_VPWR_c_3645_n 0.0035837f $X=16.955 $Y=3.455 $X2=0 $Y2=0
cc_2225 N_D[5]_M1070_g N_VPWR_c_3645_n 0.0035837f $X=17.425 $Y=3.455 $X2=0 $Y2=0
cc_2226 N_D[5]_M1113_g N_VPWR_c_3646_n 0.0035837f $X=17.895 $Y=3.455 $X2=0 $Y2=0
cc_2227 N_D[5]_M1134_g N_VPWR_c_3646_n 0.0035837f $X=18.365 $Y=3.455 $X2=0 $Y2=0
cc_2228 N_D[5]_M1046_g N_VPWR_c_3661_n 0.00573859f $X=16.955 $Y=3.455 $X2=0
+ $Y2=0
cc_2229 N_D[5]_M1070_g N_VPWR_c_3661_n 0.00445624f $X=17.425 $Y=3.455 $X2=0
+ $Y2=0
cc_2230 N_D[5]_M1113_g N_VPWR_c_3661_n 0.00445624f $X=17.895 $Y=3.455 $X2=0
+ $Y2=0
cc_2231 N_D[5]_M1134_g N_VPWR_c_3661_n 0.00579371f $X=18.365 $Y=3.455 $X2=0
+ $Y2=0
cc_2232 N_D[5]_M1046_g N_Z_c_4649_n 0.00311896f $X=16.955 $Y=3.455 $X2=0 $Y2=0
cc_2233 N_D[5]_M1070_g N_Z_c_4649_n 0.00306964f $X=17.425 $Y=3.455 $X2=0 $Y2=0
cc_2234 N_D[5]_M1113_g N_Z_c_4649_n 0.00306964f $X=17.895 $Y=3.455 $X2=0 $Y2=0
cc_2235 N_D[5]_M1134_g N_Z_c_4649_n 0.00470782f $X=18.365 $Y=3.455 $X2=0 $Y2=0
cc_2236 N_D[5]_c_2839_n N_Z_c_4649_n 0.00846955f $X=18.26 $Y=4.28 $X2=0 $Y2=0
cc_2237 N_D[5]_M1046_g N_A_2839_613#_c_5889_n 0.013247f $X=16.955 $Y=3.455 $X2=0
+ $Y2=0
cc_2238 N_D[5]_M1070_g N_A_2839_613#_c_5911_n 0.00916655f $X=17.425 $Y=3.455
+ $X2=0 $Y2=0
cc_2239 N_D[5]_M1113_g N_A_2839_613#_c_5911_n 0.00916655f $X=17.895 $Y=3.455
+ $X2=0 $Y2=0
cc_2240 N_D[5]_c_2837_n N_A_2839_613#_c_5911_n 7.15862e-19 $X=17.805 $Y=4.28
+ $X2=0 $Y2=0
cc_2241 N_D[5]_c_2839_n N_A_2839_613#_c_5911_n 0.0387168f $X=18.26 $Y=4.28 $X2=0
+ $Y2=0
cc_2242 N_D[5]_M1046_g N_A_2839_613#_c_5915_n 8.61029e-19 $X=16.955 $Y=3.455
+ $X2=0 $Y2=0
cc_2243 N_D[5]_M1070_g N_A_2839_613#_c_5915_n 5.79575e-19 $X=17.425 $Y=3.455
+ $X2=0 $Y2=0
cc_2244 N_D[5]_c_2838_n N_A_2839_613#_c_5915_n 8.03631e-19 $X=17.515 $Y=4.28
+ $X2=0 $Y2=0
cc_2245 N_D[5]_c_2839_n N_A_2839_613#_c_5915_n 0.0191156f $X=18.26 $Y=4.28 $X2=0
+ $Y2=0
cc_2246 N_D[5]_M1113_g N_A_2839_613#_c_5919_n 5.79575e-19 $X=17.895 $Y=3.455
+ $X2=0 $Y2=0
cc_2247 N_D[5]_M1134_g N_A_2839_613#_c_5919_n 0.002088f $X=18.365 $Y=3.455 $X2=0
+ $Y2=0
cc_2248 N_D[5]_c_2839_n N_A_2839_613#_c_5919_n 0.0217153f $X=18.26 $Y=4.28 $X2=0
+ $Y2=0
cc_2249 N_D[5]_c_2840_n N_A_2839_613#_c_5919_n 8.03631e-19 $X=18.365 $Y=4.28
+ $X2=0 $Y2=0
cc_2250 N_D[5]_M1046_g N_A_2839_613#_c_5891_n 0.00232998f $X=16.955 $Y=3.455
+ $X2=0 $Y2=0
cc_2251 N_D[5]_M1070_g N_A_2839_613#_c_5924_n 0.00232998f $X=17.425 $Y=3.455
+ $X2=0 $Y2=0
cc_2252 N_D[5]_M1113_g N_A_2839_613#_c_5924_n 0.00232998f $X=17.895 $Y=3.455
+ $X2=0 $Y2=0
cc_2253 N_D[5]_M1046_g N_A_2839_613#_c_5894_n 0.00333758f $X=16.955 $Y=3.455
+ $X2=0 $Y2=0
cc_2254 N_D[5]_M1046_g N_A_2839_613#_c_5927_n 0.00977623f $X=16.955 $Y=3.455
+ $X2=0 $Y2=0
cc_2255 N_D[5]_M1070_g N_A_2839_613#_c_5927_n 0.00911325f $X=17.425 $Y=3.455
+ $X2=0 $Y2=0
cc_2256 N_D[5]_M1113_g N_A_2839_613#_c_5927_n 7.05028e-19 $X=17.895 $Y=3.455
+ $X2=0 $Y2=0
cc_2257 N_D[5]_M1070_g N_A_2839_613#_c_5930_n 7.05028e-19 $X=17.425 $Y=3.455
+ $X2=0 $Y2=0
cc_2258 N_D[5]_M1113_g N_A_2839_613#_c_5930_n 0.00911325f $X=17.895 $Y=3.455
+ $X2=0 $Y2=0
cc_2259 N_D[5]_M1134_g N_A_2839_613#_c_5930_n 0.00819194f $X=18.365 $Y=3.455
+ $X2=0 $Y2=0
cc_2260 N_D[5]_M1033_g N_VGND_c_6291_n 0.00321269f $X=16.98 $Y=4.88 $X2=0 $Y2=0
cc_2261 N_D[5]_M1077_g N_VGND_c_6291_n 2.6376e-19 $X=17.4 $Y=4.88 $X2=0 $Y2=0
cc_2262 N_D[5]_M1077_g N_VGND_c_6293_n 0.0019152f $X=17.4 $Y=4.88 $X2=0 $Y2=0
cc_2263 N_D[5]_M1106_g N_VGND_c_6293_n 0.00166854f $X=17.92 $Y=4.88 $X2=0 $Y2=0
cc_2264 N_D[5]_M1107_g N_VGND_c_6293_n 2.64031e-19 $X=18.34 $Y=4.88 $X2=0 $Y2=0
cc_2265 N_D[5]_M1107_g N_VGND_c_6295_n 0.0058918f $X=18.34 $Y=4.88 $X2=0 $Y2=0
cc_2266 N_D[5]_M1033_g N_VGND_c_6347_n 0.00422241f $X=16.98 $Y=4.88 $X2=0 $Y2=0
cc_2267 N_D[5]_M1077_g N_VGND_c_6347_n 0.00430643f $X=17.4 $Y=4.88 $X2=0 $Y2=0
cc_2268 N_D[5]_M1106_g N_VGND_c_6349_n 0.00422241f $X=17.92 $Y=4.88 $X2=0 $Y2=0
cc_2269 N_D[5]_M1107_g N_VGND_c_6349_n 0.00551064f $X=18.34 $Y=4.88 $X2=0 $Y2=0
cc_2270 N_D[5]_M1033_g N_VGND_c_6371_n 0.00702263f $X=16.98 $Y=4.88 $X2=0 $Y2=0
cc_2271 N_D[5]_M1077_g N_VGND_c_6371_n 0.00624811f $X=17.4 $Y=4.88 $X2=0 $Y2=0
cc_2272 N_D[5]_M1106_g N_VGND_c_6371_n 0.00593887f $X=17.92 $Y=4.88 $X2=0 $Y2=0
cc_2273 N_D[5]_M1107_g N_VGND_c_6371_n 0.0101978f $X=18.34 $Y=4.88 $X2=0 $Y2=0
cc_2274 N_D[5]_M1033_g N_A_2889_918#_c_7342_n 0.00261078f $X=16.98 $Y=4.88 $X2=0
+ $Y2=0
cc_2275 N_D[5]_M1033_g N_A_2889_918#_c_7343_n 0.0121912f $X=16.98 $Y=4.88 $X2=0
+ $Y2=0
cc_2276 N_D[5]_M1077_g N_A_2889_918#_c_7363_n 0.00900364f $X=17.4 $Y=4.88 $X2=0
+ $Y2=0
cc_2277 N_D[5]_M1106_g N_A_2889_918#_c_7363_n 0.00899636f $X=17.92 $Y=4.88 $X2=0
+ $Y2=0
cc_2278 N_D[5]_c_2837_n N_A_2889_918#_c_7363_n 0.00463549f $X=17.805 $Y=4.28
+ $X2=0 $Y2=0
cc_2279 N_D[5]_c_2839_n N_A_2889_918#_c_7363_n 0.0394855f $X=18.26 $Y=4.28 $X2=0
+ $Y2=0
cc_2280 N_D[5]_M1033_g N_A_2889_918#_c_7345_n 0.00827664f $X=16.98 $Y=4.88 $X2=0
+ $Y2=0
cc_2281 N_D[5]_M1077_g N_A_2889_918#_c_7345_n 0.00748643f $X=17.4 $Y=4.88 $X2=0
+ $Y2=0
cc_2282 N_D[5]_M1106_g N_A_2889_918#_c_7345_n 5.22365e-19 $X=17.92 $Y=4.88 $X2=0
+ $Y2=0
cc_2283 N_D[5]_c_2838_n N_A_2889_918#_c_7345_n 0.00208088f $X=17.515 $Y=4.28
+ $X2=0 $Y2=0
cc_2284 N_D[5]_c_2839_n N_A_2889_918#_c_7345_n 0.018367f $X=18.26 $Y=4.28 $X2=0
+ $Y2=0
cc_2285 N_D[5]_M1077_g N_A_2889_918#_c_7346_n 5.22365e-19 $X=17.4 $Y=4.88 $X2=0
+ $Y2=0
cc_2286 N_D[5]_M1106_g N_A_2889_918#_c_7346_n 0.00748012f $X=17.92 $Y=4.88 $X2=0
+ $Y2=0
cc_2287 N_D[5]_M1107_g N_A_2889_918#_c_7346_n 0.0073679f $X=18.34 $Y=4.88 $X2=0
+ $Y2=0
cc_2288 N_D[5]_c_2839_n N_A_2889_918#_c_7346_n 0.021403f $X=18.26 $Y=4.28 $X2=0
+ $Y2=0
cc_2289 N_D[5]_c_2840_n N_A_2889_918#_c_7346_n 0.00208088f $X=18.365 $Y=4.28
+ $X2=0 $Y2=0
cc_2290 N_D[6]_M1082_g N_D[7]_M1087_g 0.0130744f $X=18.895 $Y=1.985 $X2=0 $Y2=0
cc_2291 N_D[6]_M1108_g N_D[7]_M1117_g 0.0130744f $X=19.365 $Y=1.985 $X2=0 $Y2=0
cc_2292 N_D[6]_M1130_g N_D[7]_M1139_g 0.0130744f $X=19.835 $Y=1.985 $X2=0 $Y2=0
cc_2293 N_D[6]_M1145_g N_D[7]_M1153_g 0.0130744f $X=20.305 $Y=1.985 $X2=0 $Y2=0
cc_2294 N_D[6]_M1082_g N_VPWR_c_3614_n 0.00207065f $X=18.895 $Y=1.985 $X2=0
+ $Y2=0
cc_2295 N_D[6]_M1108_g N_VPWR_c_3616_n 0.00208662f $X=19.365 $Y=1.985 $X2=0
+ $Y2=0
cc_2296 N_D[6]_M1130_g N_VPWR_c_3616_n 0.00208662f $X=19.835 $Y=1.985 $X2=0
+ $Y2=0
cc_2297 N_D[6]_M1130_g N_VPWR_c_3618_n 0.0035837f $X=19.835 $Y=1.985 $X2=0 $Y2=0
cc_2298 N_D[6]_M1145_g N_VPWR_c_3618_n 0.0035837f $X=20.305 $Y=1.985 $X2=0 $Y2=0
cc_2299 N_D[6]_M1145_g N_VPWR_c_3619_n 0.00389633f $X=20.305 $Y=1.985 $X2=0
+ $Y2=0
cc_2300 N_D[6]_M1082_g N_VPWR_c_3647_n 0.0035837f $X=18.895 $Y=1.985 $X2=0 $Y2=0
cc_2301 N_D[6]_M1108_g N_VPWR_c_3647_n 0.0035837f $X=19.365 $Y=1.985 $X2=0 $Y2=0
cc_2302 N_D[6]_M1082_g N_VPWR_c_3661_n 0.00579371f $X=18.895 $Y=1.985 $X2=0
+ $Y2=0
cc_2303 N_D[6]_M1108_g N_VPWR_c_3661_n 0.00445624f $X=19.365 $Y=1.985 $X2=0
+ $Y2=0
cc_2304 N_D[6]_M1130_g N_VPWR_c_3661_n 0.00445624f $X=19.835 $Y=1.985 $X2=0
+ $Y2=0
cc_2305 N_D[6]_M1145_g N_VPWR_c_3661_n 0.00573859f $X=20.305 $Y=1.985 $X2=0
+ $Y2=0
cc_2306 N_D[6]_M1082_g N_Z_c_4648_n 0.00470782f $X=18.895 $Y=1.985 $X2=0 $Y2=0
cc_2307 N_D[6]_M1108_g N_Z_c_4648_n 0.00306964f $X=19.365 $Y=1.985 $X2=0 $Y2=0
cc_2308 N_D[6]_M1130_g N_Z_c_4648_n 0.00306964f $X=19.835 $Y=1.985 $X2=0 $Y2=0
cc_2309 N_D[6]_M1145_g N_Z_c_4648_n 0.00311896f $X=20.305 $Y=1.985 $X2=0 $Y2=0
cc_2310 N_D[6]_c_2936_n N_Z_c_4648_n 0.00846955f $X=20.02 $Y=1.16 $X2=0 $Y2=0
cc_2311 N_D[6]_M1108_g N_A_3797_297#_c_6025_n 0.00916655f $X=19.365 $Y=1.985
+ $X2=0 $Y2=0
cc_2312 N_D[6]_M1130_g N_A_3797_297#_c_6025_n 0.00916655f $X=19.835 $Y=1.985
+ $X2=0 $Y2=0
cc_2313 N_D[6]_c_2934_n N_A_3797_297#_c_6025_n 7.15862e-19 $X=19.745 $Y=1.16
+ $X2=0 $Y2=0
cc_2314 N_D[6]_c_2936_n N_A_3797_297#_c_6025_n 0.0387168f $X=20.02 $Y=1.16 $X2=0
+ $Y2=0
cc_2315 N_D[6]_M1145_g N_A_3797_297#_c_6020_n 0.013247f $X=20.305 $Y=1.985 $X2=0
+ $Y2=0
cc_2316 N_D[6]_M1082_g N_A_3797_297#_c_6030_n 0.002088f $X=18.895 $Y=1.985 $X2=0
+ $Y2=0
cc_2317 N_D[6]_M1108_g N_A_3797_297#_c_6030_n 5.79575e-19 $X=19.365 $Y=1.985
+ $X2=0 $Y2=0
cc_2318 N_D[6]_c_2935_n N_A_3797_297#_c_6030_n 8.03631e-19 $X=19.455 $Y=1.16
+ $X2=0 $Y2=0
cc_2319 N_D[6]_c_2936_n N_A_3797_297#_c_6030_n 0.0217153f $X=20.02 $Y=1.16 $X2=0
+ $Y2=0
cc_2320 N_D[6]_M1130_g N_A_3797_297#_c_6034_n 5.79575e-19 $X=19.835 $Y=1.985
+ $X2=0 $Y2=0
cc_2321 N_D[6]_M1145_g N_A_3797_297#_c_6034_n 8.61029e-19 $X=20.305 $Y=1.985
+ $X2=0 $Y2=0
cc_2322 N_D[6]_c_2936_n N_A_3797_297#_c_6034_n 0.0191156f $X=20.02 $Y=1.16 $X2=0
+ $Y2=0
cc_2323 N_D[6]_c_2937_n N_A_3797_297#_c_6034_n 8.03631e-19 $X=20.305 $Y=1.16
+ $X2=0 $Y2=0
cc_2324 N_D[6]_M1108_g N_A_3797_297#_c_6038_n 0.00232998f $X=19.365 $Y=1.985
+ $X2=0 $Y2=0
cc_2325 N_D[6]_M1130_g N_A_3797_297#_c_6038_n 0.00232998f $X=19.835 $Y=1.985
+ $X2=0 $Y2=0
cc_2326 N_D[6]_M1145_g N_A_3797_297#_c_6021_n 0.00232998f $X=20.305 $Y=1.985
+ $X2=0 $Y2=0
cc_2327 N_D[6]_M1082_g N_A_3797_297#_c_6041_n 0.00819194f $X=18.895 $Y=1.985
+ $X2=0 $Y2=0
cc_2328 N_D[6]_M1108_g N_A_3797_297#_c_6041_n 0.00911325f $X=19.365 $Y=1.985
+ $X2=0 $Y2=0
cc_2329 N_D[6]_M1130_g N_A_3797_297#_c_6041_n 7.05028e-19 $X=19.835 $Y=1.985
+ $X2=0 $Y2=0
cc_2330 N_D[6]_M1108_g N_A_3797_297#_c_6044_n 7.05028e-19 $X=19.365 $Y=1.985
+ $X2=0 $Y2=0
cc_2331 N_D[6]_M1130_g N_A_3797_297#_c_6044_n 0.00911325f $X=19.835 $Y=1.985
+ $X2=0 $Y2=0
cc_2332 N_D[6]_M1145_g N_A_3797_297#_c_6044_n 0.00977623f $X=20.305 $Y=1.985
+ $X2=0 $Y2=0
cc_2333 N_D[6]_M1145_g N_A_3797_297#_c_6022_n 0.00333758f $X=20.305 $Y=1.985
+ $X2=0 $Y2=0
cc_2334 N_D[6]_M1005_g N_VGND_c_6294_n 0.0058918f $X=18.92 $Y=0.56 $X2=0 $Y2=0
cc_2335 N_D[6]_M1005_g N_VGND_c_6296_n 2.64031e-19 $X=18.92 $Y=0.56 $X2=0 $Y2=0
cc_2336 N_D[6]_M1081_g N_VGND_c_6296_n 0.00166854f $X=19.34 $Y=0.56 $X2=0 $Y2=0
cc_2337 N_D[6]_M1111_g N_VGND_c_6296_n 0.0019152f $X=19.86 $Y=0.56 $X2=0 $Y2=0
cc_2338 N_D[6]_M1111_g N_VGND_c_6298_n 0.00430643f $X=19.86 $Y=0.56 $X2=0 $Y2=0
cc_2339 N_D[6]_M1159_g N_VGND_c_6298_n 0.00422241f $X=20.28 $Y=0.56 $X2=0 $Y2=0
cc_2340 N_D[6]_M1111_g N_VGND_c_6300_n 2.6376e-19 $X=19.86 $Y=0.56 $X2=0 $Y2=0
cc_2341 N_D[6]_M1159_g N_VGND_c_6300_n 0.00321269f $X=20.28 $Y=0.56 $X2=0 $Y2=0
cc_2342 N_D[6]_M1005_g N_VGND_c_6350_n 0.00551064f $X=18.92 $Y=0.56 $X2=0 $Y2=0
cc_2343 N_D[6]_M1081_g N_VGND_c_6350_n 0.00422241f $X=19.34 $Y=0.56 $X2=0 $Y2=0
cc_2344 N_D[6]_M1005_g N_VGND_c_6370_n 0.0101978f $X=18.92 $Y=0.56 $X2=0 $Y2=0
cc_2345 N_D[6]_M1081_g N_VGND_c_6370_n 0.00593887f $X=19.34 $Y=0.56 $X2=0 $Y2=0
cc_2346 N_D[6]_M1111_g N_VGND_c_6370_n 0.00624811f $X=19.86 $Y=0.56 $X2=0 $Y2=0
cc_2347 N_D[6]_M1159_g N_VGND_c_6370_n 0.00702263f $X=20.28 $Y=0.56 $X2=0 $Y2=0
cc_2348 N_D[6]_M1005_g N_A_3799_47#_c_7428_n 0.00514241f $X=18.92 $Y=0.56 $X2=0
+ $Y2=0
cc_2349 N_D[6]_M1081_g N_A_3799_47#_c_7428_n 0.00661134f $X=19.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2350 N_D[6]_M1111_g N_A_3799_47#_c_7428_n 5.22365e-19 $X=19.86 $Y=0.56 $X2=0
+ $Y2=0
cc_2351 N_D[6]_M1081_g N_A_3799_47#_c_7431_n 0.00899636f $X=19.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2352 N_D[6]_M1111_g N_A_3799_47#_c_7431_n 0.00900364f $X=19.86 $Y=0.56 $X2=0
+ $Y2=0
cc_2353 N_D[6]_c_2934_n N_A_3799_47#_c_7431_n 0.00463549f $X=19.745 $Y=1.16
+ $X2=0 $Y2=0
cc_2354 N_D[6]_c_2936_n N_A_3799_47#_c_7431_n 0.0394855f $X=20.02 $Y=1.16 $X2=0
+ $Y2=0
cc_2355 N_D[6]_M1005_g N_A_3799_47#_c_7420_n 0.00222549f $X=18.92 $Y=0.56 $X2=0
+ $Y2=0
cc_2356 N_D[6]_M1081_g N_A_3799_47#_c_7420_n 8.68782e-19 $X=19.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2357 N_D[6]_c_2935_n N_A_3799_47#_c_7420_n 0.00208088f $X=19.455 $Y=1.16
+ $X2=0 $Y2=0
cc_2358 N_D[6]_c_2936_n N_A_3799_47#_c_7420_n 0.021403f $X=20.02 $Y=1.16 $X2=0
+ $Y2=0
cc_2359 N_D[6]_M1081_g N_A_3799_47#_c_7439_n 5.22365e-19 $X=19.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2360 N_D[6]_M1111_g N_A_3799_47#_c_7439_n 0.00661764f $X=19.86 $Y=0.56 $X2=0
+ $Y2=0
cc_2361 N_D[6]_M1159_g N_A_3799_47#_c_7439_n 0.00699463f $X=20.28 $Y=0.56 $X2=0
+ $Y2=0
cc_2362 N_D[6]_M1159_g N_A_3799_47#_c_7421_n 0.0121912f $X=20.28 $Y=0.56 $X2=0
+ $Y2=0
cc_2363 N_D[6]_M1159_g N_A_3799_47#_c_7422_n 0.00261078f $X=20.28 $Y=0.56 $X2=0
+ $Y2=0
cc_2364 N_D[6]_M1111_g N_A_3799_47#_c_7427_n 8.68782e-19 $X=19.86 $Y=0.56 $X2=0
+ $Y2=0
cc_2365 N_D[6]_M1159_g N_A_3799_47#_c_7427_n 0.00128201f $X=20.28 $Y=0.56 $X2=0
+ $Y2=0
cc_2366 N_D[6]_c_2936_n N_A_3799_47#_c_7427_n 0.018367f $X=20.02 $Y=1.16 $X2=0
+ $Y2=0
cc_2367 N_D[6]_c_2937_n N_A_3799_47#_c_7427_n 0.00208088f $X=20.305 $Y=1.16
+ $X2=0 $Y2=0
cc_2368 N_D[7]_M1087_g N_VPWR_c_3615_n 0.00207065f $X=18.895 $Y=3.455 $X2=0
+ $Y2=0
cc_2369 N_D[7]_M1117_g N_VPWR_c_3617_n 0.00208662f $X=19.365 $Y=3.455 $X2=0
+ $Y2=0
cc_2370 N_D[7]_M1139_g N_VPWR_c_3617_n 0.00208662f $X=19.835 $Y=3.455 $X2=0
+ $Y2=0
cc_2371 N_D[7]_M1139_g N_VPWR_c_3618_n 0.0035837f $X=19.835 $Y=3.455 $X2=0 $Y2=0
cc_2372 N_D[7]_M1153_g N_VPWR_c_3618_n 0.0035837f $X=20.305 $Y=3.455 $X2=0 $Y2=0
cc_2373 N_D[7]_M1153_g N_VPWR_c_3620_n 0.00389633f $X=20.305 $Y=3.455 $X2=0
+ $Y2=0
cc_2374 N_D[7]_M1087_g N_VPWR_c_3647_n 0.0035837f $X=18.895 $Y=3.455 $X2=0 $Y2=0
cc_2375 N_D[7]_M1117_g N_VPWR_c_3647_n 0.0035837f $X=19.365 $Y=3.455 $X2=0 $Y2=0
cc_2376 N_D[7]_M1087_g N_VPWR_c_3661_n 0.00579371f $X=18.895 $Y=3.455 $X2=0
+ $Y2=0
cc_2377 N_D[7]_M1117_g N_VPWR_c_3661_n 0.00445624f $X=19.365 $Y=3.455 $X2=0
+ $Y2=0
cc_2378 N_D[7]_M1139_g N_VPWR_c_3661_n 0.00445624f $X=19.835 $Y=3.455 $X2=0
+ $Y2=0
cc_2379 N_D[7]_M1153_g N_VPWR_c_3661_n 0.00573859f $X=20.305 $Y=3.455 $X2=0
+ $Y2=0
cc_2380 N_D[7]_M1087_g N_Z_c_4649_n 0.00470782f $X=18.895 $Y=3.455 $X2=0 $Y2=0
cc_2381 N_D[7]_M1117_g N_Z_c_4649_n 0.00306964f $X=19.365 $Y=3.455 $X2=0 $Y2=0
cc_2382 N_D[7]_M1139_g N_Z_c_4649_n 0.00306964f $X=19.835 $Y=3.455 $X2=0 $Y2=0
cc_2383 N_D[7]_M1153_g N_Z_c_4649_n 0.00311896f $X=20.305 $Y=3.455 $X2=0 $Y2=0
cc_2384 N_D[7]_c_3037_n N_Z_c_4649_n 0.00846955f $X=20.02 $Y=4.28 $X2=0 $Y2=0
cc_2385 N_D[7]_M1117_g N_A_3797_591#_c_6147_n 0.00916655f $X=19.365 $Y=3.455
+ $X2=0 $Y2=0
cc_2386 N_D[7]_M1139_g N_A_3797_591#_c_6147_n 0.00916655f $X=19.835 $Y=3.455
+ $X2=0 $Y2=0
cc_2387 N_D[7]_c_3035_n N_A_3797_591#_c_6147_n 7.15862e-19 $X=19.745 $Y=4.28
+ $X2=0 $Y2=0
cc_2388 N_D[7]_c_3037_n N_A_3797_591#_c_6147_n 0.0387168f $X=20.02 $Y=4.28 $X2=0
+ $Y2=0
cc_2389 N_D[7]_M1153_g N_A_3797_591#_c_6142_n 0.013247f $X=20.305 $Y=3.455 $X2=0
+ $Y2=0
cc_2390 N_D[7]_M1087_g N_A_3797_591#_c_6152_n 0.002088f $X=18.895 $Y=3.455 $X2=0
+ $Y2=0
cc_2391 N_D[7]_M1117_g N_A_3797_591#_c_6152_n 5.79575e-19 $X=19.365 $Y=3.455
+ $X2=0 $Y2=0
cc_2392 N_D[7]_c_3036_n N_A_3797_591#_c_6152_n 8.03631e-19 $X=19.455 $Y=4.28
+ $X2=0 $Y2=0
cc_2393 N_D[7]_c_3037_n N_A_3797_591#_c_6152_n 0.0217153f $X=20.02 $Y=4.28 $X2=0
+ $Y2=0
cc_2394 N_D[7]_M1139_g N_A_3797_591#_c_6156_n 5.79575e-19 $X=19.835 $Y=3.455
+ $X2=0 $Y2=0
cc_2395 N_D[7]_M1153_g N_A_3797_591#_c_6156_n 8.61029e-19 $X=20.305 $Y=3.455
+ $X2=0 $Y2=0
cc_2396 N_D[7]_c_3037_n N_A_3797_591#_c_6156_n 0.0191156f $X=20.02 $Y=4.28 $X2=0
+ $Y2=0
cc_2397 N_D[7]_c_3038_n N_A_3797_591#_c_6156_n 8.03631e-19 $X=20.305 $Y=4.28
+ $X2=0 $Y2=0
cc_2398 N_D[7]_M1117_g N_A_3797_591#_c_6160_n 0.00232998f $X=19.365 $Y=3.455
+ $X2=0 $Y2=0
cc_2399 N_D[7]_M1139_g N_A_3797_591#_c_6160_n 0.00232998f $X=19.835 $Y=3.455
+ $X2=0 $Y2=0
cc_2400 N_D[7]_M1153_g N_A_3797_591#_c_6143_n 0.00232998f $X=20.305 $Y=3.455
+ $X2=0 $Y2=0
cc_2401 N_D[7]_M1087_g N_A_3797_591#_c_6163_n 0.00819194f $X=18.895 $Y=3.455
+ $X2=0 $Y2=0
cc_2402 N_D[7]_M1117_g N_A_3797_591#_c_6163_n 0.00911325f $X=19.365 $Y=3.455
+ $X2=0 $Y2=0
cc_2403 N_D[7]_M1139_g N_A_3797_591#_c_6163_n 7.05028e-19 $X=19.835 $Y=3.455
+ $X2=0 $Y2=0
cc_2404 N_D[7]_M1117_g N_A_3797_591#_c_6166_n 7.05028e-19 $X=19.365 $Y=3.455
+ $X2=0 $Y2=0
cc_2405 N_D[7]_M1139_g N_A_3797_591#_c_6166_n 0.00911325f $X=19.835 $Y=3.455
+ $X2=0 $Y2=0
cc_2406 N_D[7]_M1153_g N_A_3797_591#_c_6166_n 0.00977623f $X=20.305 $Y=3.455
+ $X2=0 $Y2=0
cc_2407 N_D[7]_M1153_g N_A_3797_591#_c_6144_n 0.00333758f $X=20.305 $Y=3.455
+ $X2=0 $Y2=0
cc_2408 N_D[7]_M1014_g N_VGND_c_6295_n 0.0058918f $X=18.92 $Y=4.88 $X2=0 $Y2=0
cc_2409 N_D[7]_M1014_g N_VGND_c_6297_n 2.64031e-19 $X=18.92 $Y=4.88 $X2=0 $Y2=0
cc_2410 N_D[7]_M1025_g N_VGND_c_6297_n 0.00166854f $X=19.34 $Y=4.88 $X2=0 $Y2=0
cc_2411 N_D[7]_M1026_g N_VGND_c_6297_n 0.0019152f $X=19.86 $Y=4.88 $X2=0 $Y2=0
cc_2412 N_D[7]_M1026_g N_VGND_c_6299_n 0.00430643f $X=19.86 $Y=4.88 $X2=0 $Y2=0
cc_2413 N_D[7]_M1098_g N_VGND_c_6299_n 0.00422241f $X=20.28 $Y=4.88 $X2=0 $Y2=0
cc_2414 N_D[7]_M1026_g N_VGND_c_6301_n 2.6376e-19 $X=19.86 $Y=4.88 $X2=0 $Y2=0
cc_2415 N_D[7]_M1098_g N_VGND_c_6301_n 0.00321269f $X=20.28 $Y=4.88 $X2=0 $Y2=0
cc_2416 N_D[7]_M1014_g N_VGND_c_6351_n 0.00551064f $X=18.92 $Y=4.88 $X2=0 $Y2=0
cc_2417 N_D[7]_M1025_g N_VGND_c_6351_n 0.00422241f $X=19.34 $Y=4.88 $X2=0 $Y2=0
cc_2418 N_D[7]_M1014_g N_VGND_c_6371_n 0.0101978f $X=18.92 $Y=4.88 $X2=0 $Y2=0
cc_2419 N_D[7]_M1025_g N_VGND_c_6371_n 0.00593887f $X=19.34 $Y=4.88 $X2=0 $Y2=0
cc_2420 N_D[7]_M1026_g N_VGND_c_6371_n 0.00624811f $X=19.86 $Y=4.88 $X2=0 $Y2=0
cc_2421 N_D[7]_M1098_g N_VGND_c_6371_n 0.00702263f $X=20.28 $Y=4.88 $X2=0 $Y2=0
cc_2422 N_D[7]_M1025_g N_A_3799_911#_c_7511_n 0.00899636f $X=19.34 $Y=4.88 $X2=0
+ $Y2=0
cc_2423 N_D[7]_M1026_g N_A_3799_911#_c_7511_n 0.00900364f $X=19.86 $Y=4.88 $X2=0
+ $Y2=0
cc_2424 N_D[7]_c_3035_n N_A_3799_911#_c_7511_n 0.00463549f $X=19.745 $Y=4.28
+ $X2=0 $Y2=0
cc_2425 N_D[7]_c_3037_n N_A_3799_911#_c_7511_n 0.0394855f $X=20.02 $Y=4.28 $X2=0
+ $Y2=0
cc_2426 N_D[7]_M1098_g N_A_3799_911#_c_7503_n 0.0121912f $X=20.28 $Y=4.88 $X2=0
+ $Y2=0
cc_2427 N_D[7]_M1098_g N_A_3799_911#_c_7504_n 0.00261078f $X=20.28 $Y=4.88 $X2=0
+ $Y2=0
cc_2428 N_D[7]_M1014_g N_A_3799_911#_c_7509_n 0.0073679f $X=18.92 $Y=4.88 $X2=0
+ $Y2=0
cc_2429 N_D[7]_M1025_g N_A_3799_911#_c_7509_n 0.00748012f $X=19.34 $Y=4.88 $X2=0
+ $Y2=0
cc_2430 N_D[7]_M1026_g N_A_3799_911#_c_7509_n 5.22365e-19 $X=19.86 $Y=4.88 $X2=0
+ $Y2=0
cc_2431 N_D[7]_c_3036_n N_A_3799_911#_c_7509_n 0.00208088f $X=19.455 $Y=4.28
+ $X2=0 $Y2=0
cc_2432 N_D[7]_c_3037_n N_A_3799_911#_c_7509_n 0.021403f $X=20.02 $Y=4.28 $X2=0
+ $Y2=0
cc_2433 N_D[7]_M1025_g N_A_3799_911#_c_7510_n 5.22365e-19 $X=19.34 $Y=4.88 $X2=0
+ $Y2=0
cc_2434 N_D[7]_M1026_g N_A_3799_911#_c_7510_n 0.00748643f $X=19.86 $Y=4.88 $X2=0
+ $Y2=0
cc_2435 N_D[7]_M1098_g N_A_3799_911#_c_7510_n 0.00827664f $X=20.28 $Y=4.88 $X2=0
+ $Y2=0
cc_2436 N_D[7]_c_3037_n N_A_3799_911#_c_7510_n 0.018367f $X=20.02 $Y=4.28 $X2=0
+ $Y2=0
cc_2437 N_D[7]_c_3038_n N_A_3799_911#_c_7510_n 0.00208088f $X=20.305 $Y=4.28
+ $X2=0 $Y2=0
cc_2438 N_A_4239_265#_c_3131_n N_A_4239_793#_c_3246_n 0.0129371f $X=21.295
+ $Y=1.475 $X2=0 $Y2=0
cc_2439 N_A_4239_265#_c_3134_n N_A_4239_793#_c_3249_n 0.0129371f $X=21.765
+ $Y=1.475 $X2=0 $Y2=0
cc_2440 N_A_4239_265#_c_3136_n N_A_4239_793#_c_3251_n 0.0129371f $X=22.235
+ $Y=1.475 $X2=0 $Y2=0
cc_2441 N_A_4239_265#_c_3138_n N_A_4239_793#_c_3253_n 0.0129371f $X=22.705
+ $Y=1.475 $X2=0 $Y2=0
cc_2442 N_A_4239_265#_c_3133_n N_S[6]_c_3360_n 0.00507426f $X=21.385 $Y=1.4
+ $X2=-0.19 $Y2=-0.24
cc_2443 N_A_4239_265#_c_3132_n N_S[6]_c_3363_n 0.00509391f $X=21.675 $Y=1.4
+ $X2=0 $Y2=0
cc_2444 N_A_4239_265#_c_3135_n N_S[6]_c_3365_n 0.00509204f $X=22.145 $Y=1.4
+ $X2=0 $Y2=0
cc_2445 N_A_4239_265#_c_3137_n N_S[6]_c_3367_n 0.00507688f $X=22.615 $Y=1.4
+ $X2=0 $Y2=0
cc_2446 N_A_4239_265#_c_3126_n N_S[6]_c_3369_n 6.53442e-19 $X=23.985 $Y=0.445
+ $X2=0 $Y2=0
cc_2447 N_A_4239_265#_c_3124_n N_S[6]_c_3371_n 0.0103812f $X=23.82 $Y=1.23 $X2=0
+ $Y2=0
cc_2448 N_A_4239_265#_c_3125_n N_S[6]_c_3371_n 0.0179529f $X=23.275 $Y=1.23
+ $X2=0 $Y2=0
cc_2449 N_A_4239_265#_c_3124_n N_S[6]_c_3372_n 0.0250056f $X=23.82 $Y=1.23 $X2=0
+ $Y2=0
cc_2450 N_A_4239_265#_c_3125_n N_S[6]_c_3372_n 0.0175393f $X=23.275 $Y=1.23
+ $X2=0 $Y2=0
cc_2451 N_A_4239_265#_c_3127_n N_S[6]_c_3372_n 0.0085951f $X=23.905 $Y=1.065
+ $X2=0 $Y2=0
cc_2452 N_A_4239_265#_c_3129_n N_S[6]_c_3372_n 0.00322131f $X=23.905 $Y=1.23
+ $X2=0 $Y2=0
cc_2453 N_A_4239_265#_c_3145_n N_S[6]_c_3372_n 0.00255921f $X=23.985 $Y=1.605
+ $X2=0 $Y2=0
cc_2454 N_A_4239_265#_c_3130_n N_S[6]_c_3372_n 0.00262132f $X=23.025 $Y=1.23
+ $X2=0 $Y2=0
cc_2455 N_A_4239_265#_c_3143_n N_S[6]_c_3383_n 0.0123982f $X=23.985 $Y=1.77
+ $X2=0 $Y2=0
cc_2456 N_A_4239_265#_c_3145_n N_S[6]_c_3383_n 0.00762115f $X=23.985 $Y=1.605
+ $X2=0 $Y2=0
cc_2457 N_A_4239_265#_c_3126_n N_S[6]_c_3373_n 0.00603996f $X=23.985 $Y=0.445
+ $X2=0 $Y2=0
cc_2458 N_A_4239_265#_c_3128_n N_S[6]_c_3373_n 9.67113e-19 $X=23.945 $Y=0.825
+ $X2=0 $Y2=0
cc_2459 N_A_4239_265#_c_3127_n N_S[6]_c_3374_n 0.00429801f $X=23.905 $Y=1.065
+ $X2=0 $Y2=0
cc_2460 N_A_4239_265#_c_3128_n N_S[6]_c_3374_n 0.0111895f $X=23.945 $Y=0.825
+ $X2=0 $Y2=0
cc_2461 N_A_4239_265#_c_3126_n N_S[6]_c_3375_n 0.00207203f $X=23.985 $Y=0.445
+ $X2=0 $Y2=0
cc_2462 N_A_4239_265#_c_3127_n N_S[6]_c_3376_n 0.00289358f $X=23.905 $Y=1.065
+ $X2=0 $Y2=0
cc_2463 N_A_4239_265#_c_3143_n N_S[6]_c_3376_n 0.0133753f $X=23.985 $Y=1.77
+ $X2=0 $Y2=0
cc_2464 N_A_4239_265#_c_3129_n N_S[6]_c_3376_n 0.00416423f $X=23.905 $Y=1.23
+ $X2=0 $Y2=0
cc_2465 N_A_4239_265#_c_3145_n N_S[6]_c_3376_n 0.00454075f $X=23.985 $Y=1.605
+ $X2=0 $Y2=0
cc_2466 N_A_4239_265#_c_3127_n N_S[6]_c_3380_n 0.00268644f $X=23.905 $Y=1.065
+ $X2=0 $Y2=0
cc_2467 N_A_4239_265#_c_3128_n N_S[6]_c_3380_n 0.00426435f $X=23.945 $Y=0.825
+ $X2=0 $Y2=0
cc_2468 N_A_4239_265#_c_3127_n S[6] 0.00541767f $X=23.905 $Y=1.065 $X2=0 $Y2=0
cc_2469 N_A_4239_265#_c_3129_n S[6] 0.0228692f $X=23.905 $Y=1.23 $X2=0 $Y2=0
cc_2470 N_A_4239_265#_c_3131_n N_VPWR_c_3619_n 0.00324472f $X=21.295 $Y=1.475
+ $X2=0 $Y2=0
cc_2471 N_A_4239_265#_c_3138_n N_VPWR_c_3621_n 0.00377407f $X=22.705 $Y=1.475
+ $X2=0 $Y2=0
cc_2472 N_A_4239_265#_c_3124_n N_VPWR_c_3621_n 0.0208071f $X=23.82 $Y=1.23 $X2=0
+ $Y2=0
cc_2473 N_A_4239_265#_c_3125_n N_VPWR_c_3621_n 6.4101e-19 $X=23.275 $Y=1.23
+ $X2=0 $Y2=0
cc_2474 N_A_4239_265#_c_3143_n N_VPWR_c_3621_n 0.0302744f $X=23.985 $Y=1.77
+ $X2=0 $Y2=0
cc_2475 N_A_4239_265#_c_3143_n N_VPWR_c_3623_n 0.03379f $X=23.985 $Y=1.77 $X2=0
+ $Y2=0
cc_2476 N_A_4239_265#_c_3143_n N_VPWR_c_3649_n 0.0233824f $X=23.985 $Y=1.77
+ $X2=0 $Y2=0
cc_2477 N_A_4239_265#_c_3131_n N_VPWR_c_3661_n 0.00473731f $X=21.295 $Y=1.475
+ $X2=0 $Y2=0
cc_2478 N_A_4239_265#_c_3134_n N_VPWR_c_3661_n 0.00362156f $X=21.765 $Y=1.475
+ $X2=0 $Y2=0
cc_2479 N_A_4239_265#_c_3136_n N_VPWR_c_3661_n 0.00362156f $X=22.235 $Y=1.475
+ $X2=0 $Y2=0
cc_2480 N_A_4239_265#_c_3138_n N_VPWR_c_3661_n 0.00473731f $X=22.705 $Y=1.475
+ $X2=0 $Y2=0
cc_2481 N_A_4239_265#_c_3143_n N_VPWR_c_3661_n 0.0124581f $X=23.985 $Y=1.77
+ $X2=0 $Y2=0
cc_2482 N_A_4239_265#_c_3135_n N_Z_c_4604_n 0.00762343f $X=22.145 $Y=1.4 $X2=0
+ $Y2=0
cc_2483 N_A_4239_265#_c_3139_n N_Z_c_4604_n 0.00704092f $X=21.765 $Y=1.4 $X2=0
+ $Y2=0
cc_2484 N_A_4239_265#_c_3133_n N_Z_c_4629_n 0.00248496f $X=21.385 $Y=1.4 $X2=0
+ $Y2=0
cc_2485 N_A_4239_265#_c_3132_n N_Z_c_4632_n 0.00678861f $X=21.675 $Y=1.4 $X2=0
+ $Y2=0
cc_2486 N_A_4239_265#_c_3133_n N_Z_c_4632_n 0.00239476f $X=21.385 $Y=1.4 $X2=0
+ $Y2=0
cc_2487 N_A_4239_265#_c_3139_n N_Z_c_4632_n 2.98555e-19 $X=21.765 $Y=1.4 $X2=0
+ $Y2=0
cc_2488 N_A_4239_265#_c_3135_n N_Z_c_4634_n 0.00145542f $X=22.145 $Y=1.4 $X2=0
+ $Y2=0
cc_2489 N_A_4239_265#_c_3137_n N_Z_c_4634_n 0.00597584f $X=22.615 $Y=1.4 $X2=0
+ $Y2=0
cc_2490 N_A_4239_265#_c_3140_n N_Z_c_4634_n 0.00909323f $X=22.235 $Y=1.4 $X2=0
+ $Y2=0
cc_2491 N_A_4239_265#_c_3124_n N_Z_c_4634_n 0.0266078f $X=23.82 $Y=1.23 $X2=0
+ $Y2=0
cc_2492 N_A_4239_265#_c_3130_n N_Z_c_4634_n 0.00747617f $X=23.025 $Y=1.23 $X2=0
+ $Y2=0
cc_2493 N_A_4239_265#_c_3131_n N_Z_c_4648_n 0.00834829f $X=21.295 $Y=1.475 $X2=0
+ $Y2=0
cc_2494 N_A_4239_265#_c_3134_n Z 0.00372458f $X=21.765 $Y=1.475 $X2=0 $Y2=0
cc_2495 N_A_4239_265#_c_3136_n Z 0.00372248f $X=22.235 $Y=1.475 $X2=0 $Y2=0
cc_2496 N_A_4239_265#_c_3131_n N_Z_c_4656_n 0.0199111f $X=21.295 $Y=1.475 $X2=0
+ $Y2=0
cc_2497 N_A_4239_265#_c_3132_n N_Z_c_4656_n 0.00560592f $X=21.675 $Y=1.4 $X2=0
+ $Y2=0
cc_2498 N_A_4239_265#_c_3133_n N_Z_c_4656_n 0.00474497f $X=21.385 $Y=1.4 $X2=0
+ $Y2=0
cc_2499 N_A_4239_265#_c_3134_n N_Z_c_4656_n 0.0181262f $X=21.765 $Y=1.475 $X2=0
+ $Y2=0
cc_2500 N_A_4239_265#_c_3136_n N_Z_c_4656_n 9.74366e-19 $X=22.235 $Y=1.475 $X2=0
+ $Y2=0
cc_2501 N_A_4239_265#_c_3139_n N_Z_c_4656_n 0.00415268f $X=21.765 $Y=1.4 $X2=0
+ $Y2=0
cc_2502 N_A_4239_265#_c_3134_n N_Z_c_4657_n 9.74366e-19 $X=21.765 $Y=1.475 $X2=0
+ $Y2=0
cc_2503 N_A_4239_265#_c_3136_n N_Z_c_4657_n 0.0181262f $X=22.235 $Y=1.475 $X2=0
+ $Y2=0
cc_2504 N_A_4239_265#_c_3137_n N_Z_c_4657_n 0.00560592f $X=22.615 $Y=1.4 $X2=0
+ $Y2=0
cc_2505 N_A_4239_265#_c_3138_n N_Z_c_4657_n 0.0226667f $X=22.705 $Y=1.475 $X2=0
+ $Y2=0
cc_2506 N_A_4239_265#_c_3140_n N_Z_c_4657_n 0.00181273f $X=22.235 $Y=1.4 $X2=0
+ $Y2=0
cc_2507 N_A_4239_265#_c_3124_n N_Z_c_4657_n 0.00240108f $X=23.82 $Y=1.23 $X2=0
+ $Y2=0
cc_2508 N_A_4239_265#_c_3130_n N_Z_c_4657_n 0.00425035f $X=23.025 $Y=1.23 $X2=0
+ $Y2=0
cc_2509 N_A_4239_265#_c_3131_n N_A_3797_297#_c_6020_n 0.00151141f $X=21.295
+ $Y=1.475 $X2=0 $Y2=0
cc_2510 N_A_4239_265#_c_3131_n N_A_3797_297#_c_6049_n 0.00307958f $X=21.295
+ $Y=1.475 $X2=0 $Y2=0
cc_2511 N_A_4239_265#_c_3134_n N_A_3797_297#_c_6049_n 0.00307958f $X=21.765
+ $Y=1.475 $X2=0 $Y2=0
cc_2512 N_A_4239_265#_c_3136_n N_A_3797_297#_c_6051_n 0.00307958f $X=22.235
+ $Y=1.475 $X2=0 $Y2=0
cc_2513 N_A_4239_265#_c_3138_n N_A_3797_297#_c_6051_n 0.00799829f $X=22.705
+ $Y=1.475 $X2=0 $Y2=0
cc_2514 N_A_4239_265#_c_3131_n N_A_3797_297#_c_6022_n 0.00554566f $X=21.295
+ $Y=1.475 $X2=0 $Y2=0
cc_2515 N_A_4239_265#_c_3134_n N_A_3797_297#_c_6023_n 0.00210632f $X=21.765
+ $Y=1.475 $X2=0 $Y2=0
cc_2516 N_A_4239_265#_c_3135_n N_A_3797_297#_c_6023_n 0.00251792f $X=22.145
+ $Y=1.4 $X2=0 $Y2=0
cc_2517 N_A_4239_265#_c_3136_n N_A_3797_297#_c_6023_n 0.00210632f $X=22.235
+ $Y=1.475 $X2=0 $Y2=0
cc_2518 N_A_4239_265#_c_3138_n N_A_3797_297#_c_6024_n 0.00483827f $X=22.705
+ $Y=1.475 $X2=0 $Y2=0
cc_2519 N_A_4239_265#_c_3124_n N_A_3797_297#_c_6024_n 0.0229374f $X=23.82
+ $Y=1.23 $X2=0 $Y2=0
cc_2520 N_A_4239_265#_c_3125_n N_A_3797_297#_c_6024_n 5.74251e-19 $X=23.275
+ $Y=1.23 $X2=0 $Y2=0
cc_2521 N_A_4239_265#_c_3130_n N_A_3797_297#_c_6024_n 0.00561627f $X=23.025
+ $Y=1.23 $X2=0 $Y2=0
cc_2522 N_A_4239_265#_c_3124_n N_VGND_c_6302_n 0.0123065f $X=23.82 $Y=1.23 $X2=0
+ $Y2=0
cc_2523 N_A_4239_265#_c_3125_n N_VGND_c_6302_n 2.04129e-19 $X=23.275 $Y=1.23
+ $X2=0 $Y2=0
cc_2524 N_A_4239_265#_c_3126_n N_VGND_c_6352_n 0.0129994f $X=23.985 $Y=0.445
+ $X2=0 $Y2=0
cc_2525 N_A_4239_265#_M1032_d N_VGND_c_6370_n 0.00394793f $X=23.85 $Y=0.235
+ $X2=0 $Y2=0
cc_2526 N_A_4239_265#_c_3126_n N_VGND_c_6370_n 0.00927134f $X=23.985 $Y=0.445
+ $X2=0 $Y2=0
cc_2527 N_A_4239_265#_c_3139_n N_A_3799_47#_c_7448_n 7.0477e-19 $X=21.765 $Y=1.4
+ $X2=0 $Y2=0
cc_2528 N_A_4239_265#_c_3124_n N_A_3799_47#_c_7426_n 0.0028695f $X=23.82 $Y=1.23
+ $X2=0 $Y2=0
cc_2529 N_A_4239_265#_c_3130_n N_A_3799_47#_c_7426_n 0.00589316f $X=23.025
+ $Y=1.23 $X2=0 $Y2=0
cc_2530 N_A_4239_793#_c_3248_n N_S[7]_c_3470_n 0.00507426f $X=21.385 $Y=4.04
+ $X2=-0.19 $Y2=-0.24
cc_2531 N_A_4239_793#_c_3247_n N_S[7]_c_3473_n 0.00509391f $X=21.675 $Y=4.04
+ $X2=0 $Y2=0
cc_2532 N_A_4239_793#_c_3250_n N_S[7]_c_3475_n 0.00509204f $X=22.145 $Y=4.04
+ $X2=0 $Y2=0
cc_2533 N_A_4239_793#_c_3252_n N_S[7]_c_3477_n 0.00507688f $X=22.615 $Y=4.04
+ $X2=0 $Y2=0
cc_2534 N_A_4239_793#_c_3241_n N_S[7]_c_3479_n 6.53442e-19 $X=23.945 $Y=4.74
+ $X2=0 $Y2=0
cc_2535 N_A_4239_793#_c_3239_n N_S[7]_c_3481_n 0.0103812f $X=23.82 $Y=4.21 $X2=0
+ $Y2=0
cc_2536 N_A_4239_793#_c_3240_n N_S[7]_c_3481_n 0.0179529f $X=23.275 $Y=4.21
+ $X2=0 $Y2=0
cc_2537 N_A_4239_793#_c_3259_n N_S[7]_c_3491_n 0.00508008f $X=23.905 $Y=4.045
+ $X2=0 $Y2=0
cc_2538 N_A_4239_793#_c_3245_n N_S[7]_c_3491_n 0.00262132f $X=23.025 $Y=4.21
+ $X2=0 $Y2=0
cc_2539 N_A_4239_793#_c_3239_n N_S[7]_c_3482_n 0.0250056f $X=23.82 $Y=4.21 $X2=0
+ $Y2=0
cc_2540 N_A_4239_793#_c_3240_n N_S[7]_c_3482_n 0.0175393f $X=23.275 $Y=4.21
+ $X2=0 $Y2=0
cc_2541 N_A_4239_793#_c_3259_n N_S[7]_c_3482_n 0.00255921f $X=23.905 $Y=4.045
+ $X2=0 $Y2=0
cc_2542 N_A_4239_793#_c_3243_n N_S[7]_c_3482_n 0.00322131f $X=23.905 $Y=4.21
+ $X2=0 $Y2=0
cc_2543 N_A_4239_793#_c_3244_n N_S[7]_c_3482_n 0.0085951f $X=23.945 $Y=4.615
+ $X2=0 $Y2=0
cc_2544 N_A_4239_793#_c_3258_n N_S[7]_c_3493_n 0.010234f $X=23.985 $Y=3.14 $X2=0
+ $Y2=0
cc_2545 N_A_4239_793#_c_3259_n N_S[7]_c_3493_n 0.00254107f $X=23.905 $Y=4.045
+ $X2=0 $Y2=0
cc_2546 N_A_4239_793#_c_3260_n N_S[7]_c_3493_n 0.00216424f $X=23.985 $Y=3.835
+ $X2=0 $Y2=0
cc_2547 N_A_4239_793#_c_3241_n N_S[7]_c_3483_n 9.67113e-19 $X=23.945 $Y=4.74
+ $X2=0 $Y2=0
cc_2548 N_A_4239_793#_c_3242_n N_S[7]_c_3483_n 0.00603996f $X=23.985 $Y=4.995
+ $X2=0 $Y2=0
cc_2549 N_A_4239_793#_c_3241_n N_S[7]_c_3484_n 0.0111895f $X=23.945 $Y=4.74
+ $X2=0 $Y2=0
cc_2550 N_A_4239_793#_c_3244_n N_S[7]_c_3484_n 0.00429801f $X=23.945 $Y=4.615
+ $X2=0 $Y2=0
cc_2551 N_A_4239_793#_c_3259_n N_S[7]_c_3485_n 0.00336772f $X=23.905 $Y=4.045
+ $X2=0 $Y2=0
cc_2552 N_A_4239_793#_c_3241_n N_S[7]_c_3485_n 0.00207203f $X=23.945 $Y=4.74
+ $X2=0 $Y2=0
cc_2553 N_A_4239_793#_c_3260_n N_S[7]_c_3485_n 5.48523e-19 $X=23.985 $Y=3.835
+ $X2=0 $Y2=0
cc_2554 N_A_4239_793#_c_3243_n N_S[7]_c_3485_n 0.00416423f $X=23.905 $Y=4.21
+ $X2=0 $Y2=0
cc_2555 N_A_4239_793#_c_3244_n N_S[7]_c_3485_n 0.00289358f $X=23.945 $Y=4.615
+ $X2=0 $Y2=0
cc_2556 N_A_4239_793#_c_3258_n N_S[7]_c_3495_n 0.0097833f $X=23.985 $Y=3.14
+ $X2=0 $Y2=0
cc_2557 N_A_4239_793#_c_3259_n N_S[7]_c_3495_n 0.00117303f $X=23.905 $Y=4.045
+ $X2=0 $Y2=0
cc_2558 N_A_4239_793#_c_3260_n N_S[7]_c_3495_n 0.00304348f $X=23.985 $Y=3.835
+ $X2=0 $Y2=0
cc_2559 N_A_4239_793#_c_3241_n N_S[7]_c_3489_n 0.00426435f $X=23.945 $Y=4.74
+ $X2=0 $Y2=0
cc_2560 N_A_4239_793#_c_3244_n N_S[7]_c_3489_n 0.00268644f $X=23.945 $Y=4.615
+ $X2=0 $Y2=0
cc_2561 N_A_4239_793#_c_3243_n S[7] 0.0228692f $X=23.905 $Y=4.21 $X2=0 $Y2=0
cc_2562 N_A_4239_793#_c_3244_n S[7] 0.00541767f $X=23.945 $Y=4.615 $X2=0 $Y2=0
cc_2563 N_A_4239_793#_c_3246_n N_VPWR_c_3620_n 0.00324472f $X=21.295 $Y=3.965
+ $X2=0 $Y2=0
cc_2564 N_A_4239_793#_c_3253_n N_VPWR_c_3622_n 0.00377407f $X=22.705 $Y=3.965
+ $X2=0 $Y2=0
cc_2565 N_A_4239_793#_c_3239_n N_VPWR_c_3622_n 0.0208071f $X=23.82 $Y=4.21 $X2=0
+ $Y2=0
cc_2566 N_A_4239_793#_c_3240_n N_VPWR_c_3622_n 6.4101e-19 $X=23.275 $Y=4.21
+ $X2=0 $Y2=0
cc_2567 N_A_4239_793#_c_3258_n N_VPWR_c_3622_n 0.0302744f $X=23.985 $Y=3.14
+ $X2=0 $Y2=0
cc_2568 N_A_4239_793#_c_3258_n N_VPWR_c_3624_n 0.03379f $X=23.985 $Y=3.14 $X2=0
+ $Y2=0
cc_2569 N_A_4239_793#_c_3258_n N_VPWR_c_3649_n 0.0233824f $X=23.985 $Y=3.14
+ $X2=0 $Y2=0
cc_2570 N_A_4239_793#_c_3246_n N_VPWR_c_3661_n 0.00473731f $X=21.295 $Y=3.965
+ $X2=0 $Y2=0
cc_2571 N_A_4239_793#_c_3249_n N_VPWR_c_3661_n 0.00362156f $X=21.765 $Y=3.965
+ $X2=0 $Y2=0
cc_2572 N_A_4239_793#_c_3251_n N_VPWR_c_3661_n 0.00362156f $X=22.235 $Y=3.965
+ $X2=0 $Y2=0
cc_2573 N_A_4239_793#_c_3253_n N_VPWR_c_3661_n 0.00473731f $X=22.705 $Y=3.965
+ $X2=0 $Y2=0
cc_2574 N_A_4239_793#_c_3258_n N_VPWR_c_3661_n 0.0124581f $X=23.985 $Y=3.14
+ $X2=0 $Y2=0
cc_2575 N_A_4239_793#_c_3250_n N_Z_c_4605_n 0.00762343f $X=22.145 $Y=4.04 $X2=0
+ $Y2=0
cc_2576 N_A_4239_793#_c_3254_n N_Z_c_4605_n 0.00704092f $X=21.765 $Y=4.04 $X2=0
+ $Y2=0
cc_2577 N_A_4239_793#_c_3248_n N_Z_c_4630_n 0.00248496f $X=21.385 $Y=4.04 $X2=0
+ $Y2=0
cc_2578 N_A_4239_793#_c_3247_n N_Z_c_4633_n 0.00678861f $X=21.675 $Y=4.04 $X2=0
+ $Y2=0
cc_2579 N_A_4239_793#_c_3248_n N_Z_c_4633_n 0.00239476f $X=21.385 $Y=4.04 $X2=0
+ $Y2=0
cc_2580 N_A_4239_793#_c_3254_n N_Z_c_4633_n 2.98555e-19 $X=21.765 $Y=4.04 $X2=0
+ $Y2=0
cc_2581 N_A_4239_793#_c_3250_n N_Z_c_4635_n 0.00145542f $X=22.145 $Y=4.04 $X2=0
+ $Y2=0
cc_2582 N_A_4239_793#_c_3252_n N_Z_c_4635_n 0.00597584f $X=22.615 $Y=4.04 $X2=0
+ $Y2=0
cc_2583 N_A_4239_793#_c_3255_n N_Z_c_4635_n 0.00909323f $X=22.235 $Y=4.04 $X2=0
+ $Y2=0
cc_2584 N_A_4239_793#_c_3239_n N_Z_c_4635_n 0.0266078f $X=23.82 $Y=4.21 $X2=0
+ $Y2=0
cc_2585 N_A_4239_793#_c_3245_n N_Z_c_4635_n 0.00747617f $X=23.025 $Y=4.21 $X2=0
+ $Y2=0
cc_2586 N_A_4239_793#_c_3246_n N_Z_c_4649_n 0.00834829f $X=21.295 $Y=3.965 $X2=0
+ $Y2=0
cc_2587 N_A_4239_793#_c_3249_n Z 0.00372458f $X=21.765 $Y=3.965 $X2=0 $Y2=0
cc_2588 N_A_4239_793#_c_3251_n Z 0.00372248f $X=22.235 $Y=3.965 $X2=0 $Y2=0
cc_2589 N_A_4239_793#_c_3246_n N_Z_c_4656_n 0.0199111f $X=21.295 $Y=3.965 $X2=0
+ $Y2=0
cc_2590 N_A_4239_793#_c_3247_n N_Z_c_4656_n 0.00560592f $X=21.675 $Y=4.04 $X2=0
+ $Y2=0
cc_2591 N_A_4239_793#_c_3248_n N_Z_c_4656_n 0.00474497f $X=21.385 $Y=4.04 $X2=0
+ $Y2=0
cc_2592 N_A_4239_793#_c_3249_n N_Z_c_4656_n 0.0181262f $X=21.765 $Y=3.965 $X2=0
+ $Y2=0
cc_2593 N_A_4239_793#_c_3251_n N_Z_c_4656_n 9.74366e-19 $X=22.235 $Y=3.965 $X2=0
+ $Y2=0
cc_2594 N_A_4239_793#_c_3254_n N_Z_c_4656_n 0.00415268f $X=21.765 $Y=4.04 $X2=0
+ $Y2=0
cc_2595 N_A_4239_793#_c_3249_n N_Z_c_4657_n 9.74366e-19 $X=21.765 $Y=3.965 $X2=0
+ $Y2=0
cc_2596 N_A_4239_793#_c_3251_n N_Z_c_4657_n 0.0181262f $X=22.235 $Y=3.965 $X2=0
+ $Y2=0
cc_2597 N_A_4239_793#_c_3252_n N_Z_c_4657_n 0.00560592f $X=22.615 $Y=4.04 $X2=0
+ $Y2=0
cc_2598 N_A_4239_793#_c_3253_n N_Z_c_4657_n 0.0226667f $X=22.705 $Y=3.965 $X2=0
+ $Y2=0
cc_2599 N_A_4239_793#_c_3255_n N_Z_c_4657_n 0.00181273f $X=22.235 $Y=4.04 $X2=0
+ $Y2=0
cc_2600 N_A_4239_793#_c_3239_n N_Z_c_4657_n 0.00240108f $X=23.82 $Y=4.21 $X2=0
+ $Y2=0
cc_2601 N_A_4239_793#_c_3245_n N_Z_c_4657_n 0.00425035f $X=23.025 $Y=4.21 $X2=0
+ $Y2=0
cc_2602 N_A_4239_793#_c_3246_n N_A_3797_591#_c_6142_n 0.00151141f $X=21.295
+ $Y=3.965 $X2=0 $Y2=0
cc_2603 N_A_4239_793#_c_3246_n N_A_3797_591#_c_6171_n 0.00307958f $X=21.295
+ $Y=3.965 $X2=0 $Y2=0
cc_2604 N_A_4239_793#_c_3249_n N_A_3797_591#_c_6171_n 0.00307958f $X=21.765
+ $Y=3.965 $X2=0 $Y2=0
cc_2605 N_A_4239_793#_c_3251_n N_A_3797_591#_c_6173_n 0.00307958f $X=22.235
+ $Y=3.965 $X2=0 $Y2=0
cc_2606 N_A_4239_793#_c_3253_n N_A_3797_591#_c_6173_n 0.00799829f $X=22.705
+ $Y=3.965 $X2=0 $Y2=0
cc_2607 N_A_4239_793#_c_3246_n N_A_3797_591#_c_6144_n 0.00554566f $X=21.295
+ $Y=3.965 $X2=0 $Y2=0
cc_2608 N_A_4239_793#_c_3249_n N_A_3797_591#_c_6145_n 0.00210632f $X=21.765
+ $Y=3.965 $X2=0 $Y2=0
cc_2609 N_A_4239_793#_c_3250_n N_A_3797_591#_c_6145_n 0.00251792f $X=22.145
+ $Y=4.04 $X2=0 $Y2=0
cc_2610 N_A_4239_793#_c_3251_n N_A_3797_591#_c_6145_n 0.00210632f $X=22.235
+ $Y=3.965 $X2=0 $Y2=0
cc_2611 N_A_4239_793#_c_3253_n N_A_3797_591#_c_6146_n 0.00483827f $X=22.705
+ $Y=3.965 $X2=0 $Y2=0
cc_2612 N_A_4239_793#_c_3239_n N_A_3797_591#_c_6146_n 0.0229374f $X=23.82
+ $Y=4.21 $X2=0 $Y2=0
cc_2613 N_A_4239_793#_c_3240_n N_A_3797_591#_c_6146_n 5.74251e-19 $X=23.275
+ $Y=4.21 $X2=0 $Y2=0
cc_2614 N_A_4239_793#_c_3245_n N_A_3797_591#_c_6146_n 0.00561627f $X=23.025
+ $Y=4.21 $X2=0 $Y2=0
cc_2615 N_A_4239_793#_c_3239_n N_VGND_c_6303_n 0.0123065f $X=23.82 $Y=4.21 $X2=0
+ $Y2=0
cc_2616 N_A_4239_793#_c_3240_n N_VGND_c_6303_n 2.04129e-19 $X=23.275 $Y=4.21
+ $X2=0 $Y2=0
cc_2617 N_A_4239_793#_c_3242_n N_VGND_c_6353_n 0.0129994f $X=23.985 $Y=4.995
+ $X2=0 $Y2=0
cc_2618 N_A_4239_793#_M1114_d N_VGND_c_6371_n 0.00394793f $X=23.85 $Y=4.785
+ $X2=0 $Y2=0
cc_2619 N_A_4239_793#_c_3242_n N_VGND_c_6371_n 0.00927134f $X=23.985 $Y=4.995
+ $X2=0 $Y2=0
cc_2620 N_A_4239_793#_c_3254_n N_A_3799_911#_c_7527_n 7.0477e-19 $X=21.765
+ $Y=4.04 $X2=0 $Y2=0
cc_2621 N_A_4239_793#_c_3239_n N_A_3799_911#_c_7508_n 0.0028695f $X=23.82
+ $Y=4.21 $X2=0 $Y2=0
cc_2622 N_A_4239_793#_c_3245_n N_A_3799_911#_c_7508_n 0.00589316f $X=23.025
+ $Y=4.21 $X2=0 $Y2=0
cc_2623 N_S[6]_c_3383_n N_S[7]_c_3493_n 0.0130744f $X=23.75 $Y=1.55 $X2=0 $Y2=0
cc_2624 N_S[6]_c_3376_n N_S[7]_c_3495_n 0.0130744f $X=24.22 $Y=1.55 $X2=0 $Y2=0
cc_2625 N_S[6]_c_3383_n N_VPWR_c_3621_n 0.00929376f $X=23.75 $Y=1.55 $X2=0 $Y2=0
cc_2626 N_S[6]_c_3376_n N_VPWR_c_3623_n 0.0161848f $X=24.22 $Y=1.55 $X2=0 $Y2=0
cc_2627 S[6] N_VPWR_c_3623_n 0.017333f $X=24.525 $Y=1.105 $X2=0 $Y2=0
cc_2628 N_S[6]_c_3383_n N_VPWR_c_3649_n 0.0035837f $X=23.75 $Y=1.55 $X2=0 $Y2=0
cc_2629 N_S[6]_c_3376_n N_VPWR_c_3649_n 0.0035837f $X=24.22 $Y=1.55 $X2=0 $Y2=0
cc_2630 N_S[6]_c_3383_n N_VPWR_c_3661_n 0.0118174f $X=23.75 $Y=1.55 $X2=0 $Y2=0
cc_2631 N_S[6]_c_3376_n N_VPWR_c_3661_n 0.0114704f $X=24.22 $Y=1.55 $X2=0 $Y2=0
cc_2632 N_S[6]_c_3360_n N_Z_c_4603_n 0.002324f $X=21.22 $Y=0.255 $X2=0 $Y2=0
cc_2633 N_S[6]_c_3363_n N_Z_c_4603_n 0.00283489f $X=21.64 $Y=0.255 $X2=0 $Y2=0
cc_2634 N_S[6]_c_3363_n N_Z_c_4604_n 3.10191e-19 $X=21.64 $Y=0.255 $X2=0 $Y2=0
cc_2635 N_S[6]_c_3365_n N_Z_c_4604_n 0.00190704f $X=22.06 $Y=0.255 $X2=0 $Y2=0
cc_2636 N_S[6]_c_3363_n N_Z_c_4606_n 6.35774e-19 $X=21.64 $Y=0.255 $X2=0 $Y2=0
cc_2637 N_S[6]_c_3365_n N_Z_c_4606_n 0.0077801f $X=22.06 $Y=0.255 $X2=0 $Y2=0
cc_2638 N_S[6]_c_3367_n N_Z_c_4606_n 0.0134253f $X=22.48 $Y=0.255 $X2=0 $Y2=0
cc_2639 N_S[6]_c_3360_n N_Z_c_4629_n 0.00443615f $X=21.22 $Y=0.255 $X2=0 $Y2=0
cc_2640 N_S[6]_c_3363_n N_Z_c_4629_n 0.00462308f $X=21.64 $Y=0.255 $X2=0 $Y2=0
cc_2641 N_S[6]_c_3365_n N_Z_c_4629_n 6.35664e-19 $X=22.06 $Y=0.255 $X2=0 $Y2=0
cc_2642 N_S[6]_c_3363_n N_Z_c_4632_n 0.00180363f $X=21.64 $Y=0.255 $X2=0 $Y2=0
cc_2643 N_S[6]_c_3367_n N_Z_c_4634_n 0.00216436f $X=22.48 $Y=0.255 $X2=0 $Y2=0
cc_2644 N_S[6]_c_3360_n N_A_3797_297#_c_6020_n 0.00168571f $X=21.22 $Y=0.255
+ $X2=0 $Y2=0
cc_2645 N_S[6]_c_3383_n N_A_3797_297#_c_6024_n 0.00249814f $X=23.75 $Y=1.55
+ $X2=0 $Y2=0
cc_2646 N_S[6]_c_3360_n N_VGND_c_6300_n 5.5039e-19 $X=21.22 $Y=0.255 $X2=0 $Y2=0
cc_2647 N_S[6]_c_3362_n N_VGND_c_6300_n 0.0028166f $X=21.295 $Y=0.18 $X2=0 $Y2=0
cc_2648 N_S[6]_c_3368_n N_VGND_c_6302_n 0.00862298f $X=23.165 $Y=0.18 $X2=0
+ $Y2=0
cc_2649 N_S[6]_c_3370_n N_VGND_c_6302_n 0.00525833f $X=23.65 $Y=0.81 $X2=0 $Y2=0
cc_2650 N_S[6]_c_3373_n N_VGND_c_6302_n 0.00173127f $X=23.775 $Y=0.735 $X2=0
+ $Y2=0
cc_2651 N_S[6]_c_3375_n N_VGND_c_6305_n 0.00374526f $X=24.195 $Y=0.735 $X2=0
+ $Y2=0
cc_2652 N_S[6]_c_3376_n N_VGND_c_6305_n 0.00578076f $X=24.22 $Y=1.55 $X2=0 $Y2=0
cc_2653 S[6] N_VGND_c_6305_n 0.0116413f $X=24.525 $Y=1.105 $X2=0 $Y2=0
cc_2654 N_S[6]_c_3362_n N_VGND_c_6336_n 0.0559651f $X=21.295 $Y=0.18 $X2=0 $Y2=0
cc_2655 N_S[6]_c_3373_n N_VGND_c_6352_n 0.00542362f $X=23.775 $Y=0.735 $X2=0
+ $Y2=0
cc_2656 N_S[6]_c_3374_n N_VGND_c_6352_n 2.16067e-19 $X=24.12 $Y=0.81 $X2=0 $Y2=0
cc_2657 N_S[6]_c_3375_n N_VGND_c_6352_n 0.00585385f $X=24.195 $Y=0.735 $X2=0
+ $Y2=0
cc_2658 N_S[6]_c_3361_n N_VGND_c_6370_n 0.00642387f $X=21.565 $Y=0.18 $X2=0
+ $Y2=0
cc_2659 N_S[6]_c_3362_n N_VGND_c_6370_n 0.00591981f $X=21.295 $Y=0.18 $X2=0
+ $Y2=0
cc_2660 N_S[6]_c_3364_n N_VGND_c_6370_n 0.0064237f $X=21.985 $Y=0.18 $X2=0 $Y2=0
cc_2661 N_S[6]_c_3366_n N_VGND_c_6370_n 0.00642387f $X=22.405 $Y=0.18 $X2=0
+ $Y2=0
cc_2662 N_S[6]_c_3368_n N_VGND_c_6370_n 0.0345801f $X=23.165 $Y=0.18 $X2=0 $Y2=0
cc_2663 N_S[6]_c_3373_n N_VGND_c_6370_n 0.00990284f $X=23.775 $Y=0.735 $X2=0
+ $Y2=0
cc_2664 N_S[6]_c_3375_n N_VGND_c_6370_n 0.0117149f $X=24.195 $Y=0.735 $X2=0
+ $Y2=0
cc_2665 N_S[6]_c_3377_n N_VGND_c_6370_n 0.00366655f $X=21.64 $Y=0.18 $X2=0 $Y2=0
cc_2666 N_S[6]_c_3378_n N_VGND_c_6370_n 0.00366655f $X=22.06 $Y=0.18 $X2=0 $Y2=0
cc_2667 N_S[6]_c_3379_n N_VGND_c_6370_n 0.00366655f $X=22.48 $Y=0.18 $X2=0 $Y2=0
cc_2668 N_S[6]_c_3360_n N_A_3799_47#_c_7421_n 0.00206084f $X=21.22 $Y=0.255
+ $X2=0 $Y2=0
cc_2669 N_S[6]_c_3360_n N_A_3799_47#_c_7423_n 0.0139014f $X=21.22 $Y=0.255 $X2=0
+ $Y2=0
cc_2670 N_S[6]_c_3361_n N_A_3799_47#_c_7423_n 0.00211351f $X=21.565 $Y=0.18
+ $X2=0 $Y2=0
cc_2671 N_S[6]_c_3363_n N_A_3799_47#_c_7423_n 0.0106826f $X=21.64 $Y=0.255 $X2=0
+ $Y2=0
cc_2672 N_S[6]_c_3365_n N_A_3799_47#_c_7425_n 0.0106844f $X=22.06 $Y=0.255 $X2=0
+ $Y2=0
cc_2673 N_S[6]_c_3366_n N_A_3799_47#_c_7425_n 0.00211351f $X=22.405 $Y=0.18
+ $X2=0 $Y2=0
cc_2674 N_S[6]_c_3367_n N_A_3799_47#_c_7425_n 0.0112916f $X=22.48 $Y=0.255 $X2=0
+ $Y2=0
cc_2675 N_S[6]_c_3368_n N_A_3799_47#_c_7425_n 0.00685838f $X=23.165 $Y=0.18
+ $X2=0 $Y2=0
cc_2676 N_S[6]_c_3369_n N_A_3799_47#_c_7425_n 0.00189496f $X=23.24 $Y=0.735
+ $X2=0 $Y2=0
cc_2677 N_S[6]_c_3369_n N_A_3799_47#_c_7426_n 0.00529837f $X=23.24 $Y=0.735
+ $X2=0 $Y2=0
cc_2678 N_S[6]_c_3364_n N_A_3799_47#_c_7461_n 0.0034777f $X=21.985 $Y=0.18 $X2=0
+ $Y2=0
cc_2679 N_S[7]_c_3493_n N_VPWR_c_3622_n 0.00929376f $X=23.75 $Y=3.89 $X2=0 $Y2=0
cc_2680 N_S[7]_c_3485_n N_VPWR_c_3624_n 0.00652399f $X=24.195 $Y=4.705 $X2=0
+ $Y2=0
cc_2681 N_S[7]_c_3495_n N_VPWR_c_3624_n 0.00966078f $X=24.22 $Y=3.89 $X2=0 $Y2=0
cc_2682 S[7] N_VPWR_c_3624_n 0.017333f $X=24.525 $Y=4.165 $X2=0 $Y2=0
cc_2683 N_S[7]_c_3493_n N_VPWR_c_3649_n 0.0035837f $X=23.75 $Y=3.89 $X2=0 $Y2=0
cc_2684 N_S[7]_c_3495_n N_VPWR_c_3649_n 0.0035837f $X=24.22 $Y=3.89 $X2=0 $Y2=0
cc_2685 N_S[7]_c_3493_n N_VPWR_c_3661_n 0.0118174f $X=23.75 $Y=3.89 $X2=0 $Y2=0
cc_2686 N_S[7]_c_3495_n N_VPWR_c_3661_n 0.0114704f $X=24.22 $Y=3.89 $X2=0 $Y2=0
cc_2687 N_S[7]_c_3473_n N_Z_c_4605_n 3.10191e-19 $X=21.64 $Y=5.185 $X2=0 $Y2=0
cc_2688 N_S[7]_c_3475_n N_Z_c_4605_n 0.00190704f $X=22.06 $Y=5.185 $X2=0 $Y2=0
cc_2689 N_S[7]_c_3473_n N_Z_c_4607_n 6.35774e-19 $X=21.64 $Y=5.185 $X2=0 $Y2=0
cc_2690 N_S[7]_c_3475_n N_Z_c_4607_n 0.0077801f $X=22.06 $Y=5.185 $X2=0 $Y2=0
cc_2691 N_S[7]_c_3477_n N_Z_c_4607_n 0.0134253f $X=22.48 $Y=5.185 $X2=0 $Y2=0
cc_2692 N_S[7]_c_3470_n N_Z_c_4630_n 0.00443615f $X=21.22 $Y=5.185 $X2=0 $Y2=0
cc_2693 N_S[7]_c_3473_n N_Z_c_4630_n 0.00462308f $X=21.64 $Y=5.185 $X2=0 $Y2=0
cc_2694 N_S[7]_c_3470_n N_Z_c_4631_n 0.002324f $X=21.22 $Y=5.185 $X2=0 $Y2=0
cc_2695 N_S[7]_c_3473_n N_Z_c_4631_n 0.00283489f $X=21.64 $Y=5.185 $X2=0 $Y2=0
cc_2696 N_S[7]_c_3475_n N_Z_c_4631_n 6.35664e-19 $X=22.06 $Y=5.185 $X2=0 $Y2=0
cc_2697 N_S[7]_c_3473_n N_Z_c_4633_n 0.00180363f $X=21.64 $Y=5.185 $X2=0 $Y2=0
cc_2698 N_S[7]_c_3477_n N_Z_c_4635_n 0.00216436f $X=22.48 $Y=5.185 $X2=0 $Y2=0
cc_2699 N_S[7]_c_3470_n N_A_3797_591#_c_6142_n 0.00168571f $X=21.22 $Y=5.185
+ $X2=0 $Y2=0
cc_2700 N_S[7]_c_3493_n N_A_3797_591#_c_6146_n 0.00249814f $X=23.75 $Y=3.89
+ $X2=0 $Y2=0
cc_2701 N_S[7]_c_3470_n N_VGND_c_6301_n 5.5039e-19 $X=21.22 $Y=5.185 $X2=0 $Y2=0
cc_2702 N_S[7]_c_3472_n N_VGND_c_6301_n 0.0028166f $X=21.295 $Y=5.26 $X2=0 $Y2=0
cc_2703 N_S[7]_c_3479_n N_VGND_c_6303_n 0.00862298f $X=23.24 $Y=5.185 $X2=0
+ $Y2=0
cc_2704 N_S[7]_c_3480_n N_VGND_c_6303_n 0.00525833f $X=23.65 $Y=4.63 $X2=0 $Y2=0
cc_2705 N_S[7]_c_3483_n N_VGND_c_6303_n 0.00173127f $X=23.775 $Y=4.705 $X2=0
+ $Y2=0
cc_2706 N_S[7]_c_3485_n N_VGND_c_6307_n 0.00952602f $X=24.195 $Y=4.705 $X2=0
+ $Y2=0
cc_2707 S[7] N_VGND_c_6307_n 0.0116413f $X=24.525 $Y=4.165 $X2=0 $Y2=0
cc_2708 N_S[7]_c_3472_n N_VGND_c_6338_n 0.0559651f $X=21.295 $Y=5.26 $X2=0 $Y2=0
cc_2709 N_S[7]_c_3483_n N_VGND_c_6353_n 0.00542362f $X=23.775 $Y=4.705 $X2=0
+ $Y2=0
cc_2710 N_S[7]_c_3484_n N_VGND_c_6353_n 2.16067e-19 $X=24.12 $Y=4.63 $X2=0 $Y2=0
cc_2711 N_S[7]_c_3485_n N_VGND_c_6353_n 0.00585385f $X=24.195 $Y=4.705 $X2=0
+ $Y2=0
cc_2712 N_S[7]_c_3471_n N_VGND_c_6371_n 0.00642387f $X=21.565 $Y=5.26 $X2=0
+ $Y2=0
cc_2713 N_S[7]_c_3472_n N_VGND_c_6371_n 0.00591981f $X=21.295 $Y=5.26 $X2=0
+ $Y2=0
cc_2714 N_S[7]_c_3474_n N_VGND_c_6371_n 0.0064237f $X=21.985 $Y=5.26 $X2=0 $Y2=0
cc_2715 N_S[7]_c_3476_n N_VGND_c_6371_n 0.00642387f $X=22.405 $Y=5.26 $X2=0
+ $Y2=0
cc_2716 N_S[7]_c_3478_n N_VGND_c_6371_n 0.0345801f $X=23.165 $Y=5.26 $X2=0 $Y2=0
cc_2717 N_S[7]_c_3483_n N_VGND_c_6371_n 0.00990284f $X=23.775 $Y=4.705 $X2=0
+ $Y2=0
cc_2718 N_S[7]_c_3485_n N_VGND_c_6371_n 0.0117149f $X=24.195 $Y=4.705 $X2=0
+ $Y2=0
cc_2719 N_S[7]_c_3486_n N_VGND_c_6371_n 0.00366655f $X=21.64 $Y=5.26 $X2=0 $Y2=0
cc_2720 N_S[7]_c_3487_n N_VGND_c_6371_n 0.00366655f $X=22.06 $Y=5.26 $X2=0 $Y2=0
cc_2721 N_S[7]_c_3488_n N_VGND_c_6371_n 0.00366655f $X=22.48 $Y=5.26 $X2=0 $Y2=0
cc_2722 N_S[7]_c_3470_n N_A_3799_911#_c_7503_n 0.00206084f $X=21.22 $Y=5.185
+ $X2=0 $Y2=0
cc_2723 N_S[7]_c_3470_n N_A_3799_911#_c_7505_n 0.0139014f $X=21.22 $Y=5.185
+ $X2=0 $Y2=0
cc_2724 N_S[7]_c_3471_n N_A_3799_911#_c_7505_n 0.00211351f $X=21.565 $Y=5.26
+ $X2=0 $Y2=0
cc_2725 N_S[7]_c_3473_n N_A_3799_911#_c_7505_n 0.0106826f $X=21.64 $Y=5.185
+ $X2=0 $Y2=0
cc_2726 N_S[7]_c_3475_n N_A_3799_911#_c_7507_n 0.0106844f $X=22.06 $Y=5.185
+ $X2=0 $Y2=0
cc_2727 N_S[7]_c_3476_n N_A_3799_911#_c_7507_n 0.00211351f $X=22.405 $Y=5.26
+ $X2=0 $Y2=0
cc_2728 N_S[7]_c_3477_n N_A_3799_911#_c_7507_n 0.0112916f $X=22.48 $Y=5.185
+ $X2=0 $Y2=0
cc_2729 N_S[7]_c_3478_n N_A_3799_911#_c_7507_n 0.00685838f $X=23.165 $Y=5.26
+ $X2=0 $Y2=0
cc_2730 N_S[7]_c_3479_n N_A_3799_911#_c_7507_n 0.00189496f $X=23.24 $Y=5.185
+ $X2=0 $Y2=0
cc_2731 N_S[7]_c_3481_n N_A_3799_911#_c_7508_n 0.00529837f $X=23.315 $Y=4.63
+ $X2=0 $Y2=0
cc_2732 N_S[7]_c_3474_n N_A_3799_911#_c_7540_n 0.0034777f $X=21.985 $Y=5.26
+ $X2=0 $Y2=0
cc_2733 N_VPWR_c_3661_n N_A_355_311#_M1012_d 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2734 N_VPWR_c_3661_n N_A_355_311#_M1086_d 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2735 N_VPWR_M1012_s N_A_355_311#_c_4334_n 0.00715085f $X=4.175 $Y=1.485 $X2=0
+ $Y2=0
cc_2736 N_VPWR_c_3590_n N_A_355_311#_c_4334_n 0.0152464f $X=4.3 $Y=2 $X2=0 $Y2=0
cc_2737 N_VPWR_M1049_s N_A_355_311#_c_4356_n 0.00331615f $X=5.095 $Y=1.485 $X2=0
+ $Y2=0
cc_2738 N_VPWR_c_3592_n N_A_355_311#_c_4356_n 0.0130979f $X=5.24 $Y=2 $X2=0
+ $Y2=0
cc_2739 N_VPWR_c_3661_n N_A_355_311#_c_4343_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2740 N_VPWR_c_3588_n N_A_355_311#_c_4385_n 0.00167067f $X=1.325 $Y=1.77 $X2=0
+ $Y2=0
cc_2741 N_VPWR_c_3661_n N_A_355_311#_c_4385_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2742 N_VPWR_c_3661_n N_A_355_311#_c_4345_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2743 N_VPWR_c_3661_n N_A_355_311#_c_4388_n 0.0296491f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2744 N_VPWR_c_3590_n N_A_355_311#_c_4336_n 0.0156478f $X=4.3 $Y=2 $X2=0 $Y2=0
cc_2745 N_VPWR_c_3628_n N_A_355_311#_c_4336_n 0.00115812f $X=4.165 $Y=2.72 $X2=0
+ $Y2=0
cc_2746 N_VPWR_c_3641_n N_A_355_311#_c_4336_n 8.30334e-19 $X=5.105 $Y=2.72 $X2=0
+ $Y2=0
cc_2747 N_VPWR_c_3661_n N_A_355_311#_c_4336_n 0.0605692f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2748 N_VPWR_c_3590_n N_A_355_311#_c_4393_n 6.69936e-19 $X=4.3 $Y=2 $X2=0
+ $Y2=0
cc_2749 N_VPWR_c_3661_n N_A_355_311#_c_4393_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2750 N_VPWR_c_3592_n N_A_355_311#_c_4369_n 0.0153177f $X=5.24 $Y=2 $X2=0
+ $Y2=0
cc_2751 N_VPWR_c_3641_n N_A_355_311#_c_4369_n 8.30334e-19 $X=5.105 $Y=2.72 $X2=0
+ $Y2=0
cc_2752 N_VPWR_c_3642_n N_A_355_311#_c_4369_n 8.30334e-19 $X=6.045 $Y=2.72 $X2=0
+ $Y2=0
cc_2753 N_VPWR_c_3661_n N_A_355_311#_c_4369_n 0.0558368f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2754 N_VPWR_c_3590_n N_A_355_311#_c_4399_n 6.68271e-19 $X=4.3 $Y=2 $X2=0
+ $Y2=0
cc_2755 N_VPWR_c_3592_n N_A_355_311#_c_4399_n 6.68271e-19 $X=5.24 $Y=2 $X2=0
+ $Y2=0
cc_2756 N_VPWR_c_3661_n N_A_355_311#_c_4399_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2757 N_VPWR_c_3590_n N_A_355_311#_c_4371_n 0.0268237f $X=4.3 $Y=2 $X2=0 $Y2=0
cc_2758 N_VPWR_c_3592_n N_A_355_311#_c_4371_n 0.0268237f $X=5.24 $Y=2 $X2=0
+ $Y2=0
cc_2759 N_VPWR_c_3641_n N_A_355_311#_c_4371_n 0.0189467f $X=5.105 $Y=2.72 $X2=0
+ $Y2=0
cc_2760 N_VPWR_c_3661_n N_A_355_311#_c_4371_n 0.00300637f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2761 N_VPWR_c_3592_n N_A_355_311#_c_4406_n 6.68271e-19 $X=5.24 $Y=2 $X2=0
+ $Y2=0
cc_2762 N_VPWR_c_3594_n N_A_355_311#_c_4406_n 0.00170069f $X=6.21 $Y=1.66 $X2=0
+ $Y2=0
cc_2763 N_VPWR_c_3661_n N_A_355_311#_c_4406_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2764 N_VPWR_c_3592_n N_A_355_311#_c_4374_n 0.0268237f $X=5.24 $Y=2 $X2=0
+ $Y2=0
cc_2765 N_VPWR_c_3594_n N_A_355_311#_c_4374_n 0.031816f $X=6.21 $Y=1.66 $X2=0
+ $Y2=0
cc_2766 N_VPWR_c_3642_n N_A_355_311#_c_4374_n 0.0189467f $X=6.045 $Y=2.72 $X2=0
+ $Y2=0
cc_2767 N_VPWR_c_3661_n N_A_355_311#_c_4374_n 0.00313104f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2768 N_VPWR_c_3588_n N_A_355_311#_c_4337_n 0.0523777f $X=1.325 $Y=1.77 $X2=0
+ $Y2=0
cc_2769 N_VPWR_c_3625_n N_A_355_311#_c_4337_n 0.0213652f $X=1.49 $Y=2.72 $X2=0
+ $Y2=0
cc_2770 N_VPWR_c_3661_n N_A_355_311#_c_4337_n 0.00302891f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2771 N_VPWR_c_3661_n N_A_355_311#_c_4338_n 0.00468575f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2772 N_VPWR_c_3590_n N_A_355_311#_c_4339_n 0.0390576f $X=4.3 $Y=2 $X2=0 $Y2=0
cc_2773 N_VPWR_c_3628_n N_A_355_311#_c_4339_n 0.0213652f $X=4.165 $Y=2.72 $X2=0
+ $Y2=0
cc_2774 N_VPWR_c_3661_n N_A_355_311#_c_4339_n 0.0027766f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2775 N_VPWR_c_3661_n N_A_355_613#_M1017_d 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2776 N_VPWR_c_3661_n N_A_355_613#_M1093_d 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2777 N_VPWR_M1017_s N_A_355_613#_c_4461_n 0.00715085f $X=4.175 $Y=2.955 $X2=0
+ $Y2=0
cc_2778 N_VPWR_c_3591_n N_A_355_613#_c_4461_n 0.0152464f $X=4.3 $Y=3.1 $X2=0
+ $Y2=0
cc_2779 N_VPWR_M1055_s N_A_355_613#_c_4483_n 0.00331615f $X=5.095 $Y=2.955 $X2=0
+ $Y2=0
cc_2780 N_VPWR_c_3593_n N_A_355_613#_c_4483_n 0.0130979f $X=5.24 $Y=3.1 $X2=0
+ $Y2=0
cc_2781 N_VPWR_c_3661_n N_A_355_613#_c_4470_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2782 N_VPWR_c_3589_n N_A_355_613#_c_4512_n 0.00167067f $X=1.325 $Y=3.14 $X2=0
+ $Y2=0
cc_2783 N_VPWR_c_3661_n N_A_355_613#_c_4512_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2784 N_VPWR_c_3661_n N_A_355_613#_c_4472_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2785 N_VPWR_c_3661_n N_A_355_613#_c_4515_n 0.0296491f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2786 N_VPWR_c_3591_n N_A_355_613#_c_4463_n 0.0156478f $X=4.3 $Y=3.1 $X2=0
+ $Y2=0
cc_2787 N_VPWR_c_3628_n N_A_355_613#_c_4463_n 0.00115812f $X=4.165 $Y=2.72 $X2=0
+ $Y2=0
cc_2788 N_VPWR_c_3641_n N_A_355_613#_c_4463_n 8.30334e-19 $X=5.105 $Y=2.72 $X2=0
+ $Y2=0
cc_2789 N_VPWR_c_3661_n N_A_355_613#_c_4463_n 0.0605692f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2790 N_VPWR_c_3591_n N_A_355_613#_c_4520_n 6.69936e-19 $X=4.3 $Y=3.1 $X2=0
+ $Y2=0
cc_2791 N_VPWR_c_3661_n N_A_355_613#_c_4520_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2792 N_VPWR_c_3593_n N_A_355_613#_c_4496_n 0.0153177f $X=5.24 $Y=3.1 $X2=0
+ $Y2=0
cc_2793 N_VPWR_c_3641_n N_A_355_613#_c_4496_n 8.30334e-19 $X=5.105 $Y=2.72 $X2=0
+ $Y2=0
cc_2794 N_VPWR_c_3642_n N_A_355_613#_c_4496_n 8.30334e-19 $X=6.045 $Y=2.72 $X2=0
+ $Y2=0
cc_2795 N_VPWR_c_3661_n N_A_355_613#_c_4496_n 0.0558368f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2796 N_VPWR_c_3591_n N_A_355_613#_c_4526_n 6.68271e-19 $X=4.3 $Y=3.1 $X2=0
+ $Y2=0
cc_2797 N_VPWR_c_3593_n N_A_355_613#_c_4526_n 6.68271e-19 $X=5.24 $Y=3.1 $X2=0
+ $Y2=0
cc_2798 N_VPWR_c_3661_n N_A_355_613#_c_4526_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2799 N_VPWR_c_3593_n N_A_355_613#_c_4529_n 6.68271e-19 $X=5.24 $Y=3.1 $X2=0
+ $Y2=0
cc_2800 N_VPWR_c_3595_n N_A_355_613#_c_4529_n 0.00170069f $X=6.21 $Y=3.1 $X2=0
+ $Y2=0
cc_2801 N_VPWR_c_3661_n N_A_355_613#_c_4529_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2802 N_VPWR_c_3589_n N_A_355_613#_c_4464_n 0.0523777f $X=1.325 $Y=3.14 $X2=0
+ $Y2=0
cc_2803 N_VPWR_c_3625_n N_A_355_613#_c_4464_n 0.0213652f $X=1.49 $Y=2.72 $X2=0
+ $Y2=0
cc_2804 N_VPWR_c_3661_n N_A_355_613#_c_4464_n 0.00302891f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2805 N_VPWR_c_3661_n N_A_355_613#_c_4465_n 0.00468575f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2806 N_VPWR_c_3591_n N_A_355_613#_c_4466_n 0.0390576f $X=4.3 $Y=3.1 $X2=0
+ $Y2=0
cc_2807 N_VPWR_c_3628_n N_A_355_613#_c_4466_n 0.0213652f $X=4.165 $Y=2.72 $X2=0
+ $Y2=0
cc_2808 N_VPWR_c_3661_n N_A_355_613#_c_4466_n 0.0027766f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2809 N_VPWR_c_3591_n N_A_355_613#_c_4499_n 0.0268237f $X=4.3 $Y=3.1 $X2=0
+ $Y2=0
cc_2810 N_VPWR_c_3593_n N_A_355_613#_c_4499_n 0.0268237f $X=5.24 $Y=3.1 $X2=0
+ $Y2=0
cc_2811 N_VPWR_c_3641_n N_A_355_613#_c_4499_n 0.0189467f $X=5.105 $Y=2.72 $X2=0
+ $Y2=0
cc_2812 N_VPWR_c_3661_n N_A_355_613#_c_4499_n 0.00300637f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2813 N_VPWR_c_3593_n N_A_355_613#_c_4502_n 0.0268237f $X=5.24 $Y=3.1 $X2=0
+ $Y2=0
cc_2814 N_VPWR_c_3595_n N_A_355_613#_c_4502_n 0.031816f $X=6.21 $Y=3.1 $X2=0
+ $Y2=0
cc_2815 N_VPWR_c_3642_n N_A_355_613#_c_4502_n 0.0189467f $X=6.045 $Y=2.72 $X2=0
+ $Y2=0
cc_2816 N_VPWR_c_3661_n N_A_355_613#_c_4502_n 0.00313104f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2817 N_VPWR_M1012_s N_Z_c_4644_n 0.00213438f $X=4.175 $Y=1.485 $X2=0 $Y2=0
cc_2818 N_VPWR_M1049_s N_Z_c_4644_n 0.00236137f $X=5.095 $Y=1.485 $X2=0 $Y2=0
cc_2819 N_VPWR_M1137_s N_Z_c_4644_n 4.10081e-19 $X=6.035 $Y=1.485 $X2=0 $Y2=0
cc_2820 N_VPWR_M1090_d N_Z_c_4644_n 0.00236137f $X=7.035 $Y=1.485 $X2=0 $Y2=0
cc_2821 N_VPWR_M1158_d N_Z_c_4644_n 0.00213438f $X=7.975 $Y=1.485 $X2=0 $Y2=0
cc_2822 N_VPWR_c_3590_n N_Z_c_4644_n 0.0106064f $X=4.3 $Y=2 $X2=0 $Y2=0
cc_2823 N_VPWR_c_3592_n N_Z_c_4644_n 0.010348f $X=5.24 $Y=2 $X2=0 $Y2=0
cc_2824 N_VPWR_c_3594_n N_Z_c_4644_n 0.0326935f $X=6.21 $Y=1.66 $X2=0 $Y2=0
cc_2825 N_VPWR_c_3596_n N_Z_c_4644_n 0.010348f $X=7.18 $Y=2 $X2=0 $Y2=0
cc_2826 N_VPWR_c_3599_n N_Z_c_4644_n 0.0106064f $X=8.12 $Y=2 $X2=0 $Y2=0
cc_2827 N_VPWR_c_3661_n N_Z_c_4644_n 0.0317429f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2828 N_VPWR_M1017_s N_Z_c_4645_n 0.00213438f $X=4.175 $Y=2.955 $X2=0 $Y2=0
cc_2829 N_VPWR_M1055_s N_Z_c_4645_n 0.00236137f $X=5.095 $Y=2.955 $X2=0 $Y2=0
cc_2830 N_VPWR_M1141_s N_Z_c_4645_n 4.10081e-19 $X=6.035 $Y=2.955 $X2=0 $Y2=0
cc_2831 N_VPWR_M1076_s N_Z_c_4645_n 0.00236137f $X=7.035 $Y=2.955 $X2=0 $Y2=0
cc_2832 N_VPWR_M1120_s N_Z_c_4645_n 0.00213438f $X=7.975 $Y=2.955 $X2=0 $Y2=0
cc_2833 N_VPWR_c_3591_n N_Z_c_4645_n 0.0106064f $X=4.3 $Y=3.1 $X2=0 $Y2=0
cc_2834 N_VPWR_c_3593_n N_Z_c_4645_n 0.010348f $X=5.24 $Y=3.1 $X2=0 $Y2=0
cc_2835 N_VPWR_c_3595_n N_Z_c_4645_n 0.0326935f $X=6.21 $Y=3.1 $X2=0 $Y2=0
cc_2836 N_VPWR_c_3597_n N_Z_c_4645_n 0.010348f $X=7.18 $Y=3.1 $X2=0 $Y2=0
cc_2837 N_VPWR_c_3600_n N_Z_c_4645_n 0.0106064f $X=8.12 $Y=3.1 $X2=0 $Y2=0
cc_2838 N_VPWR_c_3661_n N_Z_c_4645_n 0.0317429f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2839 N_VPWR_M1072_d N_Z_c_4646_n 8.15553e-19 $X=10.97 $Y=1.625 $X2=0 $Y2=0
cc_2840 N_VPWR_M1115_d N_Z_c_4646_n 2.0504e-19 $X=11.89 $Y=1.625 $X2=0 $Y2=0
cc_2841 N_VPWR_M1128_d N_Z_c_4646_n 2.0504e-19 $X=12.68 $Y=1.625 $X2=0 $Y2=0
cc_2842 N_VPWR_M1155_d N_Z_c_4646_n 8.15553e-19 $X=13.6 $Y=1.625 $X2=0 $Y2=0
cc_2843 N_VPWR_c_3601_n N_Z_c_4646_n 0.0196216f $X=11.095 $Y=1.77 $X2=0 $Y2=0
cc_2844 N_VPWR_c_3603_n N_Z_c_4646_n 0.0222682f $X=12.035 $Y=1.77 $X2=0 $Y2=0
cc_2845 N_VPWR_c_3606_n N_Z_c_4646_n 0.0222682f $X=12.805 $Y=1.77 $X2=0 $Y2=0
cc_2846 N_VPWR_c_3608_n N_Z_c_4646_n 0.0196216f $X=13.745 $Y=1.77 $X2=0 $Y2=0
cc_2847 N_VPWR_c_3661_n N_Z_c_4646_n 0.164379f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2848 N_VPWR_M1007_s N_Z_c_4647_n 8.15553e-19 $X=10.97 $Y=2.995 $X2=0 $Y2=0
cc_2849 N_VPWR_M1125_s N_Z_c_4647_n 2.0504e-19 $X=11.89 $Y=2.995 $X2=0 $Y2=0
cc_2850 N_VPWR_M1018_d N_Z_c_4647_n 2.0504e-19 $X=12.68 $Y=2.995 $X2=0 $Y2=0
cc_2851 N_VPWR_M1039_d N_Z_c_4647_n 8.15553e-19 $X=13.6 $Y=2.995 $X2=0 $Y2=0
cc_2852 N_VPWR_c_3602_n N_Z_c_4647_n 0.0196216f $X=11.095 $Y=3.14 $X2=0 $Y2=0
cc_2853 N_VPWR_c_3604_n N_Z_c_4647_n 0.0222682f $X=12.035 $Y=3.14 $X2=0 $Y2=0
cc_2854 N_VPWR_c_3607_n N_Z_c_4647_n 0.0222682f $X=12.805 $Y=3.14 $X2=0 $Y2=0
cc_2855 N_VPWR_c_3609_n N_Z_c_4647_n 0.0196216f $X=13.745 $Y=3.14 $X2=0 $Y2=0
cc_2856 N_VPWR_c_3661_n N_Z_c_4647_n 0.164379f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2857 N_VPWR_M1042_d N_Z_c_4648_n 0.00213438f $X=16.595 $Y=1.485 $X2=0 $Y2=0
cc_2858 N_VPWR_M1062_d N_Z_c_4648_n 0.00236137f $X=17.515 $Y=1.485 $X2=0 $Y2=0
cc_2859 N_VPWR_M1127_d N_Z_c_4648_n 4.10081e-19 $X=18.455 $Y=1.485 $X2=0 $Y2=0
cc_2860 N_VPWR_M1108_s N_Z_c_4648_n 0.00236137f $X=19.455 $Y=1.485 $X2=0 $Y2=0
cc_2861 N_VPWR_M1145_s N_Z_c_4648_n 0.00213438f $X=20.395 $Y=1.485 $X2=0 $Y2=0
cc_2862 N_VPWR_c_3610_n N_Z_c_4648_n 0.0106064f $X=16.72 $Y=2 $X2=0 $Y2=0
cc_2863 N_VPWR_c_3612_n N_Z_c_4648_n 0.010348f $X=17.66 $Y=2 $X2=0 $Y2=0
cc_2864 N_VPWR_c_3614_n N_Z_c_4648_n 0.0326935f $X=18.63 $Y=1.66 $X2=0 $Y2=0
cc_2865 N_VPWR_c_3616_n N_Z_c_4648_n 0.010348f $X=19.6 $Y=2 $X2=0 $Y2=0
cc_2866 N_VPWR_c_3619_n N_Z_c_4648_n 0.0106064f $X=20.54 $Y=2 $X2=0 $Y2=0
cc_2867 N_VPWR_c_3661_n N_Z_c_4648_n 0.0317429f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2868 N_VPWR_M1046_d N_Z_c_4649_n 0.00213438f $X=16.595 $Y=2.955 $X2=0 $Y2=0
cc_2869 N_VPWR_M1070_d N_Z_c_4649_n 0.00236137f $X=17.515 $Y=2.955 $X2=0 $Y2=0
cc_2870 N_VPWR_M1134_d N_Z_c_4649_n 4.10081e-19 $X=18.455 $Y=2.955 $X2=0 $Y2=0
cc_2871 N_VPWR_M1117_s N_Z_c_4649_n 0.00236137f $X=19.455 $Y=2.955 $X2=0 $Y2=0
cc_2872 N_VPWR_M1153_s N_Z_c_4649_n 0.00213438f $X=20.395 $Y=2.955 $X2=0 $Y2=0
cc_2873 N_VPWR_c_3611_n N_Z_c_4649_n 0.0106064f $X=16.72 $Y=3.1 $X2=0 $Y2=0
cc_2874 N_VPWR_c_3613_n N_Z_c_4649_n 0.010348f $X=17.66 $Y=3.1 $X2=0 $Y2=0
cc_2875 N_VPWR_c_3615_n N_Z_c_4649_n 0.0326935f $X=18.63 $Y=3.1 $X2=0 $Y2=0
cc_2876 N_VPWR_c_3617_n N_Z_c_4649_n 0.010348f $X=19.6 $Y=3.1 $X2=0 $Y2=0
cc_2877 N_VPWR_c_3620_n N_Z_c_4649_n 0.0106064f $X=20.54 $Y=3.1 $X2=0 $Y2=0
cc_2878 N_VPWR_c_3661_n N_Z_c_4649_n 0.0317429f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2879 N_VPWR_c_3625_n N_Z_c_4650_n 0.0123133f $X=1.49 $Y=2.72 $X2=0 $Y2=0
cc_2880 N_VPWR_c_3661_n N_Z_c_4650_n 0.0498209f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2881 N_VPWR_c_3628_n N_Z_c_4651_n 0.0123133f $X=4.165 $Y=2.72 $X2=0 $Y2=0
cc_2882 N_VPWR_c_3661_n N_Z_c_4651_n 0.0498209f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2883 N_VPWR_c_3644_n N_Z_c_4652_n 0.0123133f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_2884 N_VPWR_c_3661_n N_Z_c_4652_n 0.0498209f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2885 N_VPWR_c_3630_n N_Z_c_4653_n 0.0123133f $X=10.93 $Y=2.72 $X2=0 $Y2=0
cc_2886 N_VPWR_c_3661_n N_Z_c_4653_n 0.0498209f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2887 N_VPWR_c_3634_n N_Z_c_4654_n 0.0123133f $X=13.91 $Y=2.72 $X2=0 $Y2=0
cc_2888 N_VPWR_c_3661_n N_Z_c_4654_n 0.0498209f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2889 N_VPWR_c_3637_n N_Z_c_4655_n 0.0123133f $X=16.585 $Y=2.72 $X2=0 $Y2=0
cc_2890 N_VPWR_c_3661_n N_Z_c_4655_n 0.0498209f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2891 N_VPWR_c_3648_n N_Z_c_4656_n 0.0123133f $X=20.93 $Y=2.72 $X2=0 $Y2=0
cc_2892 N_VPWR_c_3661_n N_Z_c_4656_n 0.0498209f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2893 N_VPWR_c_3639_n N_Z_c_4657_n 0.0123133f $X=23.35 $Y=2.72 $X2=0 $Y2=0
cc_2894 N_VPWR_c_3661_n N_Z_c_4657_n 0.0498209f $X=24.61 $Y=2.72 $X2=0 $Y2=0
cc_2895 N_VPWR_c_3661_n N_A_1313_297#_M1071_s 0.0011753f $X=24.61 $Y=2.72
+ $X2=-0.19 $Y2=1.305
cc_2896 N_VPWR_c_3661_n N_A_1313_297#_M1118_s 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2897 N_VPWR_M1090_d N_A_1313_297#_c_5507_n 0.00331615f $X=7.035 $Y=1.485
+ $X2=0 $Y2=0
cc_2898 N_VPWR_c_3596_n N_A_1313_297#_c_5507_n 0.0130979f $X=7.18 $Y=2 $X2=0
+ $Y2=0
cc_2899 N_VPWR_M1158_d N_A_1313_297#_c_5502_n 0.00715085f $X=7.975 $Y=1.485
+ $X2=0 $Y2=0
cc_2900 N_VPWR_c_3599_n N_A_1313_297#_c_5502_n 0.0152464f $X=8.12 $Y=2 $X2=0
+ $Y2=0
cc_2901 N_VPWR_c_3596_n N_A_1313_297#_c_5520_n 0.0153177f $X=7.18 $Y=2 $X2=0
+ $Y2=0
cc_2902 N_VPWR_c_3598_n N_A_1313_297#_c_5520_n 8.30334e-19 $X=7.985 $Y=2.72
+ $X2=0 $Y2=0
cc_2903 N_VPWR_c_3643_n N_A_1313_297#_c_5520_n 8.30334e-19 $X=7.045 $Y=2.72
+ $X2=0 $Y2=0
cc_2904 N_VPWR_c_3661_n N_A_1313_297#_c_5520_n 0.0558368f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2905 N_VPWR_c_3594_n N_A_1313_297#_c_5555_n 0.00170069f $X=6.21 $Y=1.66 $X2=0
+ $Y2=0
cc_2906 N_VPWR_c_3596_n N_A_1313_297#_c_5555_n 6.68271e-19 $X=7.18 $Y=2 $X2=0
+ $Y2=0
cc_2907 N_VPWR_c_3661_n N_A_1313_297#_c_5555_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2908 N_VPWR_c_3598_n N_A_1313_297#_c_5503_n 8.30334e-19 $X=7.985 $Y=2.72
+ $X2=0 $Y2=0
cc_2909 N_VPWR_c_3599_n N_A_1313_297#_c_5503_n 0.0156478f $X=8.12 $Y=2 $X2=0
+ $Y2=0
cc_2910 N_VPWR_c_3644_n N_A_1313_297#_c_5503_n 0.00115812f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_2911 N_VPWR_c_3661_n N_A_1313_297#_c_5503_n 0.0605692f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2912 N_VPWR_c_3596_n N_A_1313_297#_c_5562_n 6.68271e-19 $X=7.18 $Y=2 $X2=0
+ $Y2=0
cc_2913 N_VPWR_c_3599_n N_A_1313_297#_c_5562_n 6.68271e-19 $X=8.12 $Y=2 $X2=0
+ $Y2=0
cc_2914 N_VPWR_c_3661_n N_A_1313_297#_c_5562_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2915 N_VPWR_c_3661_n N_A_1313_297#_c_5531_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2916 N_VPWR_c_3599_n N_A_1313_297#_c_5566_n 6.69936e-19 $X=8.12 $Y=2 $X2=0
+ $Y2=0
cc_2917 N_VPWR_c_3661_n N_A_1313_297#_c_5566_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2918 N_VPWR_c_3661_n N_A_1313_297#_c_5533_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2919 N_VPWR_c_3661_n N_A_1313_297#_c_5569_n 0.0296491f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2920 N_VPWR_c_3594_n N_A_1313_297#_c_5523_n 0.031816f $X=6.21 $Y=1.66 $X2=0
+ $Y2=0
cc_2921 N_VPWR_c_3596_n N_A_1313_297#_c_5523_n 0.0268237f $X=7.18 $Y=2 $X2=0
+ $Y2=0
cc_2922 N_VPWR_c_3643_n N_A_1313_297#_c_5523_n 0.0189467f $X=7.045 $Y=2.72 $X2=0
+ $Y2=0
cc_2923 N_VPWR_c_3661_n N_A_1313_297#_c_5523_n 0.00313104f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_2924 N_VPWR_c_3596_n N_A_1313_297#_c_5526_n 0.0268237f $X=7.18 $Y=2 $X2=0
+ $Y2=0
cc_2925 N_VPWR_c_3598_n N_A_1313_297#_c_5526_n 0.0189467f $X=7.985 $Y=2.72 $X2=0
+ $Y2=0
cc_2926 N_VPWR_c_3599_n N_A_1313_297#_c_5526_n 0.0268237f $X=8.12 $Y=2 $X2=0
+ $Y2=0
cc_2927 N_VPWR_c_3661_n N_A_1313_297#_c_5526_n 0.00300637f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_2928 N_VPWR_c_3601_n N_A_1313_297#_c_5578_n 0.00167067f $X=11.095 $Y=1.77
+ $X2=0 $Y2=0
cc_2929 N_VPWR_c_3661_n N_A_1313_297#_c_5578_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2930 N_VPWR_c_3599_n N_A_1313_297#_c_5504_n 0.0390576f $X=8.12 $Y=2 $X2=0
+ $Y2=0
cc_2931 N_VPWR_c_3644_n N_A_1313_297#_c_5504_n 0.0213652f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_2932 N_VPWR_c_3661_n N_A_1313_297#_c_5504_n 0.0027766f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2933 N_VPWR_c_3661_n N_A_1313_297#_c_5505_n 0.00468575f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_2934 N_VPWR_c_3601_n N_A_1313_297#_c_5506_n 0.0505494f $X=11.095 $Y=1.77
+ $X2=0 $Y2=0
cc_2935 N_VPWR_c_3630_n N_A_1313_297#_c_5506_n 0.0213652f $X=10.93 $Y=2.72 $X2=0
+ $Y2=0
cc_2936 N_VPWR_c_3661_n N_A_1313_297#_c_5506_n 0.00284741f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_2937 N_VPWR_c_3661_n N_A_1313_591#_M1000_d 0.0011753f $X=24.61 $Y=2.72
+ $X2=-0.19 $Y2=1.305
cc_2938 N_VPWR_c_3661_n N_A_1313_591#_M1095_d 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2939 N_VPWR_M1076_s N_A_1313_591#_c_5635_n 0.00331615f $X=7.035 $Y=2.955
+ $X2=0 $Y2=0
cc_2940 N_VPWR_c_3597_n N_A_1313_591#_c_5635_n 0.0130979f $X=7.18 $Y=3.1 $X2=0
+ $Y2=0
cc_2941 N_VPWR_M1120_s N_A_1313_591#_c_5630_n 0.00715085f $X=7.975 $Y=2.955
+ $X2=0 $Y2=0
cc_2942 N_VPWR_c_3600_n N_A_1313_591#_c_5630_n 0.0152464f $X=8.12 $Y=3.1 $X2=0
+ $Y2=0
cc_2943 N_VPWR_c_3597_n N_A_1313_591#_c_5648_n 0.0153177f $X=7.18 $Y=3.1 $X2=0
+ $Y2=0
cc_2944 N_VPWR_c_3598_n N_A_1313_591#_c_5648_n 8.30334e-19 $X=7.985 $Y=2.72
+ $X2=0 $Y2=0
cc_2945 N_VPWR_c_3643_n N_A_1313_591#_c_5648_n 8.30334e-19 $X=7.045 $Y=2.72
+ $X2=0 $Y2=0
cc_2946 N_VPWR_c_3661_n N_A_1313_591#_c_5648_n 0.0558368f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2947 N_VPWR_c_3595_n N_A_1313_591#_c_5683_n 0.00170069f $X=6.21 $Y=3.1 $X2=0
+ $Y2=0
cc_2948 N_VPWR_c_3597_n N_A_1313_591#_c_5683_n 6.68271e-19 $X=7.18 $Y=3.1 $X2=0
+ $Y2=0
cc_2949 N_VPWR_c_3661_n N_A_1313_591#_c_5683_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2950 N_VPWR_c_3598_n N_A_1313_591#_c_5631_n 8.30334e-19 $X=7.985 $Y=2.72
+ $X2=0 $Y2=0
cc_2951 N_VPWR_c_3600_n N_A_1313_591#_c_5631_n 0.0156478f $X=8.12 $Y=3.1 $X2=0
+ $Y2=0
cc_2952 N_VPWR_c_3644_n N_A_1313_591#_c_5631_n 0.00115812f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_2953 N_VPWR_c_3661_n N_A_1313_591#_c_5631_n 0.0605692f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2954 N_VPWR_c_3597_n N_A_1313_591#_c_5690_n 6.68271e-19 $X=7.18 $Y=3.1 $X2=0
+ $Y2=0
cc_2955 N_VPWR_c_3600_n N_A_1313_591#_c_5690_n 6.68271e-19 $X=8.12 $Y=3.1 $X2=0
+ $Y2=0
cc_2956 N_VPWR_c_3661_n N_A_1313_591#_c_5690_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2957 N_VPWR_c_3661_n N_A_1313_591#_c_5659_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2958 N_VPWR_c_3600_n N_A_1313_591#_c_5694_n 6.69936e-19 $X=8.12 $Y=3.1 $X2=0
+ $Y2=0
cc_2959 N_VPWR_c_3661_n N_A_1313_591#_c_5694_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2960 N_VPWR_c_3661_n N_A_1313_591#_c_5661_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2961 N_VPWR_c_3661_n N_A_1313_591#_c_5697_n 0.0296491f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2962 N_VPWR_c_3602_n N_A_1313_591#_c_5698_n 0.00167067f $X=11.095 $Y=3.14
+ $X2=0 $Y2=0
cc_2963 N_VPWR_c_3661_n N_A_1313_591#_c_5698_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2964 N_VPWR_c_3595_n N_A_1313_591#_c_5651_n 0.031816f $X=6.21 $Y=3.1 $X2=0
+ $Y2=0
cc_2965 N_VPWR_c_3597_n N_A_1313_591#_c_5651_n 0.0268237f $X=7.18 $Y=3.1 $X2=0
+ $Y2=0
cc_2966 N_VPWR_c_3643_n N_A_1313_591#_c_5651_n 0.0189467f $X=7.045 $Y=2.72 $X2=0
+ $Y2=0
cc_2967 N_VPWR_c_3661_n N_A_1313_591#_c_5651_n 0.00313104f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_2968 N_VPWR_c_3597_n N_A_1313_591#_c_5654_n 0.0268237f $X=7.18 $Y=3.1 $X2=0
+ $Y2=0
cc_2969 N_VPWR_c_3598_n N_A_1313_591#_c_5654_n 0.0189467f $X=7.985 $Y=2.72 $X2=0
+ $Y2=0
cc_2970 N_VPWR_c_3600_n N_A_1313_591#_c_5654_n 0.0268237f $X=8.12 $Y=3.1 $X2=0
+ $Y2=0
cc_2971 N_VPWR_c_3661_n N_A_1313_591#_c_5654_n 0.00300637f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_2972 N_VPWR_c_3600_n N_A_1313_591#_c_5632_n 0.0390576f $X=8.12 $Y=3.1 $X2=0
+ $Y2=0
cc_2973 N_VPWR_c_3644_n N_A_1313_591#_c_5632_n 0.0213652f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_2974 N_VPWR_c_3661_n N_A_1313_591#_c_5632_n 0.0027766f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2975 N_VPWR_c_3661_n N_A_1313_591#_c_5633_n 0.00468575f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_2976 N_VPWR_c_3602_n N_A_1313_591#_c_5634_n 0.0505494f $X=11.095 $Y=3.14
+ $X2=0 $Y2=0
cc_2977 N_VPWR_c_3630_n N_A_1313_591#_c_5634_n 0.0213652f $X=10.93 $Y=2.72 $X2=0
+ $Y2=0
cc_2978 N_VPWR_c_3661_n N_A_1313_591#_c_5634_n 0.00284741f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_2979 N_VPWR_c_3661_n N_A_2839_311#_M1042_s 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2980 N_VPWR_c_3661_n N_A_2839_311#_M1105_s 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2981 N_VPWR_M1042_d N_A_2839_311#_c_5758_n 0.00715085f $X=16.595 $Y=1.485
+ $X2=0 $Y2=0
cc_2982 N_VPWR_c_3610_n N_A_2839_311#_c_5758_n 0.0152464f $X=16.72 $Y=2 $X2=0
+ $Y2=0
cc_2983 N_VPWR_M1062_d N_A_2839_311#_c_5780_n 0.00331615f $X=17.515 $Y=1.485
+ $X2=0 $Y2=0
cc_2984 N_VPWR_c_3612_n N_A_2839_311#_c_5780_n 0.0130979f $X=17.66 $Y=2 $X2=0
+ $Y2=0
cc_2985 N_VPWR_c_3661_n N_A_2839_311#_c_5767_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2986 N_VPWR_c_3608_n N_A_2839_311#_c_5809_n 0.00167067f $X=13.745 $Y=1.77
+ $X2=0 $Y2=0
cc_2987 N_VPWR_c_3661_n N_A_2839_311#_c_5809_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2988 N_VPWR_c_3661_n N_A_2839_311#_c_5769_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2989 N_VPWR_c_3661_n N_A_2839_311#_c_5812_n 0.0296491f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2990 N_VPWR_c_3610_n N_A_2839_311#_c_5760_n 0.0156478f $X=16.72 $Y=2 $X2=0
+ $Y2=0
cc_2991 N_VPWR_c_3637_n N_A_2839_311#_c_5760_n 0.00115812f $X=16.585 $Y=2.72
+ $X2=0 $Y2=0
cc_2992 N_VPWR_c_3645_n N_A_2839_311#_c_5760_n 8.30334e-19 $X=17.525 $Y=2.72
+ $X2=0 $Y2=0
cc_2993 N_VPWR_c_3661_n N_A_2839_311#_c_5760_n 0.0605692f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2994 N_VPWR_c_3610_n N_A_2839_311#_c_5817_n 6.69936e-19 $X=16.72 $Y=2 $X2=0
+ $Y2=0
cc_2995 N_VPWR_c_3661_n N_A_2839_311#_c_5817_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_2996 N_VPWR_c_3612_n N_A_2839_311#_c_5793_n 0.0153177f $X=17.66 $Y=2 $X2=0
+ $Y2=0
cc_2997 N_VPWR_c_3645_n N_A_2839_311#_c_5793_n 8.30334e-19 $X=17.525 $Y=2.72
+ $X2=0 $Y2=0
cc_2998 N_VPWR_c_3646_n N_A_2839_311#_c_5793_n 8.30334e-19 $X=18.465 $Y=2.72
+ $X2=0 $Y2=0
cc_2999 N_VPWR_c_3661_n N_A_2839_311#_c_5793_n 0.0558368f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3000 N_VPWR_c_3610_n N_A_2839_311#_c_5823_n 6.68271e-19 $X=16.72 $Y=2 $X2=0
+ $Y2=0
cc_3001 N_VPWR_c_3612_n N_A_2839_311#_c_5823_n 6.68271e-19 $X=17.66 $Y=2 $X2=0
+ $Y2=0
cc_3002 N_VPWR_c_3661_n N_A_2839_311#_c_5823_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3003 N_VPWR_c_3610_n N_A_2839_311#_c_5795_n 0.0268237f $X=16.72 $Y=2 $X2=0
+ $Y2=0
cc_3004 N_VPWR_c_3612_n N_A_2839_311#_c_5795_n 0.0268237f $X=17.66 $Y=2 $X2=0
+ $Y2=0
cc_3005 N_VPWR_c_3645_n N_A_2839_311#_c_5795_n 0.0189467f $X=17.525 $Y=2.72
+ $X2=0 $Y2=0
cc_3006 N_VPWR_c_3661_n N_A_2839_311#_c_5795_n 0.00300637f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3007 N_VPWR_c_3612_n N_A_2839_311#_c_5830_n 6.68271e-19 $X=17.66 $Y=2 $X2=0
+ $Y2=0
cc_3008 N_VPWR_c_3614_n N_A_2839_311#_c_5830_n 0.00170069f $X=18.63 $Y=1.66
+ $X2=0 $Y2=0
cc_3009 N_VPWR_c_3661_n N_A_2839_311#_c_5830_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3010 N_VPWR_c_3612_n N_A_2839_311#_c_5798_n 0.0268237f $X=17.66 $Y=2 $X2=0
+ $Y2=0
cc_3011 N_VPWR_c_3614_n N_A_2839_311#_c_5798_n 0.031816f $X=18.63 $Y=1.66 $X2=0
+ $Y2=0
cc_3012 N_VPWR_c_3646_n N_A_2839_311#_c_5798_n 0.0189467f $X=18.465 $Y=2.72
+ $X2=0 $Y2=0
cc_3013 N_VPWR_c_3661_n N_A_2839_311#_c_5798_n 0.00313104f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3014 N_VPWR_c_3608_n N_A_2839_311#_c_5761_n 0.0505494f $X=13.745 $Y=1.77
+ $X2=0 $Y2=0
cc_3015 N_VPWR_c_3634_n N_A_2839_311#_c_5761_n 0.0213652f $X=13.91 $Y=2.72 $X2=0
+ $Y2=0
cc_3016 N_VPWR_c_3661_n N_A_2839_311#_c_5761_n 0.00284741f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3017 N_VPWR_c_3661_n N_A_2839_311#_c_5762_n 0.00468575f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3018 N_VPWR_c_3610_n N_A_2839_311#_c_5763_n 0.0390576f $X=16.72 $Y=2 $X2=0
+ $Y2=0
cc_3019 N_VPWR_c_3637_n N_A_2839_311#_c_5763_n 0.0213652f $X=16.585 $Y=2.72
+ $X2=0 $Y2=0
cc_3020 N_VPWR_c_3661_n N_A_2839_311#_c_5763_n 0.0027766f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3021 N_VPWR_c_3661_n N_A_2839_613#_M1046_s 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3022 N_VPWR_c_3661_n N_A_2839_613#_M1113_s 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3023 N_VPWR_M1046_d N_A_2839_613#_c_5889_n 0.00715085f $X=16.595 $Y=2.955
+ $X2=0 $Y2=0
cc_3024 N_VPWR_c_3611_n N_A_2839_613#_c_5889_n 0.0152464f $X=16.72 $Y=3.1 $X2=0
+ $Y2=0
cc_3025 N_VPWR_M1070_d N_A_2839_613#_c_5911_n 0.00331615f $X=17.515 $Y=2.955
+ $X2=0 $Y2=0
cc_3026 N_VPWR_c_3613_n N_A_2839_613#_c_5911_n 0.0130979f $X=17.66 $Y=3.1 $X2=0
+ $Y2=0
cc_3027 N_VPWR_c_3661_n N_A_2839_613#_c_5898_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3028 N_VPWR_c_3609_n N_A_2839_613#_c_5940_n 0.00167067f $X=13.745 $Y=3.14
+ $X2=0 $Y2=0
cc_3029 N_VPWR_c_3661_n N_A_2839_613#_c_5940_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3030 N_VPWR_c_3661_n N_A_2839_613#_c_5900_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3031 N_VPWR_c_3661_n N_A_2839_613#_c_5943_n 0.0296491f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3032 N_VPWR_c_3611_n N_A_2839_613#_c_5891_n 0.0156478f $X=16.72 $Y=3.1 $X2=0
+ $Y2=0
cc_3033 N_VPWR_c_3637_n N_A_2839_613#_c_5891_n 0.00115812f $X=16.585 $Y=2.72
+ $X2=0 $Y2=0
cc_3034 N_VPWR_c_3645_n N_A_2839_613#_c_5891_n 8.30334e-19 $X=17.525 $Y=2.72
+ $X2=0 $Y2=0
cc_3035 N_VPWR_c_3661_n N_A_2839_613#_c_5891_n 0.0605692f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3036 N_VPWR_c_3611_n N_A_2839_613#_c_5948_n 6.69936e-19 $X=16.72 $Y=3.1 $X2=0
+ $Y2=0
cc_3037 N_VPWR_c_3661_n N_A_2839_613#_c_5948_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3038 N_VPWR_c_3613_n N_A_2839_613#_c_5924_n 0.0153177f $X=17.66 $Y=3.1 $X2=0
+ $Y2=0
cc_3039 N_VPWR_c_3645_n N_A_2839_613#_c_5924_n 8.30334e-19 $X=17.525 $Y=2.72
+ $X2=0 $Y2=0
cc_3040 N_VPWR_c_3646_n N_A_2839_613#_c_5924_n 8.30334e-19 $X=18.465 $Y=2.72
+ $X2=0 $Y2=0
cc_3041 N_VPWR_c_3661_n N_A_2839_613#_c_5924_n 0.0558368f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3042 N_VPWR_c_3611_n N_A_2839_613#_c_5954_n 6.68271e-19 $X=16.72 $Y=3.1 $X2=0
+ $Y2=0
cc_3043 N_VPWR_c_3613_n N_A_2839_613#_c_5954_n 6.68271e-19 $X=17.66 $Y=3.1 $X2=0
+ $Y2=0
cc_3044 N_VPWR_c_3661_n N_A_2839_613#_c_5954_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3045 N_VPWR_c_3613_n N_A_2839_613#_c_5957_n 6.68271e-19 $X=17.66 $Y=3.1 $X2=0
+ $Y2=0
cc_3046 N_VPWR_c_3615_n N_A_2839_613#_c_5957_n 0.00170069f $X=18.63 $Y=3.1 $X2=0
+ $Y2=0
cc_3047 N_VPWR_c_3661_n N_A_2839_613#_c_5957_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3048 N_VPWR_c_3609_n N_A_2839_613#_c_5892_n 0.0505494f $X=13.745 $Y=3.14
+ $X2=0 $Y2=0
cc_3049 N_VPWR_c_3634_n N_A_2839_613#_c_5892_n 0.0213652f $X=13.91 $Y=2.72 $X2=0
+ $Y2=0
cc_3050 N_VPWR_c_3661_n N_A_2839_613#_c_5892_n 0.00284741f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3051 N_VPWR_c_3661_n N_A_2839_613#_c_5893_n 0.00468575f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3052 N_VPWR_c_3611_n N_A_2839_613#_c_5894_n 0.0390576f $X=16.72 $Y=3.1 $X2=0
+ $Y2=0
cc_3053 N_VPWR_c_3637_n N_A_2839_613#_c_5894_n 0.0213652f $X=16.585 $Y=2.72
+ $X2=0 $Y2=0
cc_3054 N_VPWR_c_3661_n N_A_2839_613#_c_5894_n 0.0027766f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3055 N_VPWR_c_3611_n N_A_2839_613#_c_5927_n 0.0268237f $X=16.72 $Y=3.1 $X2=0
+ $Y2=0
cc_3056 N_VPWR_c_3613_n N_A_2839_613#_c_5927_n 0.0268237f $X=17.66 $Y=3.1 $X2=0
+ $Y2=0
cc_3057 N_VPWR_c_3645_n N_A_2839_613#_c_5927_n 0.0189467f $X=17.525 $Y=2.72
+ $X2=0 $Y2=0
cc_3058 N_VPWR_c_3661_n N_A_2839_613#_c_5927_n 0.00300637f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3059 N_VPWR_c_3613_n N_A_2839_613#_c_5930_n 0.0268237f $X=17.66 $Y=3.1 $X2=0
+ $Y2=0
cc_3060 N_VPWR_c_3615_n N_A_2839_613#_c_5930_n 0.031816f $X=18.63 $Y=3.1 $X2=0
+ $Y2=0
cc_3061 N_VPWR_c_3646_n N_A_2839_613#_c_5930_n 0.0189467f $X=18.465 $Y=2.72
+ $X2=0 $Y2=0
cc_3062 N_VPWR_c_3661_n N_A_2839_613#_c_5930_n 0.00313104f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3063 N_VPWR_c_3661_n N_A_3797_297#_M1082_d 0.0011753f $X=24.61 $Y=2.72
+ $X2=-0.19 $Y2=1.305
cc_3064 N_VPWR_c_3661_n N_A_3797_297#_M1130_d 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3065 N_VPWR_M1108_s N_A_3797_297#_c_6025_n 0.00331615f $X=19.455 $Y=1.485
+ $X2=0 $Y2=0
cc_3066 N_VPWR_c_3616_n N_A_3797_297#_c_6025_n 0.0130979f $X=19.6 $Y=2 $X2=0
+ $Y2=0
cc_3067 N_VPWR_M1145_s N_A_3797_297#_c_6020_n 0.00715085f $X=20.395 $Y=1.485
+ $X2=0 $Y2=0
cc_3068 N_VPWR_c_3619_n N_A_3797_297#_c_6020_n 0.0152464f $X=20.54 $Y=2 $X2=0
+ $Y2=0
cc_3069 N_VPWR_c_3616_n N_A_3797_297#_c_6038_n 0.0153177f $X=19.6 $Y=2 $X2=0
+ $Y2=0
cc_3070 N_VPWR_c_3618_n N_A_3797_297#_c_6038_n 8.30334e-19 $X=20.405 $Y=2.72
+ $X2=0 $Y2=0
cc_3071 N_VPWR_c_3647_n N_A_3797_297#_c_6038_n 8.30334e-19 $X=19.465 $Y=2.72
+ $X2=0 $Y2=0
cc_3072 N_VPWR_c_3661_n N_A_3797_297#_c_6038_n 0.0558368f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3073 N_VPWR_c_3614_n N_A_3797_297#_c_6073_n 0.00170069f $X=18.63 $Y=1.66
+ $X2=0 $Y2=0
cc_3074 N_VPWR_c_3616_n N_A_3797_297#_c_6073_n 6.68271e-19 $X=19.6 $Y=2 $X2=0
+ $Y2=0
cc_3075 N_VPWR_c_3661_n N_A_3797_297#_c_6073_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3076 N_VPWR_c_3618_n N_A_3797_297#_c_6021_n 8.30334e-19 $X=20.405 $Y=2.72
+ $X2=0 $Y2=0
cc_3077 N_VPWR_c_3619_n N_A_3797_297#_c_6021_n 0.0156478f $X=20.54 $Y=2 $X2=0
+ $Y2=0
cc_3078 N_VPWR_c_3648_n N_A_3797_297#_c_6021_n 0.00115812f $X=20.93 $Y=2.72
+ $X2=0 $Y2=0
cc_3079 N_VPWR_c_3661_n N_A_3797_297#_c_6021_n 0.0605692f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3080 N_VPWR_c_3616_n N_A_3797_297#_c_6080_n 6.68271e-19 $X=19.6 $Y=2 $X2=0
+ $Y2=0
cc_3081 N_VPWR_c_3619_n N_A_3797_297#_c_6080_n 6.68271e-19 $X=20.54 $Y=2 $X2=0
+ $Y2=0
cc_3082 N_VPWR_c_3661_n N_A_3797_297#_c_6080_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3083 N_VPWR_c_3661_n N_A_3797_297#_c_6049_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3084 N_VPWR_c_3619_n N_A_3797_297#_c_6084_n 6.69936e-19 $X=20.54 $Y=2 $X2=0
+ $Y2=0
cc_3085 N_VPWR_c_3661_n N_A_3797_297#_c_6084_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3086 N_VPWR_c_3661_n N_A_3797_297#_c_6051_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3087 N_VPWR_c_3661_n N_A_3797_297#_c_6087_n 0.0296491f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3088 N_VPWR_c_3614_n N_A_3797_297#_c_6041_n 0.031816f $X=18.63 $Y=1.66 $X2=0
+ $Y2=0
cc_3089 N_VPWR_c_3616_n N_A_3797_297#_c_6041_n 0.0268237f $X=19.6 $Y=2 $X2=0
+ $Y2=0
cc_3090 N_VPWR_c_3647_n N_A_3797_297#_c_6041_n 0.0189467f $X=19.465 $Y=2.72
+ $X2=0 $Y2=0
cc_3091 N_VPWR_c_3661_n N_A_3797_297#_c_6041_n 0.00313104f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3092 N_VPWR_c_3616_n N_A_3797_297#_c_6044_n 0.0268237f $X=19.6 $Y=2 $X2=0
+ $Y2=0
cc_3093 N_VPWR_c_3618_n N_A_3797_297#_c_6044_n 0.0189467f $X=20.405 $Y=2.72
+ $X2=0 $Y2=0
cc_3094 N_VPWR_c_3619_n N_A_3797_297#_c_6044_n 0.0268237f $X=20.54 $Y=2 $X2=0
+ $Y2=0
cc_3095 N_VPWR_c_3661_n N_A_3797_297#_c_6044_n 0.00300637f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3096 N_VPWR_c_3621_n N_A_3797_297#_c_6096_n 0.00167067f $X=23.515 $Y=1.77
+ $X2=0 $Y2=0
cc_3097 N_VPWR_c_3661_n N_A_3797_297#_c_6096_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3098 N_VPWR_c_3619_n N_A_3797_297#_c_6022_n 0.0390576f $X=20.54 $Y=2 $X2=0
+ $Y2=0
cc_3099 N_VPWR_c_3648_n N_A_3797_297#_c_6022_n 0.0213652f $X=20.93 $Y=2.72 $X2=0
+ $Y2=0
cc_3100 N_VPWR_c_3661_n N_A_3797_297#_c_6022_n 0.0027766f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3101 N_VPWR_c_3661_n N_A_3797_297#_c_6023_n 0.00468575f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3102 N_VPWR_c_3621_n N_A_3797_297#_c_6024_n 0.0523777f $X=23.515 $Y=1.77
+ $X2=0 $Y2=0
cc_3103 N_VPWR_c_3639_n N_A_3797_297#_c_6024_n 0.0213652f $X=23.35 $Y=2.72 $X2=0
+ $Y2=0
cc_3104 N_VPWR_c_3661_n N_A_3797_297#_c_6024_n 0.00302891f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3105 N_VPWR_c_3661_n N_A_3797_591#_M1087_d 0.0011753f $X=24.61 $Y=2.72
+ $X2=-0.19 $Y2=1.305
cc_3106 N_VPWR_c_3661_n N_A_3797_591#_M1139_d 0.0011753f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3107 N_VPWR_M1117_s N_A_3797_591#_c_6147_n 0.00331615f $X=19.455 $Y=2.955
+ $X2=0 $Y2=0
cc_3108 N_VPWR_c_3617_n N_A_3797_591#_c_6147_n 0.0130979f $X=19.6 $Y=3.1 $X2=0
+ $Y2=0
cc_3109 N_VPWR_M1153_s N_A_3797_591#_c_6142_n 0.00715085f $X=20.395 $Y=2.955
+ $X2=0 $Y2=0
cc_3110 N_VPWR_c_3620_n N_A_3797_591#_c_6142_n 0.0152464f $X=20.54 $Y=3.1 $X2=0
+ $Y2=0
cc_3111 N_VPWR_c_3617_n N_A_3797_591#_c_6160_n 0.0153177f $X=19.6 $Y=3.1 $X2=0
+ $Y2=0
cc_3112 N_VPWR_c_3618_n N_A_3797_591#_c_6160_n 8.30334e-19 $X=20.405 $Y=2.72
+ $X2=0 $Y2=0
cc_3113 N_VPWR_c_3647_n N_A_3797_591#_c_6160_n 8.30334e-19 $X=19.465 $Y=2.72
+ $X2=0 $Y2=0
cc_3114 N_VPWR_c_3661_n N_A_3797_591#_c_6160_n 0.0558368f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3115 N_VPWR_c_3615_n N_A_3797_591#_c_6195_n 0.00170069f $X=18.63 $Y=3.1 $X2=0
+ $Y2=0
cc_3116 N_VPWR_c_3617_n N_A_3797_591#_c_6195_n 6.68271e-19 $X=19.6 $Y=3.1 $X2=0
+ $Y2=0
cc_3117 N_VPWR_c_3661_n N_A_3797_591#_c_6195_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3118 N_VPWR_c_3618_n N_A_3797_591#_c_6143_n 8.30334e-19 $X=20.405 $Y=2.72
+ $X2=0 $Y2=0
cc_3119 N_VPWR_c_3620_n N_A_3797_591#_c_6143_n 0.0156478f $X=20.54 $Y=3.1 $X2=0
+ $Y2=0
cc_3120 N_VPWR_c_3648_n N_A_3797_591#_c_6143_n 0.00115812f $X=20.93 $Y=2.72
+ $X2=0 $Y2=0
cc_3121 N_VPWR_c_3661_n N_A_3797_591#_c_6143_n 0.0605692f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3122 N_VPWR_c_3617_n N_A_3797_591#_c_6202_n 6.68271e-19 $X=19.6 $Y=3.1 $X2=0
+ $Y2=0
cc_3123 N_VPWR_c_3620_n N_A_3797_591#_c_6202_n 6.68271e-19 $X=20.54 $Y=3.1 $X2=0
+ $Y2=0
cc_3124 N_VPWR_c_3661_n N_A_3797_591#_c_6202_n 0.0295747f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3125 N_VPWR_c_3661_n N_A_3797_591#_c_6171_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3126 N_VPWR_c_3620_n N_A_3797_591#_c_6206_n 6.69936e-19 $X=20.54 $Y=3.1 $X2=0
+ $Y2=0
cc_3127 N_VPWR_c_3661_n N_A_3797_591#_c_6206_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3128 N_VPWR_c_3661_n N_A_3797_591#_c_6173_n 0.0571367f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3129 N_VPWR_c_3661_n N_A_3797_591#_c_6209_n 0.0296491f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3130 N_VPWR_c_3622_n N_A_3797_591#_c_6210_n 0.00167067f $X=23.515 $Y=3.14
+ $X2=0 $Y2=0
cc_3131 N_VPWR_c_3661_n N_A_3797_591#_c_6210_n 0.0297857f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3132 N_VPWR_c_3615_n N_A_3797_591#_c_6163_n 0.031816f $X=18.63 $Y=3.1 $X2=0
+ $Y2=0
cc_3133 N_VPWR_c_3617_n N_A_3797_591#_c_6163_n 0.0268237f $X=19.6 $Y=3.1 $X2=0
+ $Y2=0
cc_3134 N_VPWR_c_3647_n N_A_3797_591#_c_6163_n 0.0189467f $X=19.465 $Y=2.72
+ $X2=0 $Y2=0
cc_3135 N_VPWR_c_3661_n N_A_3797_591#_c_6163_n 0.00313104f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3136 N_VPWR_c_3617_n N_A_3797_591#_c_6166_n 0.0268237f $X=19.6 $Y=3.1 $X2=0
+ $Y2=0
cc_3137 N_VPWR_c_3618_n N_A_3797_591#_c_6166_n 0.0189467f $X=20.405 $Y=2.72
+ $X2=0 $Y2=0
cc_3138 N_VPWR_c_3620_n N_A_3797_591#_c_6166_n 0.0268237f $X=20.54 $Y=3.1 $X2=0
+ $Y2=0
cc_3139 N_VPWR_c_3661_n N_A_3797_591#_c_6166_n 0.00300637f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3140 N_VPWR_c_3620_n N_A_3797_591#_c_6144_n 0.0390576f $X=20.54 $Y=3.1 $X2=0
+ $Y2=0
cc_3141 N_VPWR_c_3648_n N_A_3797_591#_c_6144_n 0.0213652f $X=20.93 $Y=2.72 $X2=0
+ $Y2=0
cc_3142 N_VPWR_c_3661_n N_A_3797_591#_c_6144_n 0.0027766f $X=24.61 $Y=2.72 $X2=0
+ $Y2=0
cc_3143 N_VPWR_c_3661_n N_A_3797_591#_c_6145_n 0.00468575f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3144 N_VPWR_c_3622_n N_A_3797_591#_c_6146_n 0.0523777f $X=23.515 $Y=3.14
+ $X2=0 $Y2=0
cc_3145 N_VPWR_c_3639_n N_A_3797_591#_c_6146_n 0.0213652f $X=23.35 $Y=2.72 $X2=0
+ $Y2=0
cc_3146 N_VPWR_c_3661_n N_A_3797_591#_c_6146_n 0.00302891f $X=24.61 $Y=2.72
+ $X2=0 $Y2=0
cc_3147 N_VPWR_c_3594_n N_VGND_c_6274_n 0.00950712f $X=6.21 $Y=1.66 $X2=0 $Y2=0
cc_3148 N_VPWR_c_3595_n N_VGND_c_6275_n 0.00950712f $X=6.21 $Y=3.1 $X2=0 $Y2=0
cc_3149 N_VPWR_c_3614_n N_VGND_c_6294_n 0.00950712f $X=18.63 $Y=1.66 $X2=0 $Y2=0
cc_3150 N_VPWR_c_3615_n N_VGND_c_6295_n 0.00950712f $X=18.63 $Y=3.1 $X2=0 $Y2=0
cc_3151 N_A_355_311#_c_4338_n N_A_355_613#_c_4465_n 0.00460759f $X=2.84 $Y=1.7
+ $X2=0 $Y2=0
cc_3152 N_A_355_311#_c_4338_n N_Z_c_4590_n 0.0192125f $X=2.84 $Y=1.7 $X2=0 $Y2=0
cc_3153 N_A_355_311#_c_4338_n N_Z_c_4608_n 0.0024794f $X=2.84 $Y=1.7 $X2=0 $Y2=0
cc_3154 N_A_355_311#_M1147_d N_Z_c_4644_n 2.15519e-19 $X=3.635 $Y=1.555 $X2=0
+ $Y2=0
cc_3155 N_A_355_311#_c_4334_n N_Z_c_4644_n 0.0242319f $X=4.605 $Y=1.58 $X2=0
+ $Y2=0
cc_3156 N_A_355_311#_c_4356_n N_Z_c_4644_n 0.020688f $X=5.545 $Y=1.58 $X2=0
+ $Y2=0
cc_3157 N_A_355_311#_c_4345_n N_Z_c_4644_n 0.0146113f $X=3.645 $Y=2.225 $X2=0
+ $Y2=0
cc_3158 N_A_355_311#_c_4336_n N_Z_c_4644_n 0.0521734f $X=4.625 $Y=2.225 $X2=0
+ $Y2=0
cc_3159 N_A_355_311#_c_4393_n N_Z_c_4644_n 0.0238046f $X=3.935 $Y=2.225 $X2=0
+ $Y2=0
cc_3160 N_A_355_311#_c_4369_n N_Z_c_4644_n 0.0481433f $X=5.565 $Y=2.225 $X2=0
+ $Y2=0
cc_3161 N_A_355_311#_c_4399_n N_Z_c_4644_n 0.0238869f $X=4.915 $Y=2.225 $X2=0
+ $Y2=0
cc_3162 N_A_355_311#_c_4371_n N_Z_c_4644_n 0.0205035f $X=4.77 $Y=2.225 $X2=0
+ $Y2=0
cc_3163 N_A_355_311#_c_4406_n N_Z_c_4644_n 0.0238869f $X=5.71 $Y=2.225 $X2=0
+ $Y2=0
cc_3164 N_A_355_311#_c_4374_n N_Z_c_4644_n 0.0187608f $X=5.71 $Y=2.225 $X2=0
+ $Y2=0
cc_3165 N_A_355_311#_c_4339_n N_Z_c_4644_n 0.026602f $X=3.78 $Y=1.7 $X2=0 $Y2=0
cc_3166 N_A_355_311#_c_4345_n N_Z_c_5128_n 0.0238869f $X=3.645 $Y=2.225 $X2=0
+ $Y2=0
cc_3167 N_A_355_311#_c_4338_n N_Z_c_5128_n 6.68271e-19 $X=2.84 $Y=1.7 $X2=0
+ $Y2=0
cc_3168 N_A_355_311#_c_4339_n N_Z_c_5128_n 6.74054e-19 $X=3.78 $Y=1.7 $X2=0
+ $Y2=0
cc_3169 N_A_355_311#_M1019_d N_Z_c_4693_n 3.28377e-19 $X=2.695 $Y=1.555 $X2=0
+ $Y2=0
cc_3170 N_A_355_311#_c_4343_n N_Z_c_4693_n 0.0139315f $X=2.695 $Y=2.225 $X2=0
+ $Y2=0
cc_3171 N_A_355_311#_c_4345_n N_Z_c_4693_n 0.0139315f $X=3.645 $Y=2.225 $X2=0
+ $Y2=0
cc_3172 N_A_355_311#_c_4388_n N_Z_c_4693_n 0.0236317f $X=2.985 $Y=2.225 $X2=0
+ $Y2=0
cc_3173 N_A_355_311#_c_4338_n N_Z_c_4693_n 0.0151604f $X=2.84 $Y=1.7 $X2=0 $Y2=0
cc_3174 N_A_355_311#_c_4343_n Z 0.0238869f $X=2.695 $Y=2.225 $X2=0 $Y2=0
cc_3175 N_A_355_311#_c_4337_n Z 0.00168706f $X=1.9 $Y=1.73 $X2=0 $Y2=0
cc_3176 N_A_355_311#_c_4338_n Z 6.68271e-19 $X=2.84 $Y=1.7 $X2=0 $Y2=0
cc_3177 N_A_355_311#_c_4343_n N_Z_c_4650_n 0.0181912f $X=2.695 $Y=2.225 $X2=0
+ $Y2=0
cc_3178 N_A_355_311#_c_4385_n N_Z_c_4650_n 0.0025679f $X=2.035 $Y=2.225 $X2=0
+ $Y2=0
cc_3179 N_A_355_311#_c_4388_n N_Z_c_4650_n 0.00259673f $X=2.985 $Y=2.225 $X2=0
+ $Y2=0
cc_3180 N_A_355_311#_c_4337_n N_Z_c_4650_n 0.0402246f $X=1.9 $Y=1.73 $X2=0 $Y2=0
cc_3181 N_A_355_311#_c_4338_n N_Z_c_4650_n 0.0438531f $X=2.84 $Y=1.7 $X2=0 $Y2=0
cc_3182 N_A_355_311#_c_4335_n N_Z_c_4651_n 0.00915958f $X=3.945 $Y=1.58 $X2=0
+ $Y2=0
cc_3183 N_A_355_311#_c_4345_n N_Z_c_4651_n 0.0174871f $X=3.645 $Y=2.225 $X2=0
+ $Y2=0
cc_3184 N_A_355_311#_c_4388_n N_Z_c_4651_n 0.00259673f $X=2.985 $Y=2.225 $X2=0
+ $Y2=0
cc_3185 N_A_355_311#_c_4393_n N_Z_c_4651_n 0.0025679f $X=3.935 $Y=2.225 $X2=0
+ $Y2=0
cc_3186 N_A_355_311#_c_4338_n N_Z_c_4651_n 0.0438531f $X=2.84 $Y=1.7 $X2=0 $Y2=0
cc_3187 N_A_355_311#_c_4339_n N_Z_c_4651_n 0.0383005f $X=3.78 $Y=1.7 $X2=0 $Y2=0
cc_3188 N_A_355_311#_c_4334_n N_A_405_66#_c_6931_n 0.0147893f $X=4.605 $Y=1.58
+ $X2=0 $Y2=0
cc_3189 N_A_355_311#_c_4334_n N_A_405_66#_c_6932_n 0.00239279f $X=4.605 $Y=1.58
+ $X2=0 $Y2=0
cc_3190 N_A_355_311#_c_4335_n N_A_405_66#_c_6932_n 0.00761509f $X=3.945 $Y=1.58
+ $X2=0 $Y2=0
cc_3191 N_A_355_311#_c_4360_n N_A_405_66#_c_6934_n 6.95815e-19 $X=4.77 $Y=1.66
+ $X2=0 $Y2=0
cc_3192 N_A_355_613#_c_4465_n N_Z_c_4591_n 0.0192125f $X=2.84 $Y=3.21 $X2=0
+ $Y2=0
cc_3193 N_A_355_613#_c_4465_n N_Z_c_4609_n 0.0024794f $X=2.84 $Y=3.21 $X2=0
+ $Y2=0
cc_3194 N_A_355_613#_M1123_d N_Z_c_4645_n 2.15519e-19 $X=3.635 $Y=3.065 $X2=0
+ $Y2=0
cc_3195 N_A_355_613#_c_4461_n N_Z_c_4645_n 0.0242319f $X=4.605 $Y=3.86 $X2=0
+ $Y2=0
cc_3196 N_A_355_613#_c_4483_n N_Z_c_4645_n 0.020688f $X=5.545 $Y=3.86 $X2=0
+ $Y2=0
cc_3197 N_A_355_613#_c_4472_n N_Z_c_4645_n 0.0146113f $X=3.645 $Y=3.215 $X2=0
+ $Y2=0
cc_3198 N_A_355_613#_c_4463_n N_Z_c_4645_n 0.0521734f $X=4.625 $Y=3.215 $X2=0
+ $Y2=0
cc_3199 N_A_355_613#_c_4520_n N_Z_c_4645_n 0.0238046f $X=3.935 $Y=3.215 $X2=0
+ $Y2=0
cc_3200 N_A_355_613#_c_4496_n N_Z_c_4645_n 0.0481433f $X=5.565 $Y=3.215 $X2=0
+ $Y2=0
cc_3201 N_A_355_613#_c_4526_n N_Z_c_4645_n 0.0238869f $X=4.915 $Y=3.215 $X2=0
+ $Y2=0
cc_3202 N_A_355_613#_c_4529_n N_Z_c_4645_n 0.0238869f $X=5.71 $Y=3.215 $X2=0
+ $Y2=0
cc_3203 N_A_355_613#_c_4466_n N_Z_c_4645_n 0.026602f $X=3.78 $Y=3.21 $X2=0 $Y2=0
cc_3204 N_A_355_613#_c_4499_n N_Z_c_4645_n 0.0205035f $X=4.77 $Y=3.1 $X2=0 $Y2=0
cc_3205 N_A_355_613#_c_4502_n N_Z_c_4645_n 0.0187608f $X=5.71 $Y=3.1 $X2=0 $Y2=0
cc_3206 N_A_355_613#_c_4472_n N_Z_c_5164_n 0.0238869f $X=3.645 $Y=3.215 $X2=0
+ $Y2=0
cc_3207 N_A_355_613#_c_4465_n N_Z_c_5164_n 6.68271e-19 $X=2.84 $Y=3.21 $X2=0
+ $Y2=0
cc_3208 N_A_355_613#_c_4466_n N_Z_c_5164_n 6.74054e-19 $X=3.78 $Y=3.21 $X2=0
+ $Y2=0
cc_3209 N_A_355_613#_M1080_d N_Z_c_4718_n 3.28377e-19 $X=2.695 $Y=3.065 $X2=0
+ $Y2=0
cc_3210 N_A_355_613#_c_4470_n N_Z_c_4718_n 0.0139315f $X=2.695 $Y=3.215 $X2=0
+ $Y2=0
cc_3211 N_A_355_613#_c_4472_n N_Z_c_4718_n 0.0139315f $X=3.645 $Y=3.215 $X2=0
+ $Y2=0
cc_3212 N_A_355_613#_c_4515_n N_Z_c_4718_n 0.0236317f $X=2.985 $Y=3.215 $X2=0
+ $Y2=0
cc_3213 N_A_355_613#_c_4465_n N_Z_c_4718_n 0.0151604f $X=2.84 $Y=3.21 $X2=0
+ $Y2=0
cc_3214 N_A_355_613#_c_4470_n Z 0.0238869f $X=2.695 $Y=3.215 $X2=0 $Y2=0
cc_3215 N_A_355_613#_c_4464_n Z 0.00168706f $X=1.9 $Y=3.21 $X2=0 $Y2=0
cc_3216 N_A_355_613#_c_4465_n Z 6.68271e-19 $X=2.84 $Y=3.21 $X2=0 $Y2=0
cc_3217 N_A_355_613#_c_4470_n N_Z_c_4650_n 0.0181912f $X=2.695 $Y=3.215 $X2=0
+ $Y2=0
cc_3218 N_A_355_613#_c_4512_n N_Z_c_4650_n 0.0025679f $X=2.035 $Y=3.215 $X2=0
+ $Y2=0
cc_3219 N_A_355_613#_c_4515_n N_Z_c_4650_n 0.00259673f $X=2.985 $Y=3.215 $X2=0
+ $Y2=0
cc_3220 N_A_355_613#_c_4464_n N_Z_c_4650_n 0.0402246f $X=1.9 $Y=3.21 $X2=0 $Y2=0
cc_3221 N_A_355_613#_c_4465_n N_Z_c_4650_n 0.0438531f $X=2.84 $Y=3.21 $X2=0
+ $Y2=0
cc_3222 N_A_355_613#_c_4462_n N_Z_c_4651_n 0.00915958f $X=3.945 $Y=3.86 $X2=0
+ $Y2=0
cc_3223 N_A_355_613#_c_4472_n N_Z_c_4651_n 0.0174871f $X=3.645 $Y=3.215 $X2=0
+ $Y2=0
cc_3224 N_A_355_613#_c_4515_n N_Z_c_4651_n 0.00259673f $X=2.985 $Y=3.215 $X2=0
+ $Y2=0
cc_3225 N_A_355_613#_c_4520_n N_Z_c_4651_n 0.0025679f $X=3.935 $Y=3.215 $X2=0
+ $Y2=0
cc_3226 N_A_355_613#_c_4465_n N_Z_c_4651_n 0.0438531f $X=2.84 $Y=3.21 $X2=0
+ $Y2=0
cc_3227 N_A_355_613#_c_4466_n N_Z_c_4651_n 0.0383005f $X=3.78 $Y=3.21 $X2=0
+ $Y2=0
cc_3228 N_A_355_613#_c_4461_n N_A_405_918#_c_7015_n 0.0147893f $X=4.605 $Y=3.86
+ $X2=0 $Y2=0
cc_3229 N_A_355_613#_c_4461_n N_A_405_918#_c_7016_n 0.00239279f $X=4.605 $Y=3.86
+ $X2=0 $Y2=0
cc_3230 N_A_355_613#_c_4462_n N_A_405_918#_c_7016_n 0.00761509f $X=3.945 $Y=3.86
+ $X2=0 $Y2=0
cc_3231 N_A_355_613#_c_4487_n N_A_405_918#_c_7017_n 6.95815e-19 $X=4.77 $Y=3.78
+ $X2=0 $Y2=0
cc_3232 N_Z_c_4644_n N_A_1313_297#_M1050_s 2.15519e-19 $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3233 Z N_A_1313_297#_M1073_s 3.28377e-19 $X=9.905 $Y=1.785 $X2=0 $Y2=0
cc_3234 N_Z_c_4646_n N_A_1313_297#_M1126_s 2.15519e-19 $X=14.645 $Y=1.87 $X2=0
+ $Y2=0
cc_3235 N_Z_c_4644_n N_A_1313_297#_c_5507_n 0.020688f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3236 N_Z_c_4644_n N_A_1313_297#_c_5502_n 0.0242319f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3237 N_Z_c_4652_n N_A_1313_297#_c_5502_n 0.00915958f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3238 N_Z_c_4644_n N_A_1313_297#_c_5520_n 0.0481433f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3239 N_Z_c_4644_n N_A_1313_297#_c_5555_n 0.0238869f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3240 N_Z_c_4644_n N_A_1313_297#_c_5503_n 0.0521734f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3241 N_Z_c_4644_n N_A_1313_297#_c_5562_n 0.0238869f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3242 N_Z_c_4644_n N_A_1313_297#_c_5531_n 0.0146113f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3243 N_Z_c_5197_p N_A_1313_297#_c_5531_n 0.0238869f $X=9.255 $Y=1.87 $X2=0
+ $Y2=0
cc_3244 Z N_A_1313_297#_c_5531_n 0.0139315f $X=9.905 $Y=1.785 $X2=0 $Y2=0
cc_3245 N_Z_c_4652_n N_A_1313_297#_c_5531_n 0.0174871f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3246 N_Z_c_4644_n N_A_1313_297#_c_5566_n 0.0238046f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3247 N_Z_c_4652_n N_A_1313_297#_c_5566_n 0.0025679f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3248 N_Z_c_4646_n N_A_1313_297#_c_5533_n 0.0146113f $X=14.645 $Y=1.87 $X2=0
+ $Y2=0
cc_3249 N_Z_c_5203_p N_A_1313_297#_c_5533_n 0.0238869f $X=10.195 $Y=1.87 $X2=0
+ $Y2=0
cc_3250 Z N_A_1313_297#_c_5533_n 0.0139315f $X=9.905 $Y=1.785 $X2=0 $Y2=0
cc_3251 N_Z_c_4653_n N_A_1313_297#_c_5533_n 0.0174871f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3252 Z N_A_1313_297#_c_5569_n 0.0236317f $X=9.905 $Y=1.785 $X2=0 $Y2=0
cc_3253 N_Z_c_4652_n N_A_1313_297#_c_5569_n 0.00259673f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3254 N_Z_c_4653_n N_A_1313_297#_c_5569_n 0.00259673f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3255 N_Z_c_4644_n N_A_1313_297#_c_5523_n 0.0187608f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3256 N_Z_c_4644_n N_A_1313_297#_c_5526_n 0.0205035f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3257 N_Z_c_4646_n N_A_1313_297#_c_5578_n 0.0238046f $X=14.645 $Y=1.87 $X2=0
+ $Y2=0
cc_3258 N_Z_c_4653_n N_A_1313_297#_c_5578_n 0.0025679f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3259 N_Z_c_4644_n N_A_1313_297#_c_5504_n 0.026602f $X=8.965 $Y=1.87 $X2=0
+ $Y2=0
cc_3260 N_Z_c_5197_p N_A_1313_297#_c_5504_n 6.74054e-19 $X=9.255 $Y=1.87 $X2=0
+ $Y2=0
cc_3261 N_Z_c_4652_n N_A_1313_297#_c_5504_n 0.0383005f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3262 N_Z_c_4594_n N_A_1313_297#_c_5505_n 0.0192125f $X=9.685 $Y=1.215 $X2=0
+ $Y2=0
cc_3263 N_Z_c_4620_n N_A_1313_297#_c_5505_n 0.0024794f $X=9.95 $Y=1.215 $X2=0
+ $Y2=0
cc_3264 N_Z_c_5203_p N_A_1313_297#_c_5505_n 6.68271e-19 $X=10.195 $Y=1.87 $X2=0
+ $Y2=0
cc_3265 N_Z_c_5197_p N_A_1313_297#_c_5505_n 6.68271e-19 $X=9.255 $Y=1.87 $X2=0
+ $Y2=0
cc_3266 Z N_A_1313_297#_c_5505_n 0.0151604f $X=9.905 $Y=1.785 $X2=0 $Y2=0
cc_3267 N_Z_c_4652_n N_A_1313_297#_c_5505_n 0.0438531f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3268 N_Z_c_4653_n N_A_1313_297#_c_5505_n 0.0438531f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3269 N_Z_c_4646_n N_A_1313_297#_c_5506_n 0.0169532f $X=14.645 $Y=1.87 $X2=0
+ $Y2=0
cc_3270 N_Z_c_5203_p N_A_1313_297#_c_5506_n 6.74054e-19 $X=10.195 $Y=1.87 $X2=0
+ $Y2=0
cc_3271 N_Z_c_4653_n N_A_1313_297#_c_5506_n 0.0420527f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3272 N_Z_c_4645_n N_A_1313_591#_M1031_s 2.15519e-19 $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3273 Z N_A_1313_591#_M1036_s 3.28377e-19 $X=9.905 $Y=3.485 $X2=0 $Y2=0
cc_3274 N_Z_c_4647_n N_A_1313_591#_M1152_s 2.15519e-19 $X=14.645 $Y=3.57 $X2=0
+ $Y2=0
cc_3275 N_Z_c_4645_n N_A_1313_591#_c_5635_n 0.020688f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3276 N_Z_c_4645_n N_A_1313_591#_c_5630_n 0.0242319f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3277 N_Z_c_4652_n N_A_1313_591#_c_5630_n 0.00915958f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3278 N_Z_c_4645_n N_A_1313_591#_c_5648_n 0.0481433f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3279 N_Z_c_4645_n N_A_1313_591#_c_5683_n 0.0238869f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3280 N_Z_c_4645_n N_A_1313_591#_c_5631_n 0.0521734f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3281 N_Z_c_4645_n N_A_1313_591#_c_5690_n 0.0238869f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3282 N_Z_c_4645_n N_A_1313_591#_c_5659_n 0.0146113f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3283 N_Z_c_5237_p N_A_1313_591#_c_5659_n 0.0238869f $X=9.255 $Y=3.57 $X2=0
+ $Y2=0
cc_3284 Z N_A_1313_591#_c_5659_n 0.0139315f $X=9.905 $Y=3.485 $X2=0 $Y2=0
cc_3285 N_Z_c_4652_n N_A_1313_591#_c_5659_n 0.0174871f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3286 N_Z_c_4645_n N_A_1313_591#_c_5694_n 0.0238046f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3287 N_Z_c_4652_n N_A_1313_591#_c_5694_n 0.0025679f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3288 N_Z_c_4647_n N_A_1313_591#_c_5661_n 0.0146113f $X=14.645 $Y=3.57 $X2=0
+ $Y2=0
cc_3289 N_Z_c_5243_p N_A_1313_591#_c_5661_n 0.0238869f $X=10.195 $Y=3.57 $X2=0
+ $Y2=0
cc_3290 Z N_A_1313_591#_c_5661_n 0.0139315f $X=9.905 $Y=3.485 $X2=0 $Y2=0
cc_3291 N_Z_c_4653_n N_A_1313_591#_c_5661_n 0.0174871f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3292 Z N_A_1313_591#_c_5697_n 0.0236317f $X=9.905 $Y=3.485 $X2=0 $Y2=0
cc_3293 N_Z_c_4652_n N_A_1313_591#_c_5697_n 0.00259673f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3294 N_Z_c_4653_n N_A_1313_591#_c_5697_n 0.00259673f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3295 N_Z_c_4647_n N_A_1313_591#_c_5698_n 0.0238046f $X=14.645 $Y=3.57 $X2=0
+ $Y2=0
cc_3296 N_Z_c_4653_n N_A_1313_591#_c_5698_n 0.0025679f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3297 N_Z_c_4645_n N_A_1313_591#_c_5651_n 0.0187608f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3298 N_Z_c_4645_n N_A_1313_591#_c_5654_n 0.0205035f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3299 N_Z_c_4645_n N_A_1313_591#_c_5632_n 0.026602f $X=8.965 $Y=3.57 $X2=0
+ $Y2=0
cc_3300 N_Z_c_5237_p N_A_1313_591#_c_5632_n 6.74054e-19 $X=9.255 $Y=3.57 $X2=0
+ $Y2=0
cc_3301 N_Z_c_4652_n N_A_1313_591#_c_5632_n 0.0383005f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3302 N_Z_c_4595_n N_A_1313_591#_c_5633_n 0.0192125f $X=9.685 $Y=4.225 $X2=0
+ $Y2=0
cc_3303 N_Z_c_4621_n N_A_1313_591#_c_5633_n 0.0024794f $X=9.95 $Y=4.225 $X2=0
+ $Y2=0
cc_3304 N_Z_c_5243_p N_A_1313_591#_c_5633_n 6.68271e-19 $X=10.195 $Y=3.57 $X2=0
+ $Y2=0
cc_3305 N_Z_c_5237_p N_A_1313_591#_c_5633_n 6.68271e-19 $X=9.255 $Y=3.57 $X2=0
+ $Y2=0
cc_3306 Z N_A_1313_591#_c_5633_n 0.0151604f $X=9.905 $Y=3.485 $X2=0 $Y2=0
cc_3307 N_Z_c_4652_n N_A_1313_591#_c_5633_n 0.0438531f $X=9.11 $Y=1.7 $X2=0
+ $Y2=0
cc_3308 N_Z_c_4653_n N_A_1313_591#_c_5633_n 0.0438531f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3309 N_Z_c_4647_n N_A_1313_591#_c_5634_n 0.0169532f $X=14.645 $Y=3.57 $X2=0
+ $Y2=0
cc_3310 N_Z_c_5243_p N_A_1313_591#_c_5634_n 6.74054e-19 $X=10.195 $Y=3.57 $X2=0
+ $Y2=0
cc_3311 N_Z_c_4653_n N_A_1313_591#_c_5634_n 0.0420527f $X=10.05 $Y=1.7 $X2=0
+ $Y2=0
cc_3312 N_Z_c_4646_n N_A_2839_311#_M1004_s 2.15519e-19 $X=14.645 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_3313 N_Z_c_4895_n N_A_2839_311#_M1110_s 3.28377e-19 $X=15.585 $Y=1.87 $X2=0
+ $Y2=0
cc_3314 N_Z_c_4648_n N_A_2839_311#_M1146_s 2.15519e-19 $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3315 N_Z_c_4648_n N_A_2839_311#_c_5758_n 0.0242319f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3316 N_Z_c_4655_n N_A_2839_311#_c_5759_n 0.00915958f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3317 N_Z_c_4648_n N_A_2839_311#_c_5780_n 0.020688f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3318 N_Z_c_4646_n N_A_2839_311#_c_5767_n 0.0146113f $X=14.645 $Y=1.87 $X2=0
+ $Y2=0
cc_3319 N_Z_c_4895_n N_A_2839_311#_c_5767_n 0.0139315f $X=15.585 $Y=1.87 $X2=0
+ $Y2=0
cc_3320 Z N_A_2839_311#_c_5767_n 0.0238869f $X=14.765 $Y=1.785 $X2=0 $Y2=0
cc_3321 N_Z_c_4654_n N_A_2839_311#_c_5767_n 0.0174871f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3322 N_Z_c_4646_n N_A_2839_311#_c_5809_n 0.0238046f $X=14.645 $Y=1.87 $X2=0
+ $Y2=0
cc_3323 N_Z_c_4654_n N_A_2839_311#_c_5809_n 0.0025679f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3324 N_Z_c_4648_n N_A_2839_311#_c_5769_n 0.0146113f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3325 N_Z_c_5279_p N_A_2839_311#_c_5769_n 0.0238869f $X=15.875 $Y=1.87 $X2=0
+ $Y2=0
cc_3326 N_Z_c_4895_n N_A_2839_311#_c_5769_n 0.0139315f $X=15.585 $Y=1.87 $X2=0
+ $Y2=0
cc_3327 N_Z_c_4655_n N_A_2839_311#_c_5769_n 0.0174871f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3328 N_Z_c_4895_n N_A_2839_311#_c_5812_n 0.0236317f $X=15.585 $Y=1.87 $X2=0
+ $Y2=0
cc_3329 N_Z_c_4654_n N_A_2839_311#_c_5812_n 0.00259673f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3330 N_Z_c_4655_n N_A_2839_311#_c_5812_n 0.00259673f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3331 N_Z_c_4648_n N_A_2839_311#_c_5760_n 0.0521734f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3332 N_Z_c_4648_n N_A_2839_311#_c_5817_n 0.0238046f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3333 N_Z_c_4655_n N_A_2839_311#_c_5817_n 0.0025679f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3334 N_Z_c_4648_n N_A_2839_311#_c_5793_n 0.0481433f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3335 N_Z_c_4648_n N_A_2839_311#_c_5823_n 0.0238869f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3336 N_Z_c_4648_n N_A_2839_311#_c_5795_n 0.0205035f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3337 N_Z_c_4648_n N_A_2839_311#_c_5830_n 0.0238869f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3338 N_Z_c_4648_n N_A_2839_311#_c_5798_n 0.0187608f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3339 N_Z_c_4646_n N_A_2839_311#_c_5761_n 0.0169532f $X=14.645 $Y=1.87 $X2=0
+ $Y2=0
cc_3340 Z N_A_2839_311#_c_5761_n 6.74054e-19 $X=14.765 $Y=1.785 $X2=0 $Y2=0
cc_3341 N_Z_c_4654_n N_A_2839_311#_c_5761_n 0.0420527f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3342 N_Z_c_4600_n N_A_2839_311#_c_5762_n 0.0192125f $X=15.565 $Y=1.215 $X2=0
+ $Y2=0
cc_3343 N_Z_c_4622_n N_A_2839_311#_c_5762_n 0.0024794f $X=14.89 $Y=1.215 $X2=0
+ $Y2=0
cc_3344 N_Z_c_5279_p N_A_2839_311#_c_5762_n 6.68271e-19 $X=15.875 $Y=1.87 $X2=0
+ $Y2=0
cc_3345 N_Z_c_4895_n N_A_2839_311#_c_5762_n 0.0151604f $X=15.585 $Y=1.87 $X2=0
+ $Y2=0
cc_3346 Z N_A_2839_311#_c_5762_n 6.68271e-19 $X=14.765 $Y=1.785 $X2=0 $Y2=0
cc_3347 N_Z_c_4654_n N_A_2839_311#_c_5762_n 0.0438531f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3348 N_Z_c_4655_n N_A_2839_311#_c_5762_n 0.0438531f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3349 N_Z_c_4648_n N_A_2839_311#_c_5763_n 0.026602f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3350 N_Z_c_5279_p N_A_2839_311#_c_5763_n 6.74054e-19 $X=15.875 $Y=1.87 $X2=0
+ $Y2=0
cc_3351 N_Z_c_4655_n N_A_2839_311#_c_5763_n 0.0383005f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3352 N_Z_c_4647_n N_A_2839_613#_M1021_d 2.15519e-19 $X=14.645 $Y=3.57
+ $X2=-0.19 $Y2=-0.24
cc_3353 N_Z_c_4924_n N_A_2839_613#_M1041_d 3.28377e-19 $X=15.585 $Y=3.57 $X2=0
+ $Y2=0
cc_3354 N_Z_c_4649_n N_A_2839_613#_M1078_d 2.15519e-19 $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3355 N_Z_c_4649_n N_A_2839_613#_c_5889_n 0.0242319f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3356 N_Z_c_4655_n N_A_2839_613#_c_5890_n 0.00915958f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3357 N_Z_c_4649_n N_A_2839_613#_c_5911_n 0.020688f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3358 N_Z_c_4647_n N_A_2839_613#_c_5898_n 0.0146113f $X=14.645 $Y=3.57 $X2=0
+ $Y2=0
cc_3359 N_Z_c_4924_n N_A_2839_613#_c_5898_n 0.0139315f $X=15.585 $Y=3.57 $X2=0
+ $Y2=0
cc_3360 Z N_A_2839_613#_c_5898_n 0.0238869f $X=14.765 $Y=3.485 $X2=0 $Y2=0
cc_3361 N_Z_c_4654_n N_A_2839_613#_c_5898_n 0.0174871f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3362 N_Z_c_4647_n N_A_2839_613#_c_5940_n 0.0238046f $X=14.645 $Y=3.57 $X2=0
+ $Y2=0
cc_3363 N_Z_c_4654_n N_A_2839_613#_c_5940_n 0.0025679f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3364 N_Z_c_4649_n N_A_2839_613#_c_5900_n 0.0146113f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3365 N_Z_c_5319_p N_A_2839_613#_c_5900_n 0.0238869f $X=15.875 $Y=3.57 $X2=0
+ $Y2=0
cc_3366 N_Z_c_4924_n N_A_2839_613#_c_5900_n 0.0139315f $X=15.585 $Y=3.57 $X2=0
+ $Y2=0
cc_3367 N_Z_c_4655_n N_A_2839_613#_c_5900_n 0.0174871f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3368 N_Z_c_4924_n N_A_2839_613#_c_5943_n 0.0236317f $X=15.585 $Y=3.57 $X2=0
+ $Y2=0
cc_3369 N_Z_c_4654_n N_A_2839_613#_c_5943_n 0.00259673f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3370 N_Z_c_4655_n N_A_2839_613#_c_5943_n 0.00259673f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3371 N_Z_c_4649_n N_A_2839_613#_c_5891_n 0.0521734f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3372 N_Z_c_4649_n N_A_2839_613#_c_5948_n 0.0238046f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3373 N_Z_c_4655_n N_A_2839_613#_c_5948_n 0.0025679f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3374 N_Z_c_4649_n N_A_2839_613#_c_5924_n 0.0481433f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3375 N_Z_c_4649_n N_A_2839_613#_c_5954_n 0.0238869f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3376 N_Z_c_4649_n N_A_2839_613#_c_5957_n 0.0238869f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3377 N_Z_c_4647_n N_A_2839_613#_c_5892_n 0.0169532f $X=14.645 $Y=3.57 $X2=0
+ $Y2=0
cc_3378 Z N_A_2839_613#_c_5892_n 6.74054e-19 $X=14.765 $Y=3.485 $X2=0 $Y2=0
cc_3379 N_Z_c_4654_n N_A_2839_613#_c_5892_n 0.0420527f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3380 N_Z_c_4601_n N_A_2839_613#_c_5893_n 0.0192125f $X=15.565 $Y=4.225 $X2=0
+ $Y2=0
cc_3381 N_Z_c_4623_n N_A_2839_613#_c_5893_n 0.0024794f $X=14.89 $Y=4.225 $X2=0
+ $Y2=0
cc_3382 N_Z_c_5319_p N_A_2839_613#_c_5893_n 6.68271e-19 $X=15.875 $Y=3.57 $X2=0
+ $Y2=0
cc_3383 N_Z_c_4924_n N_A_2839_613#_c_5893_n 0.0151604f $X=15.585 $Y=3.57 $X2=0
+ $Y2=0
cc_3384 Z N_A_2839_613#_c_5893_n 6.68271e-19 $X=14.765 $Y=3.485 $X2=0 $Y2=0
cc_3385 N_Z_c_4654_n N_A_2839_613#_c_5893_n 0.0438531f $X=14.79 $Y=1.7 $X2=0
+ $Y2=0
cc_3386 N_Z_c_4655_n N_A_2839_613#_c_5893_n 0.0438531f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3387 N_Z_c_4649_n N_A_2839_613#_c_5894_n 0.026602f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3388 N_Z_c_5319_p N_A_2839_613#_c_5894_n 6.74054e-19 $X=15.875 $Y=3.57 $X2=0
+ $Y2=0
cc_3389 N_Z_c_4655_n N_A_2839_613#_c_5894_n 0.0383005f $X=15.73 $Y=1.7 $X2=0
+ $Y2=0
cc_3390 N_Z_c_4649_n N_A_2839_613#_c_5927_n 0.0205035f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3391 N_Z_c_4649_n N_A_2839_613#_c_5930_n 0.0187608f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3392 N_Z_c_4648_n N_A_3797_297#_M1002_d 2.15519e-19 $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3393 Z N_A_3797_297#_M1023_d 3.28377e-19 $X=22.325 $Y=1.785 $X2=0 $Y2=0
cc_3394 N_Z_c_4648_n N_A_3797_297#_c_6025_n 0.020688f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3395 N_Z_c_4648_n N_A_3797_297#_c_6020_n 0.0242319f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3396 N_Z_c_4656_n N_A_3797_297#_c_6020_n 0.00915958f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3397 N_Z_c_4648_n N_A_3797_297#_c_6038_n 0.0481433f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3398 N_Z_c_4648_n N_A_3797_297#_c_6073_n 0.0238869f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3399 N_Z_c_4648_n N_A_3797_297#_c_6021_n 0.0521734f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3400 N_Z_c_4648_n N_A_3797_297#_c_6080_n 0.0238869f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3401 N_Z_c_4648_n N_A_3797_297#_c_6049_n 0.0146113f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3402 N_Z_c_5356_p N_A_3797_297#_c_6049_n 0.0238869f $X=21.675 $Y=1.87 $X2=0
+ $Y2=0
cc_3403 Z N_A_3797_297#_c_6049_n 0.0139315f $X=22.325 $Y=1.785 $X2=0 $Y2=0
cc_3404 N_Z_c_4656_n N_A_3797_297#_c_6049_n 0.0174871f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3405 N_Z_c_4648_n N_A_3797_297#_c_6084_n 0.0238046f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3406 N_Z_c_4656_n N_A_3797_297#_c_6084_n 0.0025679f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3407 Z N_A_3797_297#_c_6051_n 0.0378184f $X=22.325 $Y=1.785 $X2=0 $Y2=0
cc_3408 N_Z_c_4657_n N_A_3797_297#_c_6051_n 0.0181912f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3409 Z N_A_3797_297#_c_6087_n 0.0236317f $X=22.325 $Y=1.785 $X2=0 $Y2=0
cc_3410 N_Z_c_4656_n N_A_3797_297#_c_6087_n 0.00259673f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3411 N_Z_c_4657_n N_A_3797_297#_c_6087_n 0.00259673f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3412 N_Z_c_4648_n N_A_3797_297#_c_6041_n 0.0187608f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3413 N_Z_c_4648_n N_A_3797_297#_c_6044_n 0.0205035f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3414 N_Z_c_4657_n N_A_3797_297#_c_6096_n 0.0025679f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3415 N_Z_c_4648_n N_A_3797_297#_c_6022_n 0.026602f $X=21.385 $Y=1.87 $X2=0
+ $Y2=0
cc_3416 N_Z_c_5356_p N_A_3797_297#_c_6022_n 6.74054e-19 $X=21.675 $Y=1.87 $X2=0
+ $Y2=0
cc_3417 N_Z_c_4656_n N_A_3797_297#_c_6022_n 0.0383005f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3418 N_Z_c_4604_n N_A_3797_297#_c_6023_n 0.0192125f $X=22.105 $Y=1.215 $X2=0
+ $Y2=0
cc_3419 N_Z_c_4634_n N_A_3797_297#_c_6023_n 0.0024794f $X=22.37 $Y=1.215 $X2=0
+ $Y2=0
cc_3420 N_Z_c_5356_p N_A_3797_297#_c_6023_n 6.68271e-19 $X=21.675 $Y=1.87 $X2=0
+ $Y2=0
cc_3421 Z N_A_3797_297#_c_6023_n 0.0158287f $X=22.325 $Y=1.785 $X2=0 $Y2=0
cc_3422 N_Z_c_4656_n N_A_3797_297#_c_6023_n 0.0438531f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3423 N_Z_c_4657_n N_A_3797_297#_c_6023_n 0.0438531f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3424 Z N_A_3797_297#_c_6024_n 0.00168706f $X=22.325 $Y=1.785 $X2=0 $Y2=0
cc_3425 N_Z_c_4657_n N_A_3797_297#_c_6024_n 0.0402246f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3426 N_Z_c_4649_n N_A_3797_591#_M1011_d 2.15519e-19 $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3427 Z N_A_3797_591#_M1053_d 3.28377e-19 $X=22.325 $Y=3.485 $X2=0 $Y2=0
cc_3428 N_Z_c_4649_n N_A_3797_591#_c_6147_n 0.020688f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3429 N_Z_c_4649_n N_A_3797_591#_c_6142_n 0.0242319f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3430 N_Z_c_4656_n N_A_3797_591#_c_6142_n 0.00915958f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3431 N_Z_c_4649_n N_A_3797_591#_c_6160_n 0.0481433f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3432 N_Z_c_4649_n N_A_3797_591#_c_6195_n 0.0238869f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3433 N_Z_c_4649_n N_A_3797_591#_c_6143_n 0.0521734f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3434 N_Z_c_4649_n N_A_3797_591#_c_6202_n 0.0238869f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3435 N_Z_c_4649_n N_A_3797_591#_c_6171_n 0.0146113f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3436 N_Z_c_5390_p N_A_3797_591#_c_6171_n 0.0238869f $X=21.675 $Y=3.57 $X2=0
+ $Y2=0
cc_3437 Z N_A_3797_591#_c_6171_n 0.0139315f $X=22.325 $Y=3.485 $X2=0 $Y2=0
cc_3438 N_Z_c_4656_n N_A_3797_591#_c_6171_n 0.0174871f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3439 N_Z_c_4649_n N_A_3797_591#_c_6206_n 0.0238046f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3440 N_Z_c_4656_n N_A_3797_591#_c_6206_n 0.0025679f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3441 Z N_A_3797_591#_c_6173_n 0.0378184f $X=22.325 $Y=3.485 $X2=0 $Y2=0
cc_3442 N_Z_c_4657_n N_A_3797_591#_c_6173_n 0.0181912f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3443 Z N_A_3797_591#_c_6209_n 0.0236317f $X=22.325 $Y=3.485 $X2=0 $Y2=0
cc_3444 N_Z_c_4656_n N_A_3797_591#_c_6209_n 0.00259673f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3445 N_Z_c_4657_n N_A_3797_591#_c_6209_n 0.00259673f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3446 N_Z_c_4657_n N_A_3797_591#_c_6210_n 0.0025679f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3447 N_Z_c_4649_n N_A_3797_591#_c_6163_n 0.0187608f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3448 N_Z_c_4649_n N_A_3797_591#_c_6166_n 0.0205035f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3449 N_Z_c_4649_n N_A_3797_591#_c_6144_n 0.026602f $X=21.385 $Y=3.57 $X2=0
+ $Y2=0
cc_3450 N_Z_c_5390_p N_A_3797_591#_c_6144_n 6.74054e-19 $X=21.675 $Y=3.57 $X2=0
+ $Y2=0
cc_3451 N_Z_c_4656_n N_A_3797_591#_c_6144_n 0.0383005f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3452 N_Z_c_4605_n N_A_3797_591#_c_6145_n 0.0192125f $X=22.105 $Y=4.225 $X2=0
+ $Y2=0
cc_3453 N_Z_c_4635_n N_A_3797_591#_c_6145_n 0.0024794f $X=22.37 $Y=4.225 $X2=0
+ $Y2=0
cc_3454 N_Z_c_5390_p N_A_3797_591#_c_6145_n 6.68271e-19 $X=21.675 $Y=3.57 $X2=0
+ $Y2=0
cc_3455 Z N_A_3797_591#_c_6145_n 0.0158287f $X=22.325 $Y=3.485 $X2=0 $Y2=0
cc_3456 N_Z_c_4656_n N_A_3797_591#_c_6145_n 0.0438531f $X=21.53 $Y=1.7 $X2=0
+ $Y2=0
cc_3457 N_Z_c_4657_n N_A_3797_591#_c_6145_n 0.0438531f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3458 Z N_A_3797_591#_c_6146_n 0.00168706f $X=22.325 $Y=3.485 $X2=0 $Y2=0
cc_3459 N_Z_c_4657_n N_A_3797_591#_c_6146_n 0.0402246f $X=22.47 $Y=1.7 $X2=0
+ $Y2=0
cc_3460 N_Z_c_4608_n N_A_405_66#_c_6926_n 0.00158445f $X=2.47 $Y=1.215 $X2=0
+ $Y2=0
cc_3461 N_Z_M1003_s N_A_405_66#_c_6927_n 0.00165831f $X=2.435 $Y=0.33 $X2=0
+ $Y2=0
cc_3462 N_Z_c_4588_n N_A_405_66#_c_6927_n 0.015949f $X=2.57 $Y=0.68 $X2=0 $Y2=0
cc_3463 N_Z_c_4590_n N_A_405_66#_c_6927_n 0.00405549f $X=3.145 $Y=1.215 $X2=0
+ $Y2=0
cc_3464 N_Z_c_4608_n N_A_405_66#_c_6927_n 0.00443806f $X=2.47 $Y=1.215 $X2=0
+ $Y2=0
cc_3465 N_Z_c_4590_n N_A_405_66#_c_6948_n 0.00918654f $X=3.145 $Y=1.215 $X2=0
+ $Y2=0
cc_3466 N_Z_M1109_s N_A_405_66#_c_6929_n 0.00165831f $X=3.275 $Y=0.33 $X2=0
+ $Y2=0
cc_3467 N_Z_c_4590_n N_A_405_66#_c_6929_n 0.00133192f $X=3.145 $Y=1.215 $X2=0
+ $Y2=0
cc_3468 N_Z_c_4610_n N_A_405_66#_c_6929_n 0.00293855f $X=3.31 $Y=1.215 $X2=0
+ $Y2=0
cc_3469 N_Z_c_4612_n N_A_405_66#_c_6929_n 0.0157607f $X=3.41 $Y=0.68 $X2=0 $Y2=0
cc_3470 N_Z_c_4612_n N_A_405_66#_c_6932_n 0.00799417f $X=3.41 $Y=0.68 $X2=0
+ $Y2=0
cc_3471 N_Z_c_4609_n N_A_405_918#_c_7010_n 0.00158445f $X=2.47 $Y=4.225 $X2=0
+ $Y2=0
cc_3472 N_Z_M1029_s N_A_405_918#_c_7011_n 0.00165831f $X=2.435 $Y=4.59 $X2=0
+ $Y2=0
cc_3473 N_Z_c_4589_n N_A_405_918#_c_7011_n 0.015949f $X=2.57 $Y=4.76 $X2=0 $Y2=0
cc_3474 N_Z_c_4591_n N_A_405_918#_c_7011_n 0.00405549f $X=3.145 $Y=4.225 $X2=0
+ $Y2=0
cc_3475 N_Z_c_4609_n N_A_405_918#_c_7011_n 0.00443806f $X=2.47 $Y=4.225 $X2=0
+ $Y2=0
cc_3476 N_Z_c_4591_n N_A_405_918#_c_7032_n 0.00918654f $X=3.145 $Y=4.225 $X2=0
+ $Y2=0
cc_3477 N_Z_M1083_s N_A_405_918#_c_7013_n 0.00165831f $X=3.275 $Y=4.59 $X2=0
+ $Y2=0
cc_3478 N_Z_c_4591_n N_A_405_918#_c_7013_n 0.00133192f $X=3.145 $Y=4.225 $X2=0
+ $Y2=0
cc_3479 N_Z_c_4611_n N_A_405_918#_c_7013_n 0.00293855f $X=3.31 $Y=4.225 $X2=0
+ $Y2=0
cc_3480 N_Z_c_4613_n N_A_405_918#_c_7013_n 0.0157607f $X=3.41 $Y=4.76 $X2=0
+ $Y2=0
cc_3481 N_Z_c_4613_n N_A_405_918#_c_7016_n 0.00799417f $X=3.41 $Y=4.76 $X2=0
+ $Y2=0
cc_3482 N_Z_c_4615_n N_A_1315_47#_c_7093_n 0.00799417f $X=9.01 $Y=0.68 $X2=0
+ $Y2=0
cc_3483 N_Z_M1024_d N_A_1315_47#_c_7095_n 0.00165831f $X=8.875 $Y=0.33 $X2=0
+ $Y2=0
cc_3484 N_Z_c_4594_n N_A_1315_47#_c_7095_n 0.00133192f $X=9.685 $Y=1.215 $X2=0
+ $Y2=0
cc_3485 N_Z_c_4615_n N_A_1315_47#_c_7095_n 0.0157607f $X=9.01 $Y=0.68 $X2=0
+ $Y2=0
cc_3486 N_Z_c_4618_n N_A_1315_47#_c_7095_n 0.00293855f $X=9.11 $Y=1.215 $X2=0
+ $Y2=0
cc_3487 N_Z_c_4594_n N_A_1315_47#_c_7120_n 0.00918654f $X=9.685 $Y=1.215 $X2=0
+ $Y2=0
cc_3488 N_Z_M1044_d N_A_1315_47#_c_7097_n 0.00165831f $X=9.715 $Y=0.33 $X2=0
+ $Y2=0
cc_3489 N_Z_c_4594_n N_A_1315_47#_c_7097_n 0.00405549f $X=9.685 $Y=1.215 $X2=0
+ $Y2=0
cc_3490 N_Z_c_4596_n N_A_1315_47#_c_7097_n 0.015949f $X=9.85 $Y=0.68 $X2=0 $Y2=0
cc_3491 N_Z_c_4620_n N_A_1315_47#_c_7097_n 0.00443806f $X=9.95 $Y=1.215 $X2=0
+ $Y2=0
cc_3492 N_Z_c_4620_n N_A_1315_47#_c_7098_n 0.00158445f $X=9.95 $Y=1.215 $X2=0
+ $Y2=0
cc_3493 N_Z_c_4616_n N_A_1315_911#_c_7175_n 0.00799417f $X=9.01 $Y=4.76 $X2=0
+ $Y2=0
cc_3494 N_Z_M1016_d N_A_1315_911#_c_7177_n 0.00165831f $X=8.875 $Y=4.59 $X2=0
+ $Y2=0
cc_3495 N_Z_c_4595_n N_A_1315_911#_c_7177_n 0.00133192f $X=9.685 $Y=4.225 $X2=0
+ $Y2=0
cc_3496 N_Z_c_4616_n N_A_1315_911#_c_7177_n 0.0157607f $X=9.01 $Y=4.76 $X2=0
+ $Y2=0
cc_3497 N_Z_c_4619_n N_A_1315_911#_c_7177_n 0.00293855f $X=9.11 $Y=4.225 $X2=0
+ $Y2=0
cc_3498 N_Z_c_4595_n N_A_1315_911#_c_7199_n 0.00918654f $X=9.685 $Y=4.225 $X2=0
+ $Y2=0
cc_3499 N_Z_M1048_d N_A_1315_911#_c_7179_n 0.00165831f $X=9.715 $Y=4.59 $X2=0
+ $Y2=0
cc_3500 N_Z_c_4595_n N_A_1315_911#_c_7179_n 0.00405549f $X=9.685 $Y=4.225 $X2=0
+ $Y2=0
cc_3501 N_Z_c_4597_n N_A_1315_911#_c_7179_n 0.015949f $X=9.85 $Y=4.76 $X2=0
+ $Y2=0
cc_3502 N_Z_c_4621_n N_A_1315_911#_c_7179_n 0.00443806f $X=9.95 $Y=4.225 $X2=0
+ $Y2=0
cc_3503 N_Z_c_4621_n N_A_1315_911#_c_7180_n 0.00158445f $X=9.95 $Y=4.225 $X2=0
+ $Y2=0
cc_3504 N_Z_c_4622_n N_A_2889_66#_c_7254_n 0.00158445f $X=14.89 $Y=1.215 $X2=0
+ $Y2=0
cc_3505 N_Z_M1006_s N_A_2889_66#_c_7255_n 0.00165831f $X=14.855 $Y=0.33 $X2=0
+ $Y2=0
cc_3506 N_Z_c_4598_n N_A_2889_66#_c_7255_n 0.015949f $X=14.99 $Y=0.68 $X2=0
+ $Y2=0
cc_3507 N_Z_c_4600_n N_A_2889_66#_c_7255_n 0.00405549f $X=15.565 $Y=1.215 $X2=0
+ $Y2=0
cc_3508 N_Z_c_4622_n N_A_2889_66#_c_7255_n 0.00443806f $X=14.89 $Y=1.215 $X2=0
+ $Y2=0
cc_3509 N_Z_c_4600_n N_A_2889_66#_c_7276_n 0.00918654f $X=15.565 $Y=1.215 $X2=0
+ $Y2=0
cc_3510 N_Z_M1035_s N_A_2889_66#_c_7257_n 0.00165831f $X=15.695 $Y=0.33 $X2=0
+ $Y2=0
cc_3511 N_Z_c_4600_n N_A_2889_66#_c_7257_n 0.00133192f $X=15.565 $Y=1.215 $X2=0
+ $Y2=0
cc_3512 N_Z_c_4624_n N_A_2889_66#_c_7257_n 0.00293855f $X=15.73 $Y=1.215 $X2=0
+ $Y2=0
cc_3513 N_Z_c_4626_n N_A_2889_66#_c_7257_n 0.0157607f $X=15.83 $Y=0.68 $X2=0
+ $Y2=0
cc_3514 N_Z_c_4626_n N_A_2889_66#_c_7260_n 0.00799417f $X=15.83 $Y=0.68 $X2=0
+ $Y2=0
cc_3515 N_Z_c_4623_n N_A_2889_918#_c_7338_n 0.00158445f $X=14.89 $Y=4.225 $X2=0
+ $Y2=0
cc_3516 N_Z_M1009_d N_A_2889_918#_c_7339_n 0.00165831f $X=14.855 $Y=4.59 $X2=0
+ $Y2=0
cc_3517 N_Z_c_4599_n N_A_2889_918#_c_7339_n 0.015949f $X=14.99 $Y=4.76 $X2=0
+ $Y2=0
cc_3518 N_Z_c_4601_n N_A_2889_918#_c_7339_n 0.00405549f $X=15.565 $Y=4.225 $X2=0
+ $Y2=0
cc_3519 N_Z_c_4623_n N_A_2889_918#_c_7339_n 0.00443806f $X=14.89 $Y=4.225 $X2=0
+ $Y2=0
cc_3520 N_Z_c_4601_n N_A_2889_918#_c_7360_n 0.00918654f $X=15.565 $Y=4.225 $X2=0
+ $Y2=0
cc_3521 N_Z_M1112_d N_A_2889_918#_c_7341_n 0.00165831f $X=15.695 $Y=4.59 $X2=0
+ $Y2=0
cc_3522 N_Z_c_4601_n N_A_2889_918#_c_7341_n 0.00133192f $X=15.565 $Y=4.225 $X2=0
+ $Y2=0
cc_3523 N_Z_c_4625_n N_A_2889_918#_c_7341_n 0.00293855f $X=15.73 $Y=4.225 $X2=0
+ $Y2=0
cc_3524 N_Z_c_4627_n N_A_2889_918#_c_7341_n 0.0157607f $X=15.83 $Y=4.76 $X2=0
+ $Y2=0
cc_3525 N_Z_c_4627_n N_A_2889_918#_c_7344_n 0.00799417f $X=15.83 $Y=4.76 $X2=0
+ $Y2=0
cc_3526 N_Z_c_4629_n N_A_3799_47#_c_7421_n 0.00799417f $X=21.43 $Y=0.68 $X2=0
+ $Y2=0
cc_3527 N_Z_M1089_s N_A_3799_47#_c_7423_n 0.00165831f $X=21.295 $Y=0.33 $X2=0
+ $Y2=0
cc_3528 N_Z_c_4604_n N_A_3799_47#_c_7423_n 0.00133192f $X=22.105 $Y=1.215 $X2=0
+ $Y2=0
cc_3529 N_Z_c_4629_n N_A_3799_47#_c_7423_n 0.0157607f $X=21.43 $Y=0.68 $X2=0
+ $Y2=0
cc_3530 N_Z_c_4632_n N_A_3799_47#_c_7423_n 0.00293855f $X=21.53 $Y=1.215 $X2=0
+ $Y2=0
cc_3531 N_Z_c_4604_n N_A_3799_47#_c_7448_n 0.00918654f $X=22.105 $Y=1.215 $X2=0
+ $Y2=0
cc_3532 N_Z_M1122_s N_A_3799_47#_c_7425_n 0.00165831f $X=22.135 $Y=0.33 $X2=0
+ $Y2=0
cc_3533 N_Z_c_4604_n N_A_3799_47#_c_7425_n 0.00405549f $X=22.105 $Y=1.215 $X2=0
+ $Y2=0
cc_3534 N_Z_c_4606_n N_A_3799_47#_c_7425_n 0.015949f $X=22.27 $Y=0.68 $X2=0
+ $Y2=0
cc_3535 N_Z_c_4634_n N_A_3799_47#_c_7425_n 0.00443806f $X=22.37 $Y=1.215 $X2=0
+ $Y2=0
cc_3536 N_Z_c_4634_n N_A_3799_47#_c_7426_n 0.00158445f $X=22.37 $Y=1.215 $X2=0
+ $Y2=0
cc_3537 N_Z_c_4630_n N_A_3799_911#_c_7503_n 0.00799417f $X=21.43 $Y=4.76 $X2=0
+ $Y2=0
cc_3538 N_Z_M1008_d N_A_3799_911#_c_7505_n 0.00165831f $X=21.295 $Y=4.59 $X2=0
+ $Y2=0
cc_3539 N_Z_c_4605_n N_A_3799_911#_c_7505_n 0.00133192f $X=22.105 $Y=4.225 $X2=0
+ $Y2=0
cc_3540 N_Z_c_4630_n N_A_3799_911#_c_7505_n 0.0157607f $X=21.43 $Y=4.76 $X2=0
+ $Y2=0
cc_3541 N_Z_c_4633_n N_A_3799_911#_c_7505_n 0.00293855f $X=21.53 $Y=4.225 $X2=0
+ $Y2=0
cc_3542 N_Z_c_4605_n N_A_3799_911#_c_7527_n 0.00918654f $X=22.105 $Y=4.225 $X2=0
+ $Y2=0
cc_3543 N_Z_M1091_d N_A_3799_911#_c_7507_n 0.00165831f $X=22.135 $Y=4.59 $X2=0
+ $Y2=0
cc_3544 N_Z_c_4605_n N_A_3799_911#_c_7507_n 0.00405549f $X=22.105 $Y=4.225 $X2=0
+ $Y2=0
cc_3545 N_Z_c_4607_n N_A_3799_911#_c_7507_n 0.015949f $X=22.27 $Y=4.76 $X2=0
+ $Y2=0
cc_3546 N_Z_c_4635_n N_A_3799_911#_c_7507_n 0.00443806f $X=22.37 $Y=4.225 $X2=0
+ $Y2=0
cc_3547 N_Z_c_4635_n N_A_3799_911#_c_7508_n 0.00158445f $X=22.37 $Y=4.225 $X2=0
+ $Y2=0
cc_3548 N_A_1313_297#_c_5505_n N_A_1313_591#_c_5633_n 0.00460759f $X=9.58 $Y=1.7
+ $X2=0 $Y2=0
cc_3549 N_A_1313_297#_c_5502_n N_A_1315_47#_c_7093_n 0.0247972f $X=8.475 $Y=1.58
+ $X2=0 $Y2=0
cc_3550 N_A_1313_297#_c_5516_n N_A_1315_47#_c_7099_n 6.95815e-19 $X=7.65 $Y=1.66
+ $X2=0 $Y2=0
cc_3551 N_A_1313_591#_c_5630_n N_A_1315_911#_c_7175_n 0.0247972f $X=8.475
+ $Y=3.86 $X2=0 $Y2=0
cc_3552 N_A_1313_591#_c_5644_n N_A_1315_911#_c_7182_n 6.95815e-19 $X=7.65
+ $Y=3.78 $X2=0 $Y2=0
cc_3553 N_A_2839_311#_c_5762_n N_A_2839_613#_c_5893_n 0.00460759f $X=15.26
+ $Y=1.7 $X2=0 $Y2=0
cc_3554 N_A_2839_311#_c_5758_n N_A_2889_66#_c_7259_n 0.0147893f $X=17.025
+ $Y=1.58 $X2=0 $Y2=0
cc_3555 N_A_2839_311#_c_5758_n N_A_2889_66#_c_7260_n 0.00239279f $X=17.025
+ $Y=1.58 $X2=0 $Y2=0
cc_3556 N_A_2839_311#_c_5759_n N_A_2889_66#_c_7260_n 0.00761509f $X=16.365
+ $Y=1.58 $X2=0 $Y2=0
cc_3557 N_A_2839_311#_c_5784_n N_A_2889_66#_c_7262_n 6.95815e-19 $X=17.19
+ $Y=1.66 $X2=0 $Y2=0
cc_3558 N_A_2839_613#_c_5889_n N_A_2889_918#_c_7343_n 0.0147893f $X=17.025
+ $Y=3.86 $X2=0 $Y2=0
cc_3559 N_A_2839_613#_c_5889_n N_A_2889_918#_c_7344_n 0.00239279f $X=17.025
+ $Y=3.86 $X2=0 $Y2=0
cc_3560 N_A_2839_613#_c_5890_n N_A_2889_918#_c_7344_n 0.00761509f $X=16.365
+ $Y=3.86 $X2=0 $Y2=0
cc_3561 N_A_2839_613#_c_5915_n N_A_2889_918#_c_7345_n 6.95815e-19 $X=17.19
+ $Y=3.78 $X2=0 $Y2=0
cc_3562 N_A_3797_297#_c_6023_n N_A_3797_591#_c_6145_n 0.00460759f $X=22 $Y=1.7
+ $X2=0 $Y2=0
cc_3563 N_A_3797_297#_c_6020_n N_A_3799_47#_c_7421_n 0.0247972f $X=20.895
+ $Y=1.58 $X2=0 $Y2=0
cc_3564 N_A_3797_297#_c_6034_n N_A_3799_47#_c_7427_n 6.95815e-19 $X=20.07
+ $Y=1.66 $X2=0 $Y2=0
cc_3565 N_A_3797_591#_c_6142_n N_A_3799_911#_c_7503_n 0.0247972f $X=20.895
+ $Y=3.86 $X2=0 $Y2=0
cc_3566 N_A_3797_591#_c_6156_n N_A_3799_911#_c_7510_n 6.95815e-19 $X=20.07
+ $Y=3.78 $X2=0 $Y2=0
cc_3567 N_VGND_c_6370_n N_A_405_66#_M1065_d 0.00215201f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3568 N_VGND_c_6370_n N_A_405_66#_M1151_d 0.00215201f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3569 N_VGND_c_6268_n N_A_405_66#_c_6926_n 0.00696245f $X=1.275 $Y=0.445 $X2=0
+ $Y2=0
cc_3570 N_VGND_c_6312_n N_A_405_66#_c_6927_n 0.0422314f $X=4.185 $Y=0 $X2=0
+ $Y2=0
cc_3571 N_VGND_c_6370_n N_A_405_66#_c_6927_n 0.0219908f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3572 N_VGND_c_6268_n N_A_405_66#_c_6928_n 0.00694621f $X=1.275 $Y=0.445 $X2=0
+ $Y2=0
cc_3573 N_VGND_c_6312_n N_A_405_66#_c_6928_n 0.0167092f $X=4.185 $Y=0 $X2=0
+ $Y2=0
cc_3574 N_VGND_c_6370_n N_A_405_66#_c_6928_n 0.00841721f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3575 N_VGND_c_6270_n N_A_405_66#_c_6929_n 0.0147456f $X=4.35 $Y=0.38 $X2=0
+ $Y2=0
cc_3576 N_VGND_c_6312_n N_A_405_66#_c_6929_n 0.0614775f $X=4.185 $Y=0 $X2=0
+ $Y2=0
cc_3577 N_VGND_c_6370_n N_A_405_66#_c_6929_n 0.0325967f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3578 N_VGND_c_6270_n N_A_405_66#_c_6930_n 0.00959666f $X=4.35 $Y=0.38 $X2=0
+ $Y2=0
cc_3579 N_VGND_M1065_s N_A_405_66#_c_6931_n 0.00692362f $X=4.225 $Y=0.235 $X2=0
+ $Y2=0
cc_3580 N_VGND_c_6270_n N_A_405_66#_c_6931_n 0.0190091f $X=4.35 $Y=0.38 $X2=0
+ $Y2=0
cc_3581 N_VGND_c_6312_n N_A_405_66#_c_6931_n 0.00262594f $X=4.185 $Y=0 $X2=0
+ $Y2=0
cc_3582 N_VGND_c_6340_n N_A_405_66#_c_6931_n 0.0020257f $X=5.105 $Y=0 $X2=0
+ $Y2=0
cc_3583 N_VGND_c_6370_n N_A_405_66#_c_6931_n 0.00940109f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3584 N_VGND_c_6340_n N_A_405_66#_c_6951_n 0.0188215f $X=5.105 $Y=0 $X2=0
+ $Y2=0
cc_3585 N_VGND_c_6370_n N_A_405_66#_c_6951_n 0.0121968f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3586 N_VGND_M1097_s N_A_405_66#_c_6933_n 0.00501873f $X=5.055 $Y=0.235 $X2=0
+ $Y2=0
cc_3587 N_VGND_c_6272_n N_A_405_66#_c_6933_n 0.0199861f $X=5.24 $Y=0.38 $X2=0
+ $Y2=0
cc_3588 N_VGND_c_6340_n N_A_405_66#_c_6933_n 0.0020257f $X=5.105 $Y=0 $X2=0
+ $Y2=0
cc_3589 N_VGND_c_6342_n N_A_405_66#_c_6933_n 0.0020257f $X=6.045 $Y=0 $X2=0
+ $Y2=0
cc_3590 N_VGND_c_6370_n N_A_405_66#_c_6933_n 0.00880092f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3591 N_VGND_c_6342_n N_A_405_66#_c_6960_n 0.0188215f $X=6.045 $Y=0 $X2=0
+ $Y2=0
cc_3592 N_VGND_c_6370_n N_A_405_66#_c_6960_n 0.0121968f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3593 N_VGND_c_6312_n N_A_405_66#_c_6945_n 0.0113631f $X=4.185 $Y=0 $X2=0
+ $Y2=0
cc_3594 N_VGND_c_6370_n N_A_405_66#_c_6945_n 0.00572388f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3595 N_VGND_c_6371_n N_A_405_918#_M1030_d 0.00215201f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3596 N_VGND_c_6371_n N_A_405_918#_M1068_d 0.00215201f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3597 N_VGND_c_6269_n N_A_405_918#_c_7010_n 0.00696245f $X=1.275 $Y=4.995
+ $X2=0 $Y2=0
cc_3598 N_VGND_c_6314_n N_A_405_918#_c_7011_n 0.0422314f $X=4.185 $Y=5.44 $X2=0
+ $Y2=0
cc_3599 N_VGND_c_6371_n N_A_405_918#_c_7011_n 0.0219908f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3600 N_VGND_c_6269_n N_A_405_918#_c_7012_n 0.00694621f $X=1.275 $Y=4.995
+ $X2=0 $Y2=0
cc_3601 N_VGND_c_6314_n N_A_405_918#_c_7012_n 0.0167092f $X=4.185 $Y=5.44 $X2=0
+ $Y2=0
cc_3602 N_VGND_c_6371_n N_A_405_918#_c_7012_n 0.00841721f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3603 N_VGND_c_6271_n N_A_405_918#_c_7013_n 0.0147456f $X=4.35 $Y=5.06 $X2=0
+ $Y2=0
cc_3604 N_VGND_c_6314_n N_A_405_918#_c_7013_n 0.0614775f $X=4.185 $Y=5.44 $X2=0
+ $Y2=0
cc_3605 N_VGND_c_6371_n N_A_405_918#_c_7013_n 0.0325967f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3606 N_VGND_c_6271_n N_A_405_918#_c_7014_n 0.00959666f $X=4.35 $Y=5.06 $X2=0
+ $Y2=0
cc_3607 N_VGND_M1030_s N_A_405_918#_c_7015_n 0.00692362f $X=4.225 $Y=4.555 $X2=0
+ $Y2=0
cc_3608 N_VGND_c_6271_n N_A_405_918#_c_7015_n 0.0190091f $X=4.35 $Y=5.06 $X2=0
+ $Y2=0
cc_3609 N_VGND_c_6314_n N_A_405_918#_c_7015_n 0.00262594f $X=4.185 $Y=5.44 $X2=0
+ $Y2=0
cc_3610 N_VGND_c_6341_n N_A_405_918#_c_7015_n 0.0020257f $X=5.105 $Y=5.44 $X2=0
+ $Y2=0
cc_3611 N_VGND_c_6371_n N_A_405_918#_c_7015_n 0.00940109f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3612 N_VGND_M1059_s N_A_405_918#_c_7035_n 0.00501873f $X=5.055 $Y=4.555 $X2=0
+ $Y2=0
cc_3613 N_VGND_c_6273_n N_A_405_918#_c_7035_n 0.0199861f $X=5.24 $Y=5.06 $X2=0
+ $Y2=0
cc_3614 N_VGND_c_6341_n N_A_405_918#_c_7035_n 0.0020257f $X=5.105 $Y=5.44 $X2=0
+ $Y2=0
cc_3615 N_VGND_c_6343_n N_A_405_918#_c_7035_n 0.0020257f $X=6.045 $Y=5.44 $X2=0
+ $Y2=0
cc_3616 N_VGND_c_6371_n N_A_405_918#_c_7035_n 0.00880092f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3617 N_VGND_c_6314_n N_A_405_918#_c_7029_n 0.0113631f $X=4.185 $Y=5.44 $X2=0
+ $Y2=0
cc_3618 N_VGND_c_6371_n N_A_405_918#_c_7029_n 0.00572388f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3619 N_VGND_c_6341_n N_A_405_918#_c_7017_n 0.0188215f $X=5.105 $Y=5.44 $X2=0
+ $Y2=0
cc_3620 N_VGND_c_6371_n N_A_405_918#_c_7017_n 0.0121968f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3621 N_VGND_c_6343_n N_A_405_918#_c_7018_n 0.0188215f $X=6.045 $Y=5.44 $X2=0
+ $Y2=0
cc_3622 N_VGND_c_6371_n N_A_405_918#_c_7018_n 0.0121968f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3623 N_VGND_c_6370_n N_A_1315_47#_M1013_s 0.00215201f $X=24.61 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_3624 N_VGND_c_6370_n N_A_1315_47#_M1069_s 0.00215201f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3625 N_VGND_c_6344_n N_A_1315_47#_c_7100_n 0.0188215f $X=7.045 $Y=0 $X2=0
+ $Y2=0
cc_3626 N_VGND_c_6370_n N_A_1315_47#_c_7100_n 0.0121968f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3627 N_VGND_M1037_d N_A_1315_47#_c_7103_n 0.00501873f $X=6.995 $Y=0.235 $X2=0
+ $Y2=0
cc_3628 N_VGND_c_6276_n N_A_1315_47#_c_7103_n 0.0199861f $X=7.18 $Y=0.38 $X2=0
+ $Y2=0
cc_3629 N_VGND_c_6278_n N_A_1315_47#_c_7103_n 0.0020257f $X=7.985 $Y=0 $X2=0
+ $Y2=0
cc_3630 N_VGND_c_6344_n N_A_1315_47#_c_7103_n 0.0020257f $X=7.045 $Y=0 $X2=0
+ $Y2=0
cc_3631 N_VGND_c_6370_n N_A_1315_47#_c_7103_n 0.00880092f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3632 N_VGND_c_6278_n N_A_1315_47#_c_7111_n 0.0188215f $X=7.985 $Y=0 $X2=0
+ $Y2=0
cc_3633 N_VGND_c_6370_n N_A_1315_47#_c_7111_n 0.0121968f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3634 N_VGND_M1150_d N_A_1315_47#_c_7093_n 0.00692362f $X=7.935 $Y=0.235 $X2=0
+ $Y2=0
cc_3635 N_VGND_c_6278_n N_A_1315_47#_c_7093_n 0.0020257f $X=7.985 $Y=0 $X2=0
+ $Y2=0
cc_3636 N_VGND_c_6280_n N_A_1315_47#_c_7093_n 0.0190091f $X=8.07 $Y=0.38 $X2=0
+ $Y2=0
cc_3637 N_VGND_c_6316_n N_A_1315_47#_c_7093_n 0.00262594f $X=10.94 $Y=0 $X2=0
+ $Y2=0
cc_3638 N_VGND_c_6370_n N_A_1315_47#_c_7093_n 0.00940109f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3639 N_VGND_c_6280_n N_A_1315_47#_c_7094_n 0.00959666f $X=8.07 $Y=0.38 $X2=0
+ $Y2=0
cc_3640 N_VGND_c_6316_n N_A_1315_47#_c_7095_n 0.0422314f $X=10.94 $Y=0 $X2=0
+ $Y2=0
cc_3641 N_VGND_c_6370_n N_A_1315_47#_c_7095_n 0.0222193f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3642 N_VGND_c_6280_n N_A_1315_47#_c_7096_n 0.0147456f $X=8.07 $Y=0.38 $X2=0
+ $Y2=0
cc_3643 N_VGND_c_6316_n N_A_1315_47#_c_7096_n 0.0192461f $X=10.94 $Y=0 $X2=0
+ $Y2=0
cc_3644 N_VGND_c_6370_n N_A_1315_47#_c_7096_n 0.0103774f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3645 N_VGND_c_6282_n N_A_1315_47#_c_7097_n 0.00694621f $X=11.145 $Y=0.445
+ $X2=0 $Y2=0
cc_3646 N_VGND_c_6316_n N_A_1315_47#_c_7097_n 0.0589406f $X=10.94 $Y=0 $X2=0
+ $Y2=0
cc_3647 N_VGND_c_6370_n N_A_1315_47#_c_7097_n 0.030408f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3648 N_VGND_c_6282_n N_A_1315_47#_c_7098_n 0.00696245f $X=11.145 $Y=0.445
+ $X2=0 $Y2=0
cc_3649 N_VGND_c_6316_n N_A_1315_47#_c_7133_n 0.0113631f $X=10.94 $Y=0 $X2=0
+ $Y2=0
cc_3650 N_VGND_c_6370_n N_A_1315_47#_c_7133_n 0.00572388f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3651 N_VGND_c_6371_n N_A_1315_911#_M1015_d 0.00215201f $X=24.61 $Y=5.44
+ $X2=-0.19 $Y2=-0.24
cc_3652 N_VGND_c_6371_n N_A_1315_911#_M1104_d 0.00215201f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3653 N_VGND_M1047_s N_A_1315_911#_c_7183_n 0.00501873f $X=6.995 $Y=4.555
+ $X2=0 $Y2=0
cc_3654 N_VGND_c_6277_n N_A_1315_911#_c_7183_n 0.0199861f $X=7.18 $Y=5.06 $X2=0
+ $Y2=0
cc_3655 N_VGND_c_6279_n N_A_1315_911#_c_7183_n 0.0020257f $X=7.985 $Y=5.44 $X2=0
+ $Y2=0
cc_3656 N_VGND_c_6345_n N_A_1315_911#_c_7183_n 0.0020257f $X=7.045 $Y=5.44 $X2=0
+ $Y2=0
cc_3657 N_VGND_c_6371_n N_A_1315_911#_c_7183_n 0.00880092f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
cc_3658 N_VGND_M1136_s N_A_1315_911#_c_7175_n 0.00692362f $X=7.935 $Y=4.555
+ $X2=0 $Y2=0
cc_3659 N_VGND_c_6279_n N_A_1315_911#_c_7175_n 0.0020257f $X=7.985 $Y=5.44 $X2=0
+ $Y2=0
cc_3660 N_VGND_c_6281_n N_A_1315_911#_c_7175_n 0.0190091f $X=8.07 $Y=5.06 $X2=0
+ $Y2=0
cc_3661 N_VGND_c_6318_n N_A_1315_911#_c_7175_n 0.00262594f $X=10.94 $Y=5.44
+ $X2=0 $Y2=0
cc_3662 N_VGND_c_6371_n N_A_1315_911#_c_7175_n 0.00940109f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
cc_3663 N_VGND_c_6281_n N_A_1315_911#_c_7176_n 0.00959666f $X=8.07 $Y=5.06 $X2=0
+ $Y2=0
cc_3664 N_VGND_c_6318_n N_A_1315_911#_c_7177_n 0.0422314f $X=10.94 $Y=5.44 $X2=0
+ $Y2=0
cc_3665 N_VGND_c_6371_n N_A_1315_911#_c_7177_n 0.0222193f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3666 N_VGND_c_6281_n N_A_1315_911#_c_7178_n 0.0147456f $X=8.07 $Y=5.06 $X2=0
+ $Y2=0
cc_3667 N_VGND_c_6318_n N_A_1315_911#_c_7178_n 0.0192461f $X=10.94 $Y=5.44 $X2=0
+ $Y2=0
cc_3668 N_VGND_c_6371_n N_A_1315_911#_c_7178_n 0.0103774f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3669 N_VGND_c_6283_n N_A_1315_911#_c_7179_n 0.00694621f $X=11.145 $Y=4.995
+ $X2=0 $Y2=0
cc_3670 N_VGND_c_6318_n N_A_1315_911#_c_7179_n 0.0589406f $X=10.94 $Y=5.44 $X2=0
+ $Y2=0
cc_3671 N_VGND_c_6371_n N_A_1315_911#_c_7179_n 0.030408f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3672 N_VGND_c_6283_n N_A_1315_911#_c_7180_n 0.00696245f $X=11.145 $Y=4.995
+ $X2=0 $Y2=0
cc_3673 N_VGND_c_6345_n N_A_1315_911#_c_7181_n 0.0188215f $X=7.045 $Y=5.44 $X2=0
+ $Y2=0
cc_3674 N_VGND_c_6371_n N_A_1315_911#_c_7181_n 0.0121968f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3675 N_VGND_c_6279_n N_A_1315_911#_c_7182_n 0.0188215f $X=7.985 $Y=5.44 $X2=0
+ $Y2=0
cc_3676 N_VGND_c_6371_n N_A_1315_911#_c_7182_n 0.0121968f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3677 N_VGND_c_6318_n N_A_1315_911#_c_7212_n 0.0113631f $X=10.94 $Y=5.44 $X2=0
+ $Y2=0
cc_3678 N_VGND_c_6371_n N_A_1315_911#_c_7212_n 0.00572388f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
cc_3679 N_VGND_c_6370_n N_A_2889_66#_M1027_s 0.00215201f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3680 N_VGND_c_6370_n N_A_2889_66#_M1045_s 0.00215201f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3681 N_VGND_c_6288_n N_A_2889_66#_c_7254_n 0.00696245f $X=13.695 $Y=0.445
+ $X2=0 $Y2=0
cc_3682 N_VGND_c_6332_n N_A_2889_66#_c_7255_n 0.0422314f $X=16.605 $Y=0 $X2=0
+ $Y2=0
cc_3683 N_VGND_c_6370_n N_A_2889_66#_c_7255_n 0.0219908f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3684 N_VGND_c_6288_n N_A_2889_66#_c_7256_n 0.00694621f $X=13.695 $Y=0.445
+ $X2=0 $Y2=0
cc_3685 N_VGND_c_6332_n N_A_2889_66#_c_7256_n 0.0167092f $X=16.605 $Y=0 $X2=0
+ $Y2=0
cc_3686 N_VGND_c_6370_n N_A_2889_66#_c_7256_n 0.00841721f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3687 N_VGND_c_6290_n N_A_2889_66#_c_7257_n 0.0147456f $X=16.77 $Y=0.38 $X2=0
+ $Y2=0
cc_3688 N_VGND_c_6332_n N_A_2889_66#_c_7257_n 0.0614775f $X=16.605 $Y=0 $X2=0
+ $Y2=0
cc_3689 N_VGND_c_6370_n N_A_2889_66#_c_7257_n 0.0325967f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3690 N_VGND_c_6290_n N_A_2889_66#_c_7258_n 0.00959666f $X=16.77 $Y=0.38 $X2=0
+ $Y2=0
cc_3691 N_VGND_M1027_d N_A_2889_66#_c_7259_n 0.00692362f $X=16.645 $Y=0.235
+ $X2=0 $Y2=0
cc_3692 N_VGND_c_6290_n N_A_2889_66#_c_7259_n 0.0190091f $X=16.77 $Y=0.38 $X2=0
+ $Y2=0
cc_3693 N_VGND_c_6332_n N_A_2889_66#_c_7259_n 0.00262594f $X=16.605 $Y=0 $X2=0
+ $Y2=0
cc_3694 N_VGND_c_6346_n N_A_2889_66#_c_7259_n 0.0020257f $X=17.525 $Y=0 $X2=0
+ $Y2=0
cc_3695 N_VGND_c_6370_n N_A_2889_66#_c_7259_n 0.00940109f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3696 N_VGND_c_6346_n N_A_2889_66#_c_7279_n 0.0188215f $X=17.525 $Y=0 $X2=0
+ $Y2=0
cc_3697 N_VGND_c_6370_n N_A_2889_66#_c_7279_n 0.0121968f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3698 N_VGND_M1034_d N_A_2889_66#_c_7261_n 0.00501873f $X=17.475 $Y=0.235
+ $X2=0 $Y2=0
cc_3699 N_VGND_c_6292_n N_A_2889_66#_c_7261_n 0.0199861f $X=17.66 $Y=0.38 $X2=0
+ $Y2=0
cc_3700 N_VGND_c_6346_n N_A_2889_66#_c_7261_n 0.0020257f $X=17.525 $Y=0 $X2=0
+ $Y2=0
cc_3701 N_VGND_c_6348_n N_A_2889_66#_c_7261_n 0.0020257f $X=18.465 $Y=0 $X2=0
+ $Y2=0
cc_3702 N_VGND_c_6370_n N_A_2889_66#_c_7261_n 0.00880092f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3703 N_VGND_c_6348_n N_A_2889_66#_c_7288_n 0.0188215f $X=18.465 $Y=0 $X2=0
+ $Y2=0
cc_3704 N_VGND_c_6370_n N_A_2889_66#_c_7288_n 0.0121968f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3705 N_VGND_c_6332_n N_A_2889_66#_c_7273_n 0.0113631f $X=16.605 $Y=0 $X2=0
+ $Y2=0
cc_3706 N_VGND_c_6370_n N_A_2889_66#_c_7273_n 0.00572388f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3707 N_VGND_c_6371_n N_A_2889_918#_M1033_s 0.00215201f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3708 N_VGND_c_6371_n N_A_2889_918#_M1106_s 0.00215201f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3709 N_VGND_c_6289_n N_A_2889_918#_c_7338_n 0.00696245f $X=13.695 $Y=4.995
+ $X2=0 $Y2=0
cc_3710 N_VGND_c_6334_n N_A_2889_918#_c_7339_n 0.0422314f $X=16.605 $Y=5.44
+ $X2=0 $Y2=0
cc_3711 N_VGND_c_6371_n N_A_2889_918#_c_7339_n 0.0219908f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3712 N_VGND_c_6289_n N_A_2889_918#_c_7340_n 0.00694621f $X=13.695 $Y=4.995
+ $X2=0 $Y2=0
cc_3713 N_VGND_c_6334_n N_A_2889_918#_c_7340_n 0.0167092f $X=16.605 $Y=5.44
+ $X2=0 $Y2=0
cc_3714 N_VGND_c_6371_n N_A_2889_918#_c_7340_n 0.00841721f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
cc_3715 N_VGND_c_6291_n N_A_2889_918#_c_7341_n 0.0147456f $X=16.77 $Y=5.06 $X2=0
+ $Y2=0
cc_3716 N_VGND_c_6334_n N_A_2889_918#_c_7341_n 0.0614775f $X=16.605 $Y=5.44
+ $X2=0 $Y2=0
cc_3717 N_VGND_c_6371_n N_A_2889_918#_c_7341_n 0.0325967f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3718 N_VGND_c_6291_n N_A_2889_918#_c_7342_n 0.00959666f $X=16.77 $Y=5.06
+ $X2=0 $Y2=0
cc_3719 N_VGND_M1033_d N_A_2889_918#_c_7343_n 0.00692362f $X=16.645 $Y=4.555
+ $X2=0 $Y2=0
cc_3720 N_VGND_c_6291_n N_A_2889_918#_c_7343_n 0.0190091f $X=16.77 $Y=5.06 $X2=0
+ $Y2=0
cc_3721 N_VGND_c_6334_n N_A_2889_918#_c_7343_n 0.00262594f $X=16.605 $Y=5.44
+ $X2=0 $Y2=0
cc_3722 N_VGND_c_6347_n N_A_2889_918#_c_7343_n 0.0020257f $X=17.525 $Y=5.44
+ $X2=0 $Y2=0
cc_3723 N_VGND_c_6371_n N_A_2889_918#_c_7343_n 0.00940109f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
cc_3724 N_VGND_M1077_d N_A_2889_918#_c_7363_n 0.00501873f $X=17.475 $Y=4.555
+ $X2=0 $Y2=0
cc_3725 N_VGND_c_6293_n N_A_2889_918#_c_7363_n 0.0199861f $X=17.66 $Y=5.06 $X2=0
+ $Y2=0
cc_3726 N_VGND_c_6347_n N_A_2889_918#_c_7363_n 0.0020257f $X=17.525 $Y=5.44
+ $X2=0 $Y2=0
cc_3727 N_VGND_c_6349_n N_A_2889_918#_c_7363_n 0.0020257f $X=18.465 $Y=5.44
+ $X2=0 $Y2=0
cc_3728 N_VGND_c_6371_n N_A_2889_918#_c_7363_n 0.00880092f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
cc_3729 N_VGND_c_6334_n N_A_2889_918#_c_7357_n 0.0113631f $X=16.605 $Y=5.44
+ $X2=0 $Y2=0
cc_3730 N_VGND_c_6371_n N_A_2889_918#_c_7357_n 0.00572388f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
cc_3731 N_VGND_c_6347_n N_A_2889_918#_c_7345_n 0.0188215f $X=17.525 $Y=5.44
+ $X2=0 $Y2=0
cc_3732 N_VGND_c_6371_n N_A_2889_918#_c_7345_n 0.0121968f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3733 N_VGND_c_6349_n N_A_2889_918#_c_7346_n 0.0188215f $X=18.465 $Y=5.44
+ $X2=0 $Y2=0
cc_3734 N_VGND_c_6371_n N_A_2889_918#_c_7346_n 0.0121968f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3735 N_VGND_c_6370_n N_A_3799_47#_M1005_d 0.00215201f $X=24.61 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_3736 N_VGND_c_6370_n N_A_3799_47#_M1111_d 0.00215201f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3737 N_VGND_c_6350_n N_A_3799_47#_c_7428_n 0.0188215f $X=19.465 $Y=0 $X2=0
+ $Y2=0
cc_3738 N_VGND_c_6370_n N_A_3799_47#_c_7428_n 0.0121968f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3739 N_VGND_M1081_s N_A_3799_47#_c_7431_n 0.00501873f $X=19.415 $Y=0.235
+ $X2=0 $Y2=0
cc_3740 N_VGND_c_6296_n N_A_3799_47#_c_7431_n 0.0199861f $X=19.6 $Y=0.38 $X2=0
+ $Y2=0
cc_3741 N_VGND_c_6298_n N_A_3799_47#_c_7431_n 0.0020257f $X=20.405 $Y=0 $X2=0
+ $Y2=0
cc_3742 N_VGND_c_6350_n N_A_3799_47#_c_7431_n 0.0020257f $X=19.465 $Y=0 $X2=0
+ $Y2=0
cc_3743 N_VGND_c_6370_n N_A_3799_47#_c_7431_n 0.00880092f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3744 N_VGND_c_6298_n N_A_3799_47#_c_7439_n 0.0188215f $X=20.405 $Y=0 $X2=0
+ $Y2=0
cc_3745 N_VGND_c_6370_n N_A_3799_47#_c_7439_n 0.0121968f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3746 N_VGND_M1159_s N_A_3799_47#_c_7421_n 0.00692362f $X=20.355 $Y=0.235
+ $X2=0 $Y2=0
cc_3747 N_VGND_c_6298_n N_A_3799_47#_c_7421_n 0.0020257f $X=20.405 $Y=0 $X2=0
+ $Y2=0
cc_3748 N_VGND_c_6300_n N_A_3799_47#_c_7421_n 0.0190091f $X=20.49 $Y=0.38 $X2=0
+ $Y2=0
cc_3749 N_VGND_c_6336_n N_A_3799_47#_c_7421_n 0.00262594f $X=23.36 $Y=0 $X2=0
+ $Y2=0
cc_3750 N_VGND_c_6370_n N_A_3799_47#_c_7421_n 0.00940109f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3751 N_VGND_c_6300_n N_A_3799_47#_c_7422_n 0.00959666f $X=20.49 $Y=0.38 $X2=0
+ $Y2=0
cc_3752 N_VGND_c_6336_n N_A_3799_47#_c_7423_n 0.0422314f $X=23.36 $Y=0 $X2=0
+ $Y2=0
cc_3753 N_VGND_c_6370_n N_A_3799_47#_c_7423_n 0.0222193f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3754 N_VGND_c_6300_n N_A_3799_47#_c_7424_n 0.0147456f $X=20.49 $Y=0.38 $X2=0
+ $Y2=0
cc_3755 N_VGND_c_6336_n N_A_3799_47#_c_7424_n 0.0192461f $X=23.36 $Y=0 $X2=0
+ $Y2=0
cc_3756 N_VGND_c_6370_n N_A_3799_47#_c_7424_n 0.0103774f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3757 N_VGND_c_6302_n N_A_3799_47#_c_7425_n 0.00694621f $X=23.565 $Y=0.445
+ $X2=0 $Y2=0
cc_3758 N_VGND_c_6336_n N_A_3799_47#_c_7425_n 0.0589406f $X=23.36 $Y=0 $X2=0
+ $Y2=0
cc_3759 N_VGND_c_6370_n N_A_3799_47#_c_7425_n 0.030408f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3760 N_VGND_c_6302_n N_A_3799_47#_c_7426_n 0.00696245f $X=23.565 $Y=0.445
+ $X2=0 $Y2=0
cc_3761 N_VGND_c_6336_n N_A_3799_47#_c_7461_n 0.0113631f $X=23.36 $Y=0 $X2=0
+ $Y2=0
cc_3762 N_VGND_c_6370_n N_A_3799_47#_c_7461_n 0.00572388f $X=24.61 $Y=0 $X2=0
+ $Y2=0
cc_3763 N_VGND_c_6371_n N_A_3799_911#_M1014_s 0.00215201f $X=24.61 $Y=5.44
+ $X2=-0.19 $Y2=-0.24
cc_3764 N_VGND_c_6371_n N_A_3799_911#_M1026_s 0.00215201f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3765 N_VGND_M1025_d N_A_3799_911#_c_7511_n 0.00501873f $X=19.415 $Y=4.555
+ $X2=0 $Y2=0
cc_3766 N_VGND_c_6297_n N_A_3799_911#_c_7511_n 0.0199861f $X=19.6 $Y=5.06 $X2=0
+ $Y2=0
cc_3767 N_VGND_c_6299_n N_A_3799_911#_c_7511_n 0.0020257f $X=20.405 $Y=5.44
+ $X2=0 $Y2=0
cc_3768 N_VGND_c_6351_n N_A_3799_911#_c_7511_n 0.0020257f $X=19.465 $Y=5.44
+ $X2=0 $Y2=0
cc_3769 N_VGND_c_6371_n N_A_3799_911#_c_7511_n 0.00880092f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
cc_3770 N_VGND_M1098_d N_A_3799_911#_c_7503_n 0.00692362f $X=20.355 $Y=4.555
+ $X2=0 $Y2=0
cc_3771 N_VGND_c_6299_n N_A_3799_911#_c_7503_n 0.0020257f $X=20.405 $Y=5.44
+ $X2=0 $Y2=0
cc_3772 N_VGND_c_6301_n N_A_3799_911#_c_7503_n 0.0190091f $X=20.49 $Y=5.06 $X2=0
+ $Y2=0
cc_3773 N_VGND_c_6338_n N_A_3799_911#_c_7503_n 0.00262594f $X=23.36 $Y=5.44
+ $X2=0 $Y2=0
cc_3774 N_VGND_c_6371_n N_A_3799_911#_c_7503_n 0.00940109f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
cc_3775 N_VGND_c_6301_n N_A_3799_911#_c_7504_n 0.00959666f $X=20.49 $Y=5.06
+ $X2=0 $Y2=0
cc_3776 N_VGND_c_6338_n N_A_3799_911#_c_7505_n 0.0422314f $X=23.36 $Y=5.44 $X2=0
+ $Y2=0
cc_3777 N_VGND_c_6371_n N_A_3799_911#_c_7505_n 0.0222193f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3778 N_VGND_c_6301_n N_A_3799_911#_c_7506_n 0.0147456f $X=20.49 $Y=5.06 $X2=0
+ $Y2=0
cc_3779 N_VGND_c_6338_n N_A_3799_911#_c_7506_n 0.0192461f $X=23.36 $Y=5.44 $X2=0
+ $Y2=0
cc_3780 N_VGND_c_6371_n N_A_3799_911#_c_7506_n 0.0103774f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3781 N_VGND_c_6303_n N_A_3799_911#_c_7507_n 0.00694621f $X=23.565 $Y=4.995
+ $X2=0 $Y2=0
cc_3782 N_VGND_c_6338_n N_A_3799_911#_c_7507_n 0.0589406f $X=23.36 $Y=5.44 $X2=0
+ $Y2=0
cc_3783 N_VGND_c_6371_n N_A_3799_911#_c_7507_n 0.030408f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3784 N_VGND_c_6303_n N_A_3799_911#_c_7508_n 0.00696245f $X=23.565 $Y=4.995
+ $X2=0 $Y2=0
cc_3785 N_VGND_c_6351_n N_A_3799_911#_c_7509_n 0.0188215f $X=19.465 $Y=5.44
+ $X2=0 $Y2=0
cc_3786 N_VGND_c_6371_n N_A_3799_911#_c_7509_n 0.0121968f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3787 N_VGND_c_6299_n N_A_3799_911#_c_7510_n 0.0188215f $X=20.405 $Y=5.44
+ $X2=0 $Y2=0
cc_3788 N_VGND_c_6371_n N_A_3799_911#_c_7510_n 0.0121968f $X=24.61 $Y=5.44 $X2=0
+ $Y2=0
cc_3789 N_VGND_c_6338_n N_A_3799_911#_c_7540_n 0.0113631f $X=23.36 $Y=5.44 $X2=0
+ $Y2=0
cc_3790 N_VGND_c_6371_n N_A_3799_911#_c_7540_n 0.00572388f $X=24.61 $Y=5.44
+ $X2=0 $Y2=0
