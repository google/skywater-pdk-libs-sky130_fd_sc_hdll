* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_27_47# B1 a_1088_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A1 a_118_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y C1 a_1464_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 Y C1 a_886_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y A2 a_118_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_118_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_886_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_1088_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 Y A2 a_118_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_27_47# B1 a_886_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_118_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 a_886_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_118_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 VPWR A1 a_118_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_118_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 a_1464_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
