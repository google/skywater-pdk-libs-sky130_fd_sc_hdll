* File: sky130_fd_sc_hdll__or2_4.pex.spice
* Created: Wed Sep  2 08:47:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR2_4%B 1 3 4 6 7 8 14
r29 14 15 4.66022 $w=3.62e-07 $l=3.5e-08 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.555 $Y2=1.202
r30 12 14 34.6188 $w=3.62e-07 $l=2.6e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.52 $Y2=1.202
r31 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r32 7 8 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.217 $Y=0.85
+ $X2=0.217 $Y2=1.16
r33 4 15 19.0988 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.555 $Y=1.41
+ $X2=0.555 $Y2=1.202
r34 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.555 $Y=1.41
+ $X2=0.555 $Y2=1.985
r35 1 14 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_4%A 1 3 4 6 7 16
c31 4 0 1.39882e-19 $X=0.965 $Y=1.41
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r33 7 16 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=1.155
+ $Y2=1.16
r34 7 11 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=1
+ $Y2=1.16
r35 4 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=1.025 $Y2=1.16
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r37 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=1.025 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_4%A_35_297# 1 2 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 33 36 37 39 40 43 47 49 63
c114 40 0 1.07308e-19 $X=1.637 $Y=1.495
c115 39 0 1.39882e-19 $X=1.637 $Y=1.245
c116 36 0 1.05688e-19 $X=0.63 $Y=1.495
r117 63 64 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.93 $Y=1.202
+ $X2=2.955 $Y2=1.202
r118 62 63 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=2.46 $Y=1.202
+ $X2=2.93 $Y2=1.202
r119 59 60 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=1.99 $Y=1.202
+ $X2=2.435 $Y2=1.202
r120 58 59 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.965 $Y=1.202
+ $X2=1.99 $Y2=1.202
r121 55 56 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.495 $Y=1.202
+ $X2=1.52 $Y2=1.202
r122 54 58 31.0968 $w=3.72e-07 $l=2.4e-07 $layer=POLY_cond $X=1.725 $Y=1.202
+ $X2=1.965 $Y2=1.202
r123 54 56 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=1.725 $Y=1.202
+ $X2=1.52 $Y2=1.202
r124 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.16 $X2=1.725 $Y2=1.16
r125 49 51 14.6716 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=0.705 $Y=0.4
+ $X2=0.705 $Y2=0.825
r126 44 62 0.647849 $w=3.72e-07 $l=5e-09 $layer=POLY_cond $X=2.455 $Y=1.202
+ $X2=2.46 $Y2=1.202
r127 44 60 2.5914 $w=3.72e-07 $l=2e-08 $layer=POLY_cond $X=2.455 $Y=1.202
+ $X2=2.435 $Y2=1.202
r128 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.455
+ $Y=1.16 $X2=2.455 $Y2=1.16
r129 41 53 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.765 $Y=1.16
+ $X2=1.637 $Y2=1.16
r130 41 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.765 $Y=1.16
+ $X2=2.455 $Y2=1.16
r131 39 53 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.637 $Y=1.245
+ $X2=1.637 $Y2=1.16
r132 39 40 11.2985 $w=2.53e-07 $l=2.5e-07 $layer=LI1_cond $X=1.637 $Y=1.245
+ $X2=1.637 $Y2=1.495
r133 38 47 3.3845 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=0.745 $Y=1.58
+ $X2=0.45 $Y2=1.58
r134 37 40 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.51 $Y=1.58
+ $X2=1.637 $Y2=1.495
r135 37 38 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.51 $Y=1.58
+ $X2=0.745 $Y2=1.58
r136 36 47 3.19717 $w=2.95e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.63 $Y=1.495
+ $X2=0.45 $Y2=1.58
r137 36 51 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=0.63 $Y=1.495
+ $X2=0.63 $Y2=0.825
r138 31 47 3.19717 $w=2.95e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.335 $Y=1.665
+ $X2=0.45 $Y2=1.58
r139 31 33 20.3278 $w=3.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.335 $Y=1.665
+ $X2=0.335 $Y2=2.3
r140 28 64 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.955 $Y=0.995
+ $X2=2.955 $Y2=1.202
r141 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.955 $Y=0.995
+ $X2=2.955 $Y2=0.56
r142 25 63 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.93 $Y=1.41
+ $X2=2.93 $Y2=1.202
r143 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.93 $Y=1.41
+ $X2=2.93 $Y2=1.985
r144 22 62 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.46 $Y=1.41
+ $X2=2.46 $Y2=1.202
r145 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.46 $Y=1.41
+ $X2=2.46 $Y2=1.985
r146 19 60 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.435 $Y=0.995
+ $X2=2.435 $Y2=1.202
r147 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.435 $Y=0.995
+ $X2=2.435 $Y2=0.56
r148 16 59 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.202
r149 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.985
r150 13 58 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.965 $Y=0.995
+ $X2=1.965 $Y2=1.202
r151 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.965 $Y=0.995
+ $X2=1.965 $Y2=0.56
r152 10 56 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.52 $Y=1.41
+ $X2=1.52 $Y2=1.202
r153 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.52 $Y=1.41
+ $X2=1.52 $Y2=1.985
r154 7 55 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=1.202
r155 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=0.56
r156 2 47 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.485 $X2=0.32 $Y2=1.62
r157 2 33 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.485 $X2=0.32 $Y2=2.3
r158 1 49 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_4%VPWR 1 2 3 12 16 20 23 24 26 27 29 30 31 47
+ 48
r54 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 45 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 34 38 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 31 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 31 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 29 44 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.08 $Y=2.72 $X2=2.99
+ $Y2=2.72
r65 29 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.72
+ $X2=3.165 $Y2=2.72
r66 28 47 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.25 $Y=2.72 $X2=3.45
+ $Y2=2.72
r67 28 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=2.72
+ $X2=3.165 $Y2=2.72
r68 26 41 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.14 $Y=2.72 $X2=2.07
+ $Y2=2.72
r69 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.72
+ $X2=2.225 $Y2=2.72
r70 25 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.99 $Y2=2.72
r71 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.225 $Y2=2.72
r72 23 38 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.16 $Y=2.72 $X2=1.15
+ $Y2=2.72
r73 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=2.72
+ $X2=1.245 $Y2=2.72
r74 22 41 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.33 $Y=2.72
+ $X2=2.07 $Y2=2.72
r75 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=2.72
+ $X2=1.245 $Y2=2.72
r76 18 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=2.635
+ $X2=3.165 $Y2=2.72
r77 18 20 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.165 $Y=2.635
+ $X2=3.165 $Y2=2
r78 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.72
r79 14 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.34
r80 10 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=2.635
+ $X2=1.245 $Y2=2.72
r81 10 12 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.245 $Y=2.635
+ $X2=1.245 $Y2=2.01
r82 3 20 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.02
+ $Y=1.485 $X2=3.165 $Y2=2
r83 2 16 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.485 $X2=2.225 $Y2=2.34
r84 1 12 300 $w=1.7e-07 $l=6.12679e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.245 $Y2=2.01
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_4%X 1 2 3 4 15 19 20 21 25 29 32 35 37 47
c77 3 0 1.07308e-19 $X=1.61 $Y=1.485
r78 43 44 0.822102 $w=3.71e-07 $l=2.5e-08 $layer=LI1_cond $X=2.695 $Y=1.75
+ $X2=2.72 $Y2=1.75
r79 40 47 0.0657682 $w=3.71e-07 $l=3.59861e-08 $layer=LI1_cond $X=2.997 $Y=1.495
+ $X2=2.995 $Y2=1.53
r80 37 47 0.16442 $w=3.71e-07 $l=2.73861e-08 $layer=LI1_cond $X=2.99 $Y=1.555
+ $X2=2.995 $Y2=1.53
r81 37 44 8.87871 $w=3.71e-07 $l=3.5433e-07 $layer=LI1_cond $X=2.99 $Y=1.555
+ $X2=2.72 $Y2=1.75
r82 37 40 0.835104 $w=3.43e-07 $l=2.5e-08 $layer=LI1_cond $X=2.997 $Y=1.47
+ $X2=2.997 $Y2=1.495
r83 35 37 18.8733 $w=3.43e-07 $l=5.65e-07 $layer=LI1_cond $X=2.997 $Y=0.905
+ $X2=2.997 $Y2=1.47
r84 27 44 0.569786 $w=3.8e-07 $l=2.55e-07 $layer=LI1_cond $X=2.72 $Y=2.005
+ $X2=2.72 $Y2=1.75
r85 27 29 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.72 $Y=2.005
+ $X2=2.72 $Y2=2.34
r86 23 35 18.0717 $w=1.68e-07 $l=2.77e-07 $layer=LI1_cond $X=2.72 $Y=0.82
+ $X2=2.997 $Y2=0.82
r87 23 25 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.72 $Y=0.735
+ $X2=2.72 $Y2=0.4
r88 22 32 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.97 $Y=1.92 $X2=1.78
+ $Y2=1.92
r89 21 43 9.04258 $w=3.71e-07 $l=2.38642e-07 $layer=LI1_cond $X=2.53 $Y=1.92
+ $X2=2.695 $Y2=1.75
r90 21 22 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.53 $Y=1.92
+ $X2=1.97 $Y2=1.92
r91 19 23 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.53 $Y=0.82
+ $X2=2.72 $Y2=0.82
r92 19 20 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.53 $Y=0.82
+ $X2=1.97 $Y2=0.82
r93 13 20 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=1.78 $Y=0.735
+ $X2=1.97 $Y2=0.82
r94 13 15 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.78 $Y=0.735
+ $X2=1.78 $Y2=0.4
r95 4 43 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.55
+ $Y=1.485 $X2=2.695 $Y2=1.66
r96 4 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.55
+ $Y=1.485 $X2=2.695 $Y2=2.34
r97 3 32 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.61
+ $Y=1.485 $X2=1.755 $Y2=2
r98 2 25 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.51
+ $Y=0.235 $X2=2.695 $Y2=0.4
r99 1 15 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.235 $X2=1.755 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_4%VGND 1 2 3 4 13 15 19 23 27 30 31 33 34 36
+ 37 38 51 52
r58 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r59 49 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r60 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r61 46 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r62 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r63 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r64 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r65 40 55 3.93736 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r66 40 42 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=1.15
+ $Y2=0
r67 38 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r68 38 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r69 36 48 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.99
+ $Y2=0
r70 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.165
+ $Y2=0
r71 35 51 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.45
+ $Y2=0
r72 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.165
+ $Y2=0
r73 33 45 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.07
+ $Y2=0
r74 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.225
+ $Y2=0
r75 32 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.99
+ $Y2=0
r76 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.225
+ $Y2=0
r77 30 42 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.15
+ $Y2=0
r78 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.245
+ $Y2=0
r79 29 45 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.33 $Y=0 $X2=2.07
+ $Y2=0
r80 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=0 $X2=1.245
+ $Y2=0
r81 25 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=0.085
+ $X2=3.165 $Y2=0
r82 25 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.165 $Y=0.085
+ $X2=3.165 $Y2=0.4
r83 21 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0
r84 21 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0.4
r85 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r86 17 19 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.575
r87 13 55 3.14078 $w=2.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.172 $Y2=0
r88 13 15 15.606 $w=2.38e-07 $l=3.25e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.41
r89 4 27 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.03
+ $Y=0.235 $X2=3.165 $Y2=0.4
r90 3 23 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.235 $X2=2.225 $Y2=0.4
r91 2 19 182 $w=1.7e-07 $l=4.40227e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.245 $Y2=0.575
r92 1 15 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.41
.ends

