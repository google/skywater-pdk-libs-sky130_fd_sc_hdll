* File: sky130_fd_sc_hdll__diode_4.pxi.spice
* Created: Wed Sep  2 08:28:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__DIODE_4%DIODE N_DIODE_D0_noxref_neg DIODE DIODE DIODE
+ DIODE DIODE DIODE N_DIODE_c_8_n PM_SKY130_FD_SC_HDLL__DIODE_4%DIODE
x_PM_SKY130_FD_SC_HDLL__DIODE_4%VGND VGND N_VGND_c_15_n N_VGND_c_16_n
+ PM_SKY130_FD_SC_HDLL__DIODE_4%VGND
x_PM_SKY130_FD_SC_HDLL__DIODE_4%VPWR VPWR N_VPWR_c_21_n N_VPWR_c_20_n
+ PM_SKY130_FD_SC_HDLL__DIODE_4%VPWR
cc_1 VNB N_DIODE_c_8_n 0.115659f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=0.37
cc_2 VNB N_VGND_c_15_n 0.0472107f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.785
cc_3 VNB N_VGND_c_16_n 0.123857f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=2.125
cc_4 VNB N_VPWR_c_20_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=2.125
cc_5 VPB N_DIODE_c_8_n 0.178198f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=0.37
cc_6 VPB N_VPWR_c_21_n 0.0472107f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.785
cc_7 VPB N_VPWR_c_20_n 0.0563576f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=2.125
cc_8 N_DIODE_c_8_n N_VGND_c_15_n 0.117485f $X=0.285 $Y=0.37 $X2=0 $Y2=0
cc_9 N_DIODE_D0_noxref_neg N_VGND_c_16_n 0.0146005f $X=0.155 $Y=0.195 $X2=0
+ $Y2=0
cc_10 N_DIODE_c_8_n N_VGND_c_16_n 0.0642376f $X=0.285 $Y=0.37 $X2=0 $Y2=0
cc_11 N_DIODE_c_8_n N_VPWR_c_21_n 0.119588f $X=0.285 $Y=0.37 $X2=0 $Y2=0
cc_12 N_DIODE_c_8_n N_VPWR_c_20_n 0.0642376f $X=0.285 $Y=0.37 $X2=0 $Y2=0
