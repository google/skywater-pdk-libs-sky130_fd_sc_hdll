* File: sky130_fd_sc_hdll__and3b_4.spice
* Created: Thu Aug 27 18:58:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and3b_4.pex.spice"
.subckt sky130_fd_sc_hdll__and3b_4  VNB VPB B C A_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A_N	A_N
* C	C
* B	B
* VPB	VPB
* VNB	VNB
MM1009 A_162_47# N_A_98_199#_M1009_g N_A_56_297#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.138125 AS=0.23075 PD=1.075 PS=2.01 NRD=29.076 NRS=9.228 M=1
+ R=4.33333 SA=75000.3 SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1014 A_277_47# N_B_M1014_g A_162_47# VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.138125 PD=0.93 PS=1.075 NRD=15.684 NRS=29.076 M=1 R=4.33333 SA=75000.9
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_C_M1000_g A_277_47# VNB NSHORT L=0.15 W=0.65 AD=0.138125
+ AS=0.091 PD=1.075 PS=0.93 NRD=25.836 NRS=15.684 M=1 R=4.33333 SA=75001.3
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1004_d N_A_56_297#_M1004_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.138125 PD=0.98 PS=1.075 NRD=9.228 NRS=0.912 M=1 R=4.33333
+ SA=75001.9 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1004_d N_A_56_297#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=3.684 M=1 R=4.33333 SA=75002.3
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1008_d N_A_56_297#_M1008_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.10725 PD=1.03 PS=0.98 NRD=9.228 NRS=5.532 M=1 R=4.33333
+ SA=75002.8 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1008_d N_A_56_297#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.144428 PD=1.03 PS=1.28785 NRD=9.228 NRS=0 M=1 R=4.33333
+ SA=75003.3 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_A_98_199#_M1013_d N_A_N_M1013_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1743 AS=0.0933224 PD=1.67 PS=0.83215 NRD=37.14 NRS=47.76 M=1 R=2.8
+ SA=75003.9 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_98_199#_M1005_g N_A_56_297#_M1005_s VPB PHIGHVT L=0.18
+ W=1 AD=0.1975 AS=0.34 PD=1.395 PS=2.68 NRD=14.7553 NRS=10.8153 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1015 N_A_56_297#_M1015_d N_B_M1015_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.16 AS=0.1975 PD=1.32 PS=1.395 NRD=5.8903 NRS=7.8603 M=1 R=5.55556
+ SA=90000.8 SB=90002.9 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_C_M1003_g N_A_56_297#_M1015_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1875 AS=0.16 PD=1.375 PS=1.32 NRD=8.8453 NRS=1.9503 M=1 R=5.55556
+ SA=90001.3 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1003_d N_A_56_297#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1875 AS=0.155 PD=1.375 PS=1.31 NRD=9.8303 NRS=3.9203 M=1 R=5.55556
+ SA=90001.9 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_56_297#_M1002_g N_X_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.155 PD=1.29 PS=1.31 NRD=0.9653 NRS=1.9503 M=1 R=5.55556
+ SA=90002.4 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1002_d N_A_56_297#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.15 PD=1.29 PS=1.3 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90002.8
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_56_297#_M1012_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.232887 AS=0.15 PD=1.94366 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90003.3 SB=90000.4 A=0.18 P=2.36 MULT=1
MM1011 N_A_98_199#_M1011_d N_A_N_M1011_g N_VPWR_M1012_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1239 AS=0.0978127 PD=1.43 PS=0.816338 NRD=4.6886 NRS=83.4295 M=1
+ R=2.33333 SA=90003.9 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
pX17_noxref noxref_13 C C PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and3b_4.pxi.spice"
*
.ends
*
*
