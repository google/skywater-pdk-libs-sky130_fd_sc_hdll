# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nor3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.210000 1.075000 2.770000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.285000 1.075000 4.700000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.285000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.925500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 0.255000 1.385000 0.725000 ;
        RECT 1.005000 0.725000 7.245000 0.905000 ;
        RECT 1.945000 0.255000 2.325000 0.725000 ;
        RECT 3.405000 0.255000 3.785000 0.725000 ;
        RECT 4.345000 0.255000 4.725000 0.725000 ;
        RECT 5.285000 0.255000 5.665000 0.725000 ;
        RECT 5.375000 1.455000 7.245000 1.625000 ;
        RECT 5.375000 1.625000 5.625000 2.125000 ;
        RECT 6.225000 0.255000 6.605000 0.725000 ;
        RECT 6.315000 1.625000 6.565000 2.125000 ;
        RECT 6.905000 0.905000 7.245000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.110000  0.255000 0.445000 0.735000 ;
      RECT 0.110000  0.735000 0.835000 0.905000 ;
      RECT 0.110000  1.455000 5.155000 1.625000 ;
      RECT 0.110000  1.625000 0.405000 2.465000 ;
      RECT 0.625000  1.795000 0.875000 2.635000 ;
      RECT 0.665000  0.085000 0.835000 0.555000 ;
      RECT 0.665000  0.905000 0.835000 1.455000 ;
      RECT 1.095000  1.795000 4.685000 1.965000 ;
      RECT 1.095000  1.965000 1.345000 2.465000 ;
      RECT 1.565000  2.135000 1.815000 2.635000 ;
      RECT 1.605000  0.085000 1.775000 0.555000 ;
      RECT 2.035000  1.965000 2.285000 2.465000 ;
      RECT 2.505000  2.135000 2.755000 2.635000 ;
      RECT 2.545000  0.085000 3.235000 0.555000 ;
      RECT 3.025000  2.135000 3.275000 2.295000 ;
      RECT 3.025000  2.295000 7.035000 2.465000 ;
      RECT 3.495000  1.965000 3.745000 2.125000 ;
      RECT 3.965000  2.135000 4.215000 2.295000 ;
      RECT 4.005000  0.085000 4.175000 0.555000 ;
      RECT 4.435000  1.965000 4.685000 2.125000 ;
      RECT 4.905000  1.795000 5.155000 2.295000 ;
      RECT 4.945000  0.085000 5.115000 0.555000 ;
      RECT 4.985000  1.075000 6.720000 1.285000 ;
      RECT 4.985000  1.285000 5.155000 1.455000 ;
      RECT 5.845000  1.795000 6.095000 2.295000 ;
      RECT 5.885000  0.085000 6.055000 0.555000 ;
      RECT 6.785000  1.795000 7.035000 2.295000 ;
      RECT 6.825000  0.085000 6.995000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3b_4
