* File: sky130_fd_sc_hdll__o21bai_2.pex.spice
* Created: Wed Sep  2 08:44:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21BAI_2%B1_N 1 3 4 6 7 15
c26 15 0 1.63168e-19 $X=0.36 $Y=1.19
r27 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.355
+ $Y=1.16 $X2=0.355 $Y2=1.16
r28 7 15 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.23 $Y=1.16
+ $X2=0.355 $Y2=1.16
r29 4 10 39.1844 $w=3.78e-07 $l=2.23596e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.387 $Y2=1.16
r30 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.525 $Y2=0.675
r31 1 10 45.167 $w=3.78e-07 $l=3.01247e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.387 $Y2=1.16
r32 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_2%A_28_297# 1 2 7 9 10 12 13 15 16 18 19 23
+ 26 29 32 37 41
c67 41 0 1.63168e-19 $X=1.63 $Y=1.202
c68 26 0 1.6324e-19 $X=0.782 $Y=1.495
c69 16 0 1.76278e-19 $X=2.1 $Y=0.995
c70 7 0 1.11591e-19 $X=1.035 $Y=1.41
r71 41 42 63.4566 $w=3.57e-07 $l=4.7e-07 $layer=POLY_cond $X=1.63 $Y=1.202
+ $X2=2.1 $Y2=1.202
r72 40 41 16.8768 $w=3.57e-07 $l=1.25e-07 $layer=POLY_cond $X=1.505 $Y=1.202
+ $X2=1.63 $Y2=1.202
r73 32 35 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.265 $Y=1.58
+ $X2=0.265 $Y2=1.725
r74 30 40 44.5546 $w=3.57e-07 $l=3.3e-07 $layer=POLY_cond $X=1.175 $Y=1.202
+ $X2=1.505 $Y2=1.202
r75 30 38 18.902 $w=3.57e-07 $l=1.4e-07 $layer=POLY_cond $X=1.175 $Y=1.202
+ $X2=1.035 $Y2=1.202
r76 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.175
+ $Y=1.16 $X2=1.175 $Y2=1.16
r77 27 37 2.24312 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=0.915 $Y=1.16
+ $X2=0.782 $Y2=1.16
r78 27 29 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.915 $Y=1.16
+ $X2=1.175 $Y2=1.16
r79 25 37 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=0.782 $Y=1.245
+ $X2=0.782 $Y2=1.16
r80 25 26 10.8721 $w=2.63e-07 $l=2.5e-07 $layer=LI1_cond $X=0.782 $Y=1.245
+ $X2=0.782 $Y2=1.495
r81 21 37 4.18896 $w=2.17e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.735 $Y=1.075
+ $X2=0.782 $Y2=1.16
r82 21 23 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.735 $Y=1.075
+ $X2=0.735 $Y2=0.66
r83 20 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.58
+ $X2=0.265 $Y2=1.58
r84 19 26 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=0.65 $Y=1.58
+ $X2=0.782 $Y2=1.495
r85 19 20 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.65 $Y=1.58 $X2=0.35
+ $Y2=1.58
r86 16 42 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.1 $Y=0.995
+ $X2=2.1 $Y2=1.202
r87 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.1 $Y=0.995 $X2=2.1
+ $Y2=0.56
r88 13 41 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.63 $Y=0.995
+ $X2=1.63 $Y2=1.202
r89 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.63 $Y=0.995
+ $X2=1.63 $Y2=0.56
r90 10 40 18.7718 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.505 $Y=1.41
+ $X2=1.505 $Y2=1.202
r91 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.505 $Y=1.41
+ $X2=1.505 $Y2=1.985
r92 7 38 18.7718 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.035 $Y=1.41
+ $X2=1.035 $Y2=1.202
r93 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.035 $Y=1.41
+ $X2=1.035 $Y2=1.985
r94 2 35 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=1.725
r95 1 23 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.465 $X2=0.735 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_2%A2 1 3 4 6 7 9 10 12 13 20
c51 20 0 1.21795e-19 $X=3.015 $Y=1.202
r52 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.015 $Y=1.202
+ $X2=3.04 $Y2=1.202
r53 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=2.78 $Y=1.202
+ $X2=3.015 $Y2=1.202
r54 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=2.545 $Y=1.202
+ $X2=2.78 $Y2=1.202
r55 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.52 $Y=1.202
+ $X2=2.545 $Y2=1.202
r56 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.16 $X2=2.78 $Y2=1.16
r57 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.04 $Y=0.995
+ $X2=3.04 $Y2=1.202
r58 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.04 $Y=0.995
+ $X2=3.04 $Y2=0.56
r59 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=3.015 $Y2=1.202
r60 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=3.015 $Y2=1.985
r61 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.545 $Y2=1.202
r62 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.545 $Y2=1.985
r63 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.52 $Y=0.995
+ $X2=2.52 $Y2=1.202
r64 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.52 $Y=0.995 $X2=2.52
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_2%A1 1 3 4 6 7 9 10 12 13 20 25
c38 25 0 1.21795e-19 $X=3.815 $Y=1.19
r39 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.955 $Y=1.202
+ $X2=3.98 $Y2=1.202
r40 18 20 22.8316 $w=3.8e-07 $l=1.8e-07 $layer=POLY_cond $X=3.775 $Y=1.202
+ $X2=3.955 $Y2=1.202
r41 16 18 36.7842 $w=3.8e-07 $l=2.9e-07 $layer=POLY_cond $X=3.485 $Y=1.202
+ $X2=3.775 $Y2=1.202
r42 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.46 $Y=1.202
+ $X2=3.485 $Y2=1.202
r43 13 25 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=3.775 $Y=1.175
+ $X2=3.815 $Y2=1.175
r44 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=1.16 $X2=3.775 $Y2=1.16
r45 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.98 $Y=0.995
+ $X2=3.98 $Y2=1.202
r46 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.98 $Y=0.995
+ $X2=3.98 $Y2=0.56
r47 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.955 $Y=1.41
+ $X2=3.955 $Y2=1.202
r48 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.955 $Y=1.41
+ $X2=3.955 $Y2=1.985
r49 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.485 $Y2=1.202
r50 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.485 $Y2=1.985
r51 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.46 $Y=0.995
+ $X2=3.46 $Y2=1.202
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.46 $Y=0.995 $X2=3.46
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_2%VPWR 1 2 3 14 18 22 25 26 28 29 30 43 44
+ 47
c63 1 0 1.6324e-19 $X=0.59 $Y=1.485
r64 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r66 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r67 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 38 41 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r69 37 40 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r71 35 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r72 35 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r74 32 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=2.72
+ $X2=0.8 $Y2=2.72
r75 32 34 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.965 $Y=2.72
+ $X2=1.61 $Y2=2.72
r76 30 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 28 40 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.505 $Y=2.72
+ $X2=3.45 $Y2=2.72
r78 28 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.505 $Y=2.72
+ $X2=3.695 $Y2=2.72
r79 27 43 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=4.37 $Y2=2.72
r80 27 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=3.695 $Y2=2.72
r81 25 34 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.62 $Y=2.72 $X2=1.61
+ $Y2=2.72
r82 25 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.62 $Y=2.72
+ $X2=1.745 $Y2=2.72
r83 24 37 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.87 $Y=2.72 $X2=2.07
+ $Y2=2.72
r84 24 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.87 $Y=2.72
+ $X2=1.745 $Y2=2.72
r85 20 29 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.695 $Y=2.635
+ $X2=3.695 $Y2=2.72
r86 20 22 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.695 $Y=2.635
+ $X2=3.695 $Y2=2
r87 16 26 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=2.635
+ $X2=1.745 $Y2=2.72
r88 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.745 $Y=2.635
+ $X2=1.745 $Y2=1.96
r89 12 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=2.635 $X2=0.8
+ $Y2=2.72
r90 12 14 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.8 $Y=2.635
+ $X2=0.8 $Y2=1.96
r91 3 22 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.575
+ $Y=1.485 $X2=3.72 $Y2=2
r92 2 18 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.485 $X2=1.74 $Y2=1.96
r93 1 14 300 $w=1.7e-07 $l=5.70417e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.8 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_2%Y 1 2 3 12 16 20 23 24 27 31
c40 27 0 1.11591e-19 $X=1.84 $Y=0.73
r41 24 31 2.53714 $w=4.93e-07 $l=1.05e-07 $layer=LI1_cond $X=1.757 $Y=1.28
+ $X2=1.757 $Y2=1.385
r42 24 27 13.2898 $w=4.93e-07 $l=5.5e-07 $layer=LI1_cond $X=1.757 $Y=1.28
+ $X2=1.757 $Y2=0.73
r43 22 31 1.44979 $w=4.93e-07 $l=6e-08 $layer=LI1_cond $X=1.757 $Y=1.445
+ $X2=1.757 $Y2=1.385
r44 22 23 2.86771 $w=3.32e-07 $l=2.00035e-07 $layer=LI1_cond $X=1.757 $Y=1.445
+ $X2=1.595 $Y2=1.53
r45 18 20 0.235192 $w=2.43e-07 $l=5e-09 $layer=LI1_cond $X=2.777 $Y=1.615
+ $X2=2.777 $Y2=1.62
r46 17 23 3.83825 $w=1.7e-07 $l=4.1e-07 $layer=LI1_cond $X=2.005 $Y=1.53
+ $X2=1.595 $Y2=1.53
r47 16 18 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.655 $Y=1.53
+ $X2=2.777 $Y2=1.615
r48 16 17 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.655 $Y=1.53
+ $X2=2.005 $Y2=1.53
r49 12 14 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.27 $Y=1.62
+ $X2=1.27 $Y2=2.3
r50 10 23 2.86771 $w=3.32e-07 $l=3.65034e-07 $layer=LI1_cond $X=1.27 $Y=1.615
+ $X2=1.595 $Y2=1.53
r51 10 12 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.27 $Y=1.615
+ $X2=1.27 $Y2=1.62
r52 3 20 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.635
+ $Y=1.485 $X2=2.78 $Y2=1.62
r53 2 14 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.27 $Y2=2.3
r54 2 12 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.27 $Y2=1.62
r55 1 27 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.235 $X2=1.84 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_2%A_437_297# 1 2 3 12 14 15 16 17 18 20 22
r40 20 29 3.02719 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=4.242 $Y=1.665
+ $X2=4.242 $Y2=1.56
r41 20 22 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=4.242 $Y=1.665
+ $X2=4.242 $Y2=2.3
r42 19 25 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.56
+ $X2=3.25 $Y2=1.56
r43 18 29 3.94976 $w=2.1e-07 $l=1.37e-07 $layer=LI1_cond $X=4.105 $Y=1.56
+ $X2=4.242 $Y2=1.56
r44 18 19 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=4.105 $Y=1.56
+ $X2=3.335 $Y2=1.56
r45 17 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=2.295
+ $X2=3.25 $Y2=2.38
r46 16 25 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.25 $Y=1.665
+ $X2=3.25 $Y2=1.56
r47 16 17 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.25 $Y=1.665
+ $X2=3.25 $Y2=2.295
r48 14 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=2.38
+ $X2=3.25 $Y2=2.38
r49 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.165 $Y=2.38
+ $X2=2.435 $Y2=2.38
r50 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.27 $Y=2.295
+ $X2=2.435 $Y2=2.38
r51 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.27 $Y=2.295
+ $X2=2.27 $Y2=1.96
r52 3 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.485 $X2=4.19 $Y2=1.62
r53 3 22 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.485 $X2=4.19 $Y2=2.3
r54 2 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=1.485 $X2=3.25 $Y2=2.3
r55 2 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=1.485 $X2=3.25 $Y2=1.62
r56 1 12 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=2.185
+ $Y=1.485 $X2=2.31 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_2%VGND 1 2 3 10 12 16 20 23 24 26 27 28 41
+ 42
r64 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r65 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r66 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r67 36 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r68 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r69 33 36 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r70 32 35 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r71 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r72 30 45 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.175
+ $Y2=0
r73 30 32 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.69
+ $Y2=0
r74 28 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r75 28 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r76 26 38 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.45
+ $Y2=0
r77 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.72
+ $Y2=0
r78 25 41 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=4.37
+ $Y2=0
r79 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.72
+ $Y2=0
r80 23 35 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.53
+ $Y2=0
r81 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.78
+ $Y2=0
r82 22 38 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=3.45
+ $Y2=0
r83 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.78
+ $Y2=0
r84 18 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0
r85 18 20 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0.39
r86 14 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r87 14 16 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.39
r88 10 45 3.40825 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.175 $Y2=0
r89 10 12 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.66
r90 3 20 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.535
+ $Y=0.235 $X2=3.72 $Y2=0.39
r91 2 16 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.235 $X2=2.78 $Y2=0.39
r92 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.465 $X2=0.265 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_2%A_226_47# 1 2 3 4 13 15 17 19 20 21 25 27
+ 31 39
c72 20 0 1.76278e-19 $X=2.35 $Y=0.725
r73 29 31 9.53255 $w=4.03e-07 $l=3.35e-07 $layer=LI1_cond $X=4.177 $Y=0.725
+ $X2=4.177 $Y2=0.39
r74 28 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.415 $Y=0.815
+ $X2=3.225 $Y2=0.815
r75 27 29 8.21845 $w=1.8e-07 $l=2.42866e-07 $layer=LI1_cond $X=3.975 $Y=0.815
+ $X2=4.177 $Y2=0.725
r76 27 28 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.975 $Y=0.815
+ $X2=3.415 $Y2=0.815
r77 23 39 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.225 $Y=0.725
+ $X2=3.225 $Y2=0.815
r78 23 25 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.225 $Y=0.725
+ $X2=3.225 $Y2=0.39
r79 22 38 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.475 $Y=0.815
+ $X2=2.35 $Y2=0.815
r80 21 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.035 $Y=0.815
+ $X2=3.225 $Y2=0.815
r81 21 22 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.035 $Y=0.815
+ $X2=2.475 $Y2=0.815
r82 20 38 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.35 $Y=0.725 $X2=2.35
+ $Y2=0.815
r83 19 36 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=2.35 $Y=0.475
+ $X2=2.35 $Y2=0.365
r84 19 20 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.35 $Y=0.475
+ $X2=2.35 $Y2=0.725
r85 18 34 3.88917 $w=2.2e-07 $l=1.4e-07 $layer=LI1_cond $X=1.34 $Y=0.365 $X2=1.2
+ $Y2=0.365
r86 17 36 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.225 $Y=0.365
+ $X2=2.35 $Y2=0.365
r87 17 18 46.3596 $w=2.18e-07 $l=8.85e-07 $layer=LI1_cond $X=2.225 $Y=0.365
+ $X2=1.34 $Y2=0.365
r88 13 34 3.05577 $w=2.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.2 $Y=0.475 $X2=1.2
+ $Y2=0.365
r89 13 15 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=1.2 $Y=0.475
+ $X2=1.2 $Y2=0.73
r90 4 31 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.055
+ $Y=0.235 $X2=4.19 $Y2=0.39
r91 3 25 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.115
+ $Y=0.235 $X2=3.25 $Y2=0.39
r92 2 38 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.175
+ $Y=0.235 $X2=2.31 $Y2=0.73
r93 2 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.175
+ $Y=0.235 $X2=2.31 $Y2=0.39
r94 1 34 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.255 $Y2=0.39
r95 1 15 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.255 $Y2=0.73
.ends

