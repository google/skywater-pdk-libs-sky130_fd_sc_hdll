* File: sky130_fd_sc_hdll__nor2b_4.spice
* Created: Wed Sep  2 08:40:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor2b_4.pex.spice"
.subckt sky130_fd_sc_hdll__nor2b_4  VNB VPB A B_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B_N	B_N
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.182
+ AS=0.104 PD=1.86 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2 SB=75003.5
+ A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_M1008_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7 SB=75003.1
+ A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1008_d N_A_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1 SB=75002.6
+ A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_A_M1016_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1016_d N_A_459_21#_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_459_21#_M1005_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1005_d N_A_459_21#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A_459_21#_M1014_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_B_N_M1012_g N_A_459_21#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.208 AS=0.182 PD=1.94 PS=1.86 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_27_297#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1002_d N_A_M1004_g N_A_27_297#_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90003 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_27_297#_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1007_d N_A_M1013_g N_A_27_297#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1000 N_Y_M1000_d N_A_459_21#_M1000_g N_A_27_297#_M1013_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1010 N_Y_M1000_d N_A_459_21#_M1010_g N_A_27_297#_M1010_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1015_d N_A_459_21#_M1015_g N_A_27_297#_M1010_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1017 N_Y_M1015_d N_A_459_21#_M1017_g N_A_27_297#_M1017_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_B_N_M1011_g N_A_459_21#_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.28 PD=2.58 PS=2.56 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hdll__nor2b_4.pxi.spice"
*
.ends
*
*
