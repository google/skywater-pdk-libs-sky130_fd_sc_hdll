* File: sky130_fd_sc_hdll__probe_p_8.pex.spice
* Created: Wed Sep  2 08:50:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__PROBE_P_8%A 1 3 6 8 10 13 17 19 21 22 32 34
c78 32 0 8.84987e-20 $X=0.985 $Y=1.16
c79 8 0 3.25329e-19 $X=0.965 $Y=1.41
r80 34 35 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.212
+ $X2=1.435 $Y2=1.212
r81 33 34 62.4815 $w=3.24e-07 $l=4.2e-07 $layer=POLY_cond $X=0.99 $Y=1.212
+ $X2=1.41 $Y2=1.212
r82 31 33 0.743827 $w=3.24e-07 $l=5e-09 $layer=POLY_cond $X=0.985 $Y=1.212
+ $X2=0.99 $Y2=1.212
r83 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.16 $X2=0.985 $Y2=1.16
r84 29 31 2.97531 $w=3.24e-07 $l=2e-08 $layer=POLY_cond $X=0.965 $Y=1.212
+ $X2=0.985 $Y2=1.212
r85 28 29 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.212
+ $X2=0.965 $Y2=1.212
r86 27 28 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.212
+ $X2=0.52 $Y2=1.212
r87 25 27 28.2654 $w=3.24e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.212
+ $X2=0.495 $Y2=1.212
r88 25 26 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.305
+ $Y=1.16 $X2=0.305 $Y2=1.16
r89 22 32 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=1.175
+ $X2=0.985 $Y2=1.175
r90 22 26 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=0.69 $Y=1.175
+ $X2=0.305 $Y2=1.175
r91 19 35 16.5046 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.212
r92 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r93 15 34 20.7868 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.212
r94 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r95 11 33 20.7868 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=1.212
r96 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=0.56
r97 8 29 16.5046 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.212
r98 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r99 4 28 20.7868 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=1.212
r100 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=0.56
r101 1 27 16.5046 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.212
r102 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBE_P_8%A_27_47# 1 2 3 4 13 15 18 22 24 26 27 29
+ 32 36 38 40 41 43 46 50 52 54 55 57 60 64 66 68 71 77 79 80 81 82 85 91 94 96
+ 102 106 109 111 128
c273 128 0 8.84987e-20 $X=5.17 $Y=1.217
c274 52 0 1.73717e-19 $X=4.255 $Y=1.41
r275 128 129 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.217
+ $X2=5.195 $Y2=1.217
r276 127 128 62.8696 $w=3.22e-07 $l=4.2e-07 $layer=POLY_cond $X=4.75 $Y=1.217
+ $X2=5.17 $Y2=1.217
r277 126 127 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.725 $Y=1.217
+ $X2=4.75 $Y2=1.217
r278 125 126 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=4.255 $Y=1.217
+ $X2=4.725 $Y2=1.217
r279 124 125 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.217
+ $X2=4.255 $Y2=1.217
r280 121 122 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.217
+ $X2=3.81 $Y2=1.217
r281 120 121 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=3.315 $Y=1.217
+ $X2=3.785 $Y2=1.217
r282 119 120 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.217
+ $X2=3.315 $Y2=1.217
r283 118 119 62.8696 $w=3.22e-07 $l=4.2e-07 $layer=POLY_cond $X=2.87 $Y=1.217
+ $X2=3.29 $Y2=1.217
r284 117 118 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=2.87 $Y2=1.217
r285 116 117 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.845 $Y2=1.217
r286 115 116 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r287 112 113 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=1.93 $Y2=1.217
r288 103 124 52.3913 $w=3.22e-07 $l=3.5e-07 $layer=POLY_cond $X=3.88 $Y=1.217
+ $X2=4.23 $Y2=1.217
r289 103 122 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=3.88 $Y=1.217
+ $X2=3.81 $Y2=1.217
r290 102 103 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.88
+ $Y=1.16 $X2=3.88 $Y2=1.16
r291 100 115 25.4472 $w=3.22e-07 $l=1.7e-07 $layer=POLY_cond $X=2.18 $Y=1.217
+ $X2=2.35 $Y2=1.217
r292 100 113 37.4224 $w=3.22e-07 $l=2.5e-07 $layer=POLY_cond $X=2.18 $Y=1.217
+ $X2=1.93 $Y2=1.217
r293 99 102 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=2.18 $Y=1.16
+ $X2=3.88 $Y2=1.16
r294 99 100 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.18
+ $Y=1.16 $X2=2.18 $Y2=1.16
r295 97 111 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.507 $Y2=1.16
r296 97 99 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=2.18 $Y2=1.16
r297 96 106 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.445
+ $X2=1.507 $Y2=1.53
r298 95 111 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.245
+ $X2=1.507 $Y2=1.16
r299 95 96 12.6753 $w=1.73e-07 $l=2e-07 $layer=LI1_cond $X=1.507 $Y=1.245
+ $X2=1.507 $Y2=1.445
r300 94 111 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.075
+ $X2=1.507 $Y2=1.16
r301 93 109 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=0.905
+ $X2=1.507 $Y2=0.82
r302 93 94 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=1.507 $Y=0.905
+ $X2=1.507 $Y2=1.075
r303 89 109 20.0289 $w=1.68e-07 $l=3.07e-07 $layer=LI1_cond $X=1.2 $Y=0.82
+ $X2=1.507 $Y2=0.82
r304 89 91 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.2 $Y2=0.42
r305 85 87 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.2 $Y=1.63 $X2=1.2
+ $Y2=2.31
r306 83 106 20.0289 $w=1.68e-07 $l=3.07e-07 $layer=LI1_cond $X=1.2 $Y=1.53
+ $X2=1.507 $Y2=1.53
r307 83 85 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.2 $Y2=1.63
r308 81 89 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=0.82
+ $X2=1.2 $Y2=0.82
r309 81 82 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.065 $Y=0.82
+ $X2=0.445 $Y2=0.82
r310 79 83 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=1.53
+ $X2=1.2 $Y2=1.53
r311 79 80 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.035 $Y=1.53
+ $X2=0.425 $Y2=1.53
r312 75 82 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.295 $Y=0.735
+ $X2=0.445 $Y2=0.82
r313 75 77 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=0.295 $Y=0.735
+ $X2=0.295 $Y2=0.42
r314 71 73 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r315 69 80 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.425 $Y2=1.53
r316 69 71 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.63
r317 66 129 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.217
r318 66 68 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r319 62 128 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=1.217
r320 62 64 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=0.56
r321 58 127 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=1.217
r322 58 60 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=0.56
r323 55 126 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.217
r324 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r325 52 125 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.217
r326 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r327 48 124 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=1.217
r328 48 50 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=0.56
r329 44 122 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=1.217
r330 44 46 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=0.56
r331 41 121 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.217
r332 41 43 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r333 38 120 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r334 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r335 34 119 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r336 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r337 30 118 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=1.217
r338 30 32 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=0.56
r339 27 117 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r340 27 29 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r341 24 116 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r342 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r343 20 115 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r344 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
r345 16 113 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r346 16 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r347 13 112 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r348 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r349 4 87 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.31
r350 4 85 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.63
r351 3 73 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r352 3 71 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r353 2 91 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.42
r354 1 77 91 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.31 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBE_P_8%VPWR 1 2 3 4 5 6 21 23 27 29 33 35 39 41
+ 45 49 54 55 56 58 60 71 72 75 78 81 84 87
c111 45 0 1.22282e-19 $X=4.49 $Y=2
c112 4 0 1.8139e-19 $X=3.405 $Y=1.485
c113 3 0 1.8139e-19 $X=2.465 $Y=1.485
c114 2 0 1.8139e-19 $X=1.525 $Y=1.485
r115 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r116 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r117 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r118 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r119 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r120 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r121 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r123 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r125 69 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r126 69 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r127 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r128 66 87 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.49 $Y2=2.72
r129 66 68 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=5.29 $Y2=2.72
r130 60 75 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.73 $Y2=2.72
r131 58 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r132 56 60 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.595 $Y2=2.72
r133 56 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r134 54 68 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.295 $Y=2.72
+ $X2=5.29 $Y2=2.72
r135 54 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.295 $Y=2.72
+ $X2=5.445 $Y2=2.72
r136 53 71 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=5.75 $Y2=2.72
r137 53 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=5.445 $Y2=2.72
r138 49 52 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=5.445 $Y=1.66
+ $X2=5.445 $Y2=2.34
r139 47 55 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=2.635
+ $X2=5.445 $Y2=2.72
r140 47 52 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.445 $Y=2.635
+ $X2=5.445 $Y2=2.34
r141 43 87 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=2.635
+ $X2=4.49 $Y2=2.72
r142 43 45 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.49 $Y=2.635
+ $X2=4.49 $Y2=2
r143 42 84 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.55 $Y2=2.72
r144 41 87 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=2.72
+ $X2=4.49 $Y2=2.72
r145 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=2.72
+ $X2=3.685 $Y2=2.72
r146 37 84 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2.72
r147 37 39 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2
r148 36 81 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=2.61 $Y2=2.72
r149 35 84 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=3.55 $Y2=2.72
r150 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=2.745 $Y2=2.72
r151 31 81 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=2.72
r152 31 33 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=2
r153 30 78 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.67 $Y2=2.72
r154 29 81 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.475 $Y=2.72
+ $X2=2.61 $Y2=2.72
r155 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=2.72
+ $X2=1.805 $Y2=2.72
r156 25 78 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r157 25 27 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2
r158 24 75 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.73 $Y2=2.72
r159 23 78 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=1.67 $Y2=2.72
r160 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=0.865 $Y2=2.72
r161 19 75 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r162 19 21 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2
r163 6 52 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.34
r164 6 49 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.66
r165 5 45 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2
r166 4 39 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2
r167 3 33 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2
r168 2 27 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2
r169 1 21 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBE_P_8%A_399_297# 1 2 3 4 5 6 7 8 27 31 33 34
+ 35 36 39 43 45 47 51 55 59 63 65 66 67 69 72 74 75 78 80 84 88
c241 75 0 2.33346e-19 $X=3.56 $Y=1.27
c242 74 0 9.74311e-19 $X=3.56 $Y=1.27
c243 72 0 1.2638e-19 $X=3.975 $Y=1.19
r244 87 88 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=3.945 $Y=1.19
+ $X2=3.945 $Y2=1.19
r245 78 88 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=3.985 $Y=1.19
+ $X2=3.985 $Y2=1.19
r246 75 80 0.00650012 $w=3.02e-06 $l=6.75e-07 $layer=MET5_cond $X=2.76 $Y=1.27
+ $X2=2.76 $Y2=1.945
r247 74 78 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=3.985 $Y=1.19
+ $X2=3.985 $Y2=1.19
r248 74 75 0.19 $w=8e-07 $l=1.6e-06 $layer=via4_notcap2m $count=2 $X=3.56
+ $Y=1.27 $X2=3.56 $Y2=1.27
r249 72 87 0.0170272 $w=2.6e-07 $l=3e-08 $layer=MET1_cond $X=3.975 $Y=1.19
+ $X2=3.945 $Y2=1.19
r250 70 84 0.789928 $w=6.95e-07 $l=4.5e-08 $layer=LI1_cond $X=5.005 $Y=1.175
+ $X2=4.96 $Y2=1.175
r251 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.005 $Y=1.19
+ $X2=5.005 $Y2=1.19
r252 67 72 0.0749482 $w=2.6e-07 $l=1.3e-07 $layer=MET1_cond $X=4.105 $Y=1.19
+ $X2=3.975 $Y2=1.19
r253 67 69 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=4.105 $Y=1.19
+ $X2=5.005 $Y2=1.19
r254 61 84 5.10968 $w=3.3e-07 $l=4.4e-07 $layer=LI1_cond $X=4.96 $Y=1.615
+ $X2=4.96 $Y2=1.175
r255 61 63 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=4.96 $Y=1.615
+ $X2=4.96 $Y2=1.755
r256 57 84 5.10968 $w=3.3e-07 $l=4.4e-07 $layer=LI1_cond $X=4.96 $Y=0.735
+ $X2=4.96 $Y2=1.175
r257 57 59 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.96 $Y=0.735
+ $X2=4.96 $Y2=0.42
r258 53 55 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=4.02 $Y=1.615
+ $X2=4.02 $Y2=1.755
r259 49 84 16.5007 $w=6.95e-07 $l=1.13895e-06 $layer=LI1_cond $X=4.02 $Y=0.735
+ $X2=4.96 $Y2=1.175
r260 49 53 5.10968 $w=3.3e-07 $l=8.8e-07 $layer=LI1_cond $X=4.02 $Y=0.735
+ $X2=4.02 $Y2=1.615
r261 49 51 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.02 $Y=0.735
+ $X2=4.02 $Y2=0.42
r262 48 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=1.53
+ $X2=3.08 $Y2=1.53
r263 47 49 6.53734 $w=3.47e-07 $l=8.73613e-07 $layer=LI1_cond $X=3.855 $Y=1.53
+ $X2=4.02 $Y2=0.735
r264 47 48 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=1.53
+ $X2=3.245 $Y2=1.53
r265 46 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0.82
+ $X2=3.08 $Y2=0.82
r266 45 49 6.53734 $w=3.47e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.855 $Y=0.82
+ $X2=4.02 $Y2=0.735
r267 45 46 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=0.82
+ $X2=3.245 $Y2=0.82
r268 41 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=1.615
+ $X2=3.08 $Y2=1.53
r269 41 43 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.08 $Y=1.615
+ $X2=3.08 $Y2=1.755
r270 37 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.735
+ $X2=3.08 $Y2=0.82
r271 37 39 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.08 $Y=0.735
+ $X2=3.08 $Y2=0.42
r272 35 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=1.53
+ $X2=3.08 $Y2=1.53
r273 35 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=1.53
+ $X2=2.305 $Y2=1.53
r274 33 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0.82
+ $X2=3.08 $Y2=0.82
r275 33 34 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=0.82
+ $X2=2.305 $Y2=0.82
r276 29 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.14 $Y=1.615
+ $X2=2.305 $Y2=1.53
r277 29 31 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.14 $Y=1.615
+ $X2=2.14 $Y2=1.755
r278 25 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.305 $Y2=0.82
r279 25 27 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.14 $Y2=0.42
r280 8 63 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.755
r281 7 55 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.755
r282 6 43 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.755
r283 5 31 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.755
r284 4 59 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.235 $X2=4.96 $Y2=0.42
r285 3 51 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.42
r286 2 39 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.42
r287 1 27 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBE_P_8%VGND 1 2 3 4 5 6 21 25 27 31 33 37 39 43
+ 47 50 51 52 54 56 66 67 69 71 74 77 80 83 86 90
c120 43 0 2.9272e-20 $X=4.49 $Y=0.4
c121 21 0 1.28869e-20 $X=0.76 $Y=0.4
r122 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r123 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r124 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r125 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r126 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r127 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r128 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r129 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r130 69 71 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.755
+ $Y2=0
r131 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r132 64 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r133 64 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.37
+ $Y2=0
r134 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r135 61 83 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.49
+ $Y2=0
r136 61 63 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=5.29
+ $Y2=0
r137 60 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r138 60 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r139 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r140 57 71 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.755
+ $Y2=0
r141 57 59 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r142 56 74 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.505 $Y=0 $X2=1.655
+ $Y2=0
r143 56 59 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.505 $Y=0
+ $X2=1.15 $Y2=0
r144 54 72 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r145 54 90 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r146 52 69 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.235 $Y=0
+ $X2=0.615 $Y2=0
r147 52 86 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r148 50 63 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.29
+ $Y2=0
r149 50 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.42
+ $Y2=0
r150 49 66 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.545 $Y=0
+ $X2=5.75 $Y2=0
r151 49 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.545 $Y=0 $X2=5.42
+ $Y2=0
r152 45 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.42 $Y=0.085
+ $X2=5.42 $Y2=0
r153 45 47 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.42 $Y=0.085
+ $X2=5.42 $Y2=0.38
r154 41 83 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0
r155 41 43 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0.4
r156 40 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.55
+ $Y2=0
r157 39 83 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.49
+ $Y2=0
r158 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=0
+ $X2=3.685 $Y2=0
r159 35 80 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r160 35 37 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.4
r161 34 77 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.61
+ $Y2=0
r162 33 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.55
+ $Y2=0
r163 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=0
+ $X2=2.745 $Y2=0
r164 29 77 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r165 29 31 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.4
r166 28 74 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.655
+ $Y2=0
r167 27 77 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.61
+ $Y2=0
r168 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=1.805 $Y2=0
r169 23 74 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0
r170 23 25 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0.4
r171 19 71 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r172 19 21 12.965 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.4
r173 6 47 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.245
+ $Y=0.235 $X2=5.38 $Y2=0.38
r174 5 43 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.4
r175 4 37 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.4
r176 3 31 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.4
r177 2 25 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.4
r178 1 21 182 $w=1.7e-07 $l=2.33345e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.76 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBE_P_8%X 1 3
r20 1 3 0.00103039 $w=3.02e-06 $l=1.07e-07 $layer=MET5_cond $X=2.76 $Y=2.057
+ $X2=2.76 $Y2=1.95
.ends

