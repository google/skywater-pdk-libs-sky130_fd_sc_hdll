* NGSPICE file created from sky130_fd_sc_hdll__o2bb2ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_121_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=1.96e+12p ps=1.392e+07u
M1001 a_121_297# A2_N a_123_47# VNB nshort w=650000u l=150000u
+  ad=2.405e+11p pd=2.04e+06u as=3.575e+11p ps=3.7e+06u
M1002 a_503_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=8.7425e+11p pd=7.89e+06u as=7.345e+11p ps=7.46e+06u
M1003 VPWR A1_N a_121_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A1_N a_123_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_788_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=5.8e+11p ps=5.16e+06u
M1006 a_123_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_121_297# A2_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B2 a_788_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_121_297# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_503_47# a_121_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1011 a_123_47# A2_N a_121_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_121_297# a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_503_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_788_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A2_N a_121_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_121_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B2 a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND B1 a_503_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR B1 a_788_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

