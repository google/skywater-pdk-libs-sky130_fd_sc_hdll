* File: sky130_fd_sc_hdll__a211o_4.pxi.spice
* Created: Wed Sep  2 08:15:55 2020
* 
x_PM_SKY130_FD_SC_HDLL__A211O_4%A_79_204# N_A_79_204#_M1007_d
+ N_A_79_204#_M1023_d N_A_79_204#_M1016_s N_A_79_204#_M1006_s
+ N_A_79_204#_c_100_n N_A_79_204#_M1003_g N_A_79_204#_M1001_g
+ N_A_79_204#_c_101_n N_A_79_204#_M1009_g N_A_79_204#_M1004_g
+ N_A_79_204#_c_102_n N_A_79_204#_M1010_g N_A_79_204#_M1005_g
+ N_A_79_204#_c_103_n N_A_79_204#_M1020_g N_A_79_204#_M1011_g
+ N_A_79_204#_c_161_p N_A_79_204#_c_97_n N_A_79_204#_c_104_n N_A_79_204#_c_111_p
+ N_A_79_204#_c_189_p N_A_79_204#_c_105_n N_A_79_204#_c_114_p
+ N_A_79_204#_c_215_p N_A_79_204#_c_136_p N_A_79_204#_c_122_p N_A_79_204#_c_98_n
+ N_A_79_204#_c_106_n N_A_79_204#_c_107_n N_A_79_204#_c_118_p
+ N_A_79_204#_c_121_p N_A_79_204#_c_144_p N_A_79_204#_c_99_n
+ PM_SKY130_FD_SC_HDLL__A211O_4%A_79_204#
x_PM_SKY130_FD_SC_HDLL__A211O_4%B1 N_B1_M1007_g N_B1_c_253_n N_B1_M1017_g
+ N_B1_c_254_n N_B1_M1015_g N_B1_c_255_n N_B1_M1013_g N_B1_c_260_n B1
+ N_B1_c_256_n B1 N_B1_c_257_n PM_SKY130_FD_SC_HDLL__A211O_4%B1
x_PM_SKY130_FD_SC_HDLL__A211O_4%C1 N_C1_c_341_n N_C1_M1012_g N_C1_c_345_n
+ N_C1_M1006_g N_C1_c_346_n N_C1_M1022_g N_C1_c_342_n N_C1_M1023_g C1
+ N_C1_c_344_n C1 PM_SKY130_FD_SC_HDLL__A211O_4%C1
x_PM_SKY130_FD_SC_HDLL__A211O_4%A2 N_A2_c_387_n N_A2_M1000_g N_A2_M1002_g
+ N_A2_c_389_n N_A2_M1019_g N_A2_c_390_n N_A2_M1021_g N_A2_c_391_n N_A2_c_392_n
+ N_A2_c_393_n N_A2_c_428_p A2 N_A2_c_416_p A2 PM_SKY130_FD_SC_HDLL__A211O_4%A2
x_PM_SKY130_FD_SC_HDLL__A211O_4%A1 N_A1_M1016_g N_A1_c_463_n N_A1_M1008_g
+ N_A1_c_464_n N_A1_M1018_g N_A1_M1014_g A1 N_A1_c_462_n A1
+ PM_SKY130_FD_SC_HDLL__A211O_4%A1
x_PM_SKY130_FD_SC_HDLL__A211O_4%VPWR N_VPWR_M1003_d N_VPWR_M1009_d
+ N_VPWR_M1020_d N_VPWR_M1000_d N_VPWR_M1018_d N_VPWR_c_506_n N_VPWR_c_507_n
+ N_VPWR_c_508_n N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n VPWR
+ N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n N_VPWR_c_505_n N_VPWR_c_516_n
+ N_VPWR_c_517_n N_VPWR_c_518_n N_VPWR_c_519_n
+ PM_SKY130_FD_SC_HDLL__A211O_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A211O_4%X N_X_M1001_d N_X_M1005_d N_X_M1003_s
+ N_X_M1010_s N_X_c_612_n N_X_c_620_n N_X_c_615_n N_X_c_622_n N_X_c_623_n
+ N_X_c_662_p N_X_c_627_n N_X_c_655_n N_X_c_634_n N_X_c_635_n N_X_c_637_n X
+ N_X_c_614_n PM_SKY130_FD_SC_HDLL__A211O_4%X
x_PM_SKY130_FD_SC_HDLL__A211O_4%A_523_297# N_A_523_297#_M1017_d
+ N_A_523_297#_M1015_d N_A_523_297#_M1008_s N_A_523_297#_M1021_s
+ N_A_523_297#_c_677_n N_A_523_297#_c_696_n N_A_523_297#_c_699_n
+ N_A_523_297#_c_700_n N_A_523_297#_c_678_n N_A_523_297#_c_692_n
+ N_A_523_297#_c_704_n N_A_523_297#_c_679_n
+ PM_SKY130_FD_SC_HDLL__A211O_4%A_523_297#
x_PM_SKY130_FD_SC_HDLL__A211O_4%VGND N_VGND_M1001_s N_VGND_M1004_s
+ N_VGND_M1011_s N_VGND_M1012_s N_VGND_M1013_s N_VGND_M1019_d N_VGND_c_749_n
+ N_VGND_c_750_n VGND N_VGND_c_751_n N_VGND_c_752_n N_VGND_c_753_n
+ N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n N_VGND_c_758_n
+ N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n
+ PM_SKY130_FD_SC_HDLL__A211O_4%VGND
cc_1 VNB N_A_79_204#_M1001_g 0.0212264f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=0.56
cc_2 VNB N_A_79_204#_M1004_g 0.0183243f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.56
cc_3 VNB N_A_79_204#_M1005_g 0.0189261f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=0.56
cc_4 VNB N_A_79_204#_M1011_g 0.0181311f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.56
cc_5 VNB N_A_79_204#_c_97_n 0.00137203f $X=-0.19 $Y=-0.24 $X2=2.507 $Y2=1.045
cc_6 VNB N_A_79_204#_c_98_n 0.00154767f $X=-0.19 $Y=-0.24 $X2=2.502 $Y2=1.185
cc_7 VNB N_A_79_204#_c_99_n 0.0976531f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=1.215
cc_8 VNB N_B1_M1007_g 0.0185426f $X=-0.19 $Y=-0.24 $X2=5.685 $Y2=0.235
cc_9 VNB N_B1_c_253_n 0.0254542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B1_c_254_n 0.0316648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B1_c_255_n 0.0189254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B1_c_256_n 0.0038905f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_13 VNB N_B1_c_257_n 0.00218192f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.985
cc_14 VNB N_C1_c_341_n 0.0175738f $X=-0.19 $Y=-0.24 $X2=2.98 $Y2=0.235
cc_15 VNB N_C1_c_342_n 0.0186224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB C1 0.00858011f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_17 VNB N_C1_c_344_n 0.0388186f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.41
cc_18 VNB N_A2_c_387_n 0.0287331f $X=-0.19 $Y=-0.24 $X2=2.98 $Y2=0.235
cc_19 VNB N_A2_M1002_g 0.019793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_389_n 0.0226581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A2_c_390_n 0.0303585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A2_c_391_n 0.00232883f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=1.02
cc_23 VNB N_A2_c_392_n 0.00936732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A2_c_393_n 0.0133716f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_25 VNB N_A1_M1016_g 0.0187667f $X=-0.19 $Y=-0.24 $X2=5.685 $Y2=0.235
cc_26 VNB N_A1_M1014_g 0.0187667f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_27 VNB A1 0.00188191f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_28 VNB N_A1_c_462_n 0.0322087f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_29 VNB N_VPWR_c_505_n 0.30769f $X=-0.19 $Y=-0.24 $X2=2.502 $Y2=1.505
cc_30 VNB N_X_c_612_n 0.00564768f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_31 VNB X 0.0232413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_614_n 0.0154224f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.16
cc_33 VNB N_VGND_c_749_n 0.0150396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_750_n 0.0269949f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.02
cc_35 VNB N_VGND_c_751_n 0.0158235f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_36 VNB N_VGND_c_752_n 0.0127938f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=0.56
cc_37 VNB N_VGND_c_753_n 0.0221152f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=1.02
cc_38 VNB N_VGND_c_754_n 0.0204782f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.185
cc_39 VNB N_VGND_c_755_n 0.0435581f $X=-0.19 $Y=-0.24 $X2=1.91 $Y2=1.16
cc_40 VNB N_VGND_c_756_n 0.0137583f $X=-0.19 $Y=-0.24 $X2=2.617 $Y2=1.87
cc_41 VNB N_VGND_c_757_n 0.367062f $X=-0.19 $Y=-0.24 $X2=3.025 $Y2=0.71
cc_42 VNB N_VGND_c_758_n 0.0183666f $X=-0.19 $Y=-0.24 $X2=3.695 $Y2=1.955
cc_43 VNB N_VGND_c_759_n 0.00538742f $X=-0.19 $Y=-0.24 $X2=3.27 $Y2=0.71
cc_44 VNB N_VGND_c_760_n 0.0093268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_761_n 0.0129872f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.215
cc_46 VNB N_VGND_c_762_n 0.00606646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VPB N_A_79_204#_c_100_n 0.0183848f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_48 VPB N_A_79_204#_c_101_n 0.016282f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_49 VPB N_A_79_204#_c_102_n 0.0162845f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_50 VPB N_A_79_204#_c_103_n 0.018725f $X=-0.19 $Y=1.305 $X2=1.935 $Y2=1.41
cc_51 VPB N_A_79_204#_c_104_n 0.00294181f $X=-0.19 $Y=1.305 $X2=2.617 $Y2=1.87
cc_52 VPB N_A_79_204#_c_105_n 0.00294396f $X=-0.19 $Y=1.305 $X2=2.705 $Y2=1.955
cc_53 VPB N_A_79_204#_c_106_n 0.00292389f $X=-0.19 $Y=1.305 $X2=2.545 $Y2=1.505
cc_54 VPB N_A_79_204#_c_107_n 0.00891413f $X=-0.19 $Y=1.305 $X2=2.545 $Y2=1.675
cc_55 VPB N_A_79_204#_c_99_n 0.0669462f $X=-0.19 $Y=1.305 $X2=1.935 $Y2=1.215
cc_56 VPB N_B1_c_253_n 0.0324643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_B1_c_254_n 0.0292766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_B1_c_260_n 0.00856966f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_59 VPB N_B1_c_256_n 0.00291569f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_60 VPB B1 3.33201e-19 $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.02
cc_61 VPB N_B1_c_257_n 0.00180084f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_62 VPB N_C1_c_345_n 0.016139f $X=-0.19 $Y=1.305 $X2=3.545 $Y2=1.485
cc_63 VPB N_C1_c_346_n 0.016433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_C1_c_344_n 0.0210835f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_65 VPB N_A2_c_387_n 0.0307308f $X=-0.19 $Y=1.305 $X2=2.98 $Y2=0.235
cc_66 VPB N_A2_c_390_n 0.036005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A2_c_391_n 0.00156915f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.02
cc_68 VPB N_A2_c_393_n 0.00133134f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_69 VPB A2 0.00160963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A1_c_463_n 0.0173408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A1_c_464_n 0.0156833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A1_c_462_n 0.0188511f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_73 VPB N_VPWR_c_506_n 0.0102036f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.02
cc_74 VPB N_VPWR_c_507_n 0.0268854f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=0.56
cc_75 VPB N_VPWR_c_508_n 3.41097e-19 $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_76 VPB N_VPWR_c_509_n 0.016122f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=0.56
cc_77 VPB N_VPWR_c_510_n 0.00238224f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_78 VPB N_VPWR_c_511_n 0.0160838f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.02
cc_79 VPB N_VPWR_c_512_n 0.0160099f $X=-0.19 $Y=1.305 $X2=1.935 $Y2=1.41
cc_80 VPB N_VPWR_c_513_n 0.0648995f $X=-0.19 $Y=1.305 $X2=2.42 $Y2=0.56
cc_81 VPB N_VPWR_c_514_n 0.0244336f $X=-0.19 $Y=1.305 $X2=2.502 $Y2=1.325
cc_82 VPB N_VPWR_c_505_n 0.0658879f $X=-0.19 $Y=1.305 $X2=2.502 $Y2=1.505
cc_83 VPB N_VPWR_c_516_n 0.00436868f $X=-0.19 $Y=1.305 $X2=2.62 $Y2=0.71
cc_84 VPB N_VPWR_c_517_n 0.00362881f $X=-0.19 $Y=1.305 $X2=3.695 $Y2=1.955
cc_85 VPB N_VPWR_c_518_n 0.00877707f $X=-0.19 $Y=1.305 $X2=3.147 $Y2=0.485
cc_86 VPB N_VPWR_c_519_n 0.00556536f $X=-0.19 $Y=1.305 $X2=2.502 $Y2=1.185
cc_87 VPB N_X_c_615_n 0.00955713f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.02
cc_88 VPB X 0.00946501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_523_297#_c_677_n 0.0035016f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_90 VPB N_A_523_297#_c_678_n 0.013765f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_91 VPB N_A_523_297#_c_679_n 0.0240238f $X=-0.19 $Y=1.305 $X2=2.42 $Y2=1.02
cc_92 N_A_79_204#_M1011_g N_B1_M1007_g 0.0208137f $X=2.42 $Y=0.56 $X2=0 $Y2=0
cc_93 N_A_79_204#_c_97_n N_B1_M1007_g 0.00393239f $X=2.507 $Y=1.045 $X2=0 $Y2=0
cc_94 N_A_79_204#_c_111_p N_B1_M1007_g 0.012235f $X=3.025 $Y=0.71 $X2=0 $Y2=0
cc_95 N_A_79_204#_c_104_n N_B1_c_253_n 0.00588072f $X=2.617 $Y=1.87 $X2=0 $Y2=0
cc_96 N_A_79_204#_c_111_p N_B1_c_253_n 0.00260941f $X=3.025 $Y=0.71 $X2=0 $Y2=0
cc_97 N_A_79_204#_c_114_p N_B1_c_253_n 0.0168669f $X=3.695 $Y=1.955 $X2=0 $Y2=0
cc_98 N_A_79_204#_c_98_n N_B1_c_253_n 0.00207022f $X=2.502 $Y=1.185 $X2=0 $Y2=0
cc_99 N_A_79_204#_c_106_n N_B1_c_253_n 0.00121451f $X=2.545 $Y=1.505 $X2=0 $Y2=0
cc_100 N_A_79_204#_c_107_n N_B1_c_253_n 0.00140414f $X=2.545 $Y=1.675 $X2=0
+ $Y2=0
cc_101 N_A_79_204#_c_118_p N_B1_c_253_n 4.17806e-19 $X=3.147 $Y=0.71 $X2=0 $Y2=0
cc_102 N_A_79_204#_c_99_n N_B1_c_253_n 0.0201105f $X=1.935 $Y=1.215 $X2=0 $Y2=0
cc_103 N_A_79_204#_c_114_p N_B1_c_254_n 7.5355e-19 $X=3.695 $Y=1.955 $X2=0 $Y2=0
cc_104 N_A_79_204#_c_121_p N_B1_c_254_n 0.00131729f $X=4.235 $Y=0.38 $X2=0 $Y2=0
cc_105 N_A_79_204#_c_122_p N_B1_c_255_n 0.0128213f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_106 N_A_79_204#_M1006_s N_B1_c_260_n 0.00200696f $X=3.545 $Y=1.485 $X2=0
+ $Y2=0
cc_107 N_A_79_204#_c_114_p N_B1_c_260_n 0.0414396f $X=3.695 $Y=1.955 $X2=0 $Y2=0
cc_108 N_A_79_204#_c_118_p N_B1_c_260_n 0.00482114f $X=3.147 $Y=0.71 $X2=0 $Y2=0
cc_109 N_A_79_204#_c_121_p N_B1_c_260_n 0.00561844f $X=4.235 $Y=0.38 $X2=0 $Y2=0
cc_110 N_A_79_204#_c_97_n N_B1_c_256_n 0.0047176f $X=2.507 $Y=1.045 $X2=0 $Y2=0
cc_111 N_A_79_204#_c_111_p N_B1_c_256_n 0.0144926f $X=3.025 $Y=0.71 $X2=0 $Y2=0
cc_112 N_A_79_204#_c_114_p N_B1_c_256_n 0.0155858f $X=3.695 $Y=1.955 $X2=0 $Y2=0
cc_113 N_A_79_204#_c_98_n N_B1_c_256_n 0.023651f $X=2.502 $Y=1.185 $X2=0 $Y2=0
cc_114 N_A_79_204#_c_106_n N_B1_c_256_n 0.00989635f $X=2.545 $Y=1.505 $X2=0
+ $Y2=0
cc_115 N_A_79_204#_c_118_p N_B1_c_256_n 0.00647074f $X=3.147 $Y=0.71 $X2=0 $Y2=0
cc_116 N_A_79_204#_c_99_n N_B1_c_256_n 2.87201e-19 $X=1.935 $Y=1.215 $X2=0 $Y2=0
cc_117 N_A_79_204#_c_122_p N_B1_c_257_n 0.0131976f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_118 N_A_79_204#_c_121_p N_B1_c_257_n 0.014241f $X=4.235 $Y=0.38 $X2=0 $Y2=0
cc_119 N_A_79_204#_c_136_p N_C1_c_341_n 0.0126456f $X=4.04 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A_79_204#_c_114_p N_C1_c_345_n 0.00979272f $X=3.695 $Y=1.955 $X2=0
+ $Y2=0
cc_121 N_A_79_204#_c_114_p N_C1_c_346_n 0.00385452f $X=3.695 $Y=1.955 $X2=0
+ $Y2=0
cc_122 N_A_79_204#_c_136_p N_C1_c_342_n 0.0124091f $X=4.04 $Y=0.71 $X2=0 $Y2=0
cc_123 N_A_79_204#_c_136_p C1 0.0500168f $X=4.04 $Y=0.71 $X2=0 $Y2=0
cc_124 N_A_79_204#_c_136_p N_C1_c_344_n 0.00176462f $X=4.04 $Y=0.71 $X2=0 $Y2=0
cc_125 N_A_79_204#_c_122_p N_A2_c_387_n 0.00124013f $X=5.66 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_126 N_A_79_204#_c_122_p N_A2_M1002_g 0.0137471f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_127 N_A_79_204#_c_144_p N_A2_M1002_g 0.00144205f $X=5.875 $Y=0.36 $X2=0 $Y2=0
cc_128 N_A_79_204#_c_122_p N_A2_c_391_n 0.0210355f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_129 N_A_79_204#_c_122_p N_A1_M1016_g 0.0102493f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_130 N_A_79_204#_c_144_p N_A1_M1016_g 0.00801394f $X=5.875 $Y=0.36 $X2=0 $Y2=0
cc_131 N_A_79_204#_c_122_p A1 0.00742174f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_132 N_A_79_204#_c_144_p A1 0.0159169f $X=5.875 $Y=0.36 $X2=0 $Y2=0
cc_133 N_A_79_204#_c_144_p N_A1_c_462_n 0.00532608f $X=5.875 $Y=0.36 $X2=0 $Y2=0
cc_134 N_A_79_204#_c_100_n N_VPWR_c_507_n 0.012418f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_79_204#_c_101_n N_VPWR_c_507_n 6.20014e-19 $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_136 N_A_79_204#_c_100_n N_VPWR_c_508_n 6.12193e-19 $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_137 N_A_79_204#_c_101_n N_VPWR_c_508_n 0.0110019f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_A_79_204#_c_102_n N_VPWR_c_508_n 0.0110118f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_79_204#_c_103_n N_VPWR_c_508_n 6.13845e-19 $X=1.935 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_79_204#_c_102_n N_VPWR_c_509_n 0.00642146f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_79_204#_c_103_n N_VPWR_c_509_n 0.00642146f $X=1.935 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_79_204#_c_102_n N_VPWR_c_510_n 6.21524e-19 $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_143 N_A_79_204#_c_103_n N_VPWR_c_510_n 0.0124444f $X=1.935 $Y=1.41 $X2=0
+ $Y2=0
cc_144 N_A_79_204#_c_161_p N_VPWR_c_510_n 0.00743697f $X=2.385 $Y=1.185 $X2=0
+ $Y2=0
cc_145 N_A_79_204#_c_104_n N_VPWR_c_510_n 0.00189014f $X=2.617 $Y=1.87 $X2=0
+ $Y2=0
cc_146 N_A_79_204#_c_105_n N_VPWR_c_510_n 0.0104061f $X=2.705 $Y=1.955 $X2=0
+ $Y2=0
cc_147 N_A_79_204#_c_99_n N_VPWR_c_510_n 0.00409787f $X=1.935 $Y=1.215 $X2=0
+ $Y2=0
cc_148 N_A_79_204#_c_100_n N_VPWR_c_512_n 0.00622633f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_149 N_A_79_204#_c_101_n N_VPWR_c_512_n 0.00642146f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_150 N_A_79_204#_c_105_n N_VPWR_c_513_n 7.41891e-19 $X=2.705 $Y=1.955 $X2=0
+ $Y2=0
cc_151 N_A_79_204#_M1006_s N_VPWR_c_505_n 0.00240926f $X=3.545 $Y=1.485 $X2=0
+ $Y2=0
cc_152 N_A_79_204#_c_100_n N_VPWR_c_505_n 0.0104265f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_153 N_A_79_204#_c_101_n N_VPWR_c_505_n 0.0107337f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_154 N_A_79_204#_c_102_n N_VPWR_c_505_n 0.0107337f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_155 N_A_79_204#_c_103_n N_VPWR_c_505_n 0.0107337f $X=1.935 $Y=1.41 $X2=0
+ $Y2=0
cc_156 N_A_79_204#_c_105_n N_VPWR_c_505_n 0.0014742f $X=2.705 $Y=1.955 $X2=0
+ $Y2=0
cc_157 N_A_79_204#_M1001_g N_X_c_612_n 0.0176196f $X=0.915 $Y=0.56 $X2=0 $Y2=0
cc_158 N_A_79_204#_c_161_p N_X_c_612_n 0.0371314f $X=2.385 $Y=1.185 $X2=0 $Y2=0
cc_159 N_A_79_204#_c_99_n N_X_c_612_n 0.0117397f $X=1.935 $Y=1.215 $X2=0 $Y2=0
cc_160 N_A_79_204#_c_100_n N_X_c_620_n 0.021161f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_79_204#_c_161_p N_X_c_620_n 0.00649136f $X=2.385 $Y=1.185 $X2=0 $Y2=0
cc_162 N_A_79_204#_c_100_n N_X_c_622_n 0.0057123f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_79_204#_c_101_n N_X_c_623_n 0.0183884f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_79_204#_c_102_n N_X_c_623_n 0.0179391f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_79_204#_c_161_p N_X_c_623_n 0.0630823f $X=2.385 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A_79_204#_c_99_n N_X_c_623_n 0.0116685f $X=1.935 $Y=1.215 $X2=0 $Y2=0
cc_167 N_A_79_204#_M1004_g N_X_c_627_n 0.0158375f $X=1.395 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A_79_204#_M1005_g N_X_c_627_n 0.0155667f $X=1.875 $Y=0.56 $X2=0 $Y2=0
cc_169 N_A_79_204#_M1011_g N_X_c_627_n 0.00216789f $X=2.42 $Y=0.56 $X2=0 $Y2=0
cc_170 N_A_79_204#_c_161_p N_X_c_627_n 0.0634055f $X=2.385 $Y=1.185 $X2=0 $Y2=0
cc_171 N_A_79_204#_c_97_n N_X_c_627_n 0.00559455f $X=2.507 $Y=1.045 $X2=0 $Y2=0
cc_172 N_A_79_204#_c_189_p N_X_c_627_n 0.0166067f $X=2.62 $Y=0.71 $X2=0 $Y2=0
cc_173 N_A_79_204#_c_99_n N_X_c_627_n 0.00791525f $X=1.935 $Y=1.215 $X2=0 $Y2=0
cc_174 N_A_79_204#_M1011_g N_X_c_634_n 0.00545406f $X=2.42 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_79_204#_c_161_p N_X_c_635_n 0.0150142f $X=2.385 $Y=1.185 $X2=0 $Y2=0
cc_176 N_A_79_204#_c_99_n N_X_c_635_n 0.0044351f $X=1.935 $Y=1.215 $X2=0 $Y2=0
cc_177 N_A_79_204#_M1001_g N_X_c_637_n 6.14708e-19 $X=0.915 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A_79_204#_c_161_p N_X_c_637_n 0.0148656f $X=2.385 $Y=1.185 $X2=0 $Y2=0
cc_179 N_A_79_204#_c_99_n N_X_c_637_n 0.00346571f $X=1.935 $Y=1.215 $X2=0 $Y2=0
cc_180 N_A_79_204#_c_100_n X 0.00345199f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_79_204#_M1001_g X 0.00366097f $X=0.915 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A_79_204#_c_161_p X 0.021458f $X=2.385 $Y=1.185 $X2=0 $Y2=0
cc_183 N_A_79_204#_c_99_n X 0.0135966f $X=1.935 $Y=1.215 $X2=0 $Y2=0
cc_184 N_A_79_204#_c_104_n N_A_523_297#_M1017_d 0.00312401f $X=2.617 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_185 N_A_79_204#_c_105_n N_A_523_297#_M1017_d 0.00174358f $X=2.705 $Y=1.955
+ $X2=-0.19 $Y2=-0.24
cc_186 N_A_79_204#_c_114_p N_A_523_297#_M1017_d 0.0031205f $X=3.695 $Y=1.955
+ $X2=-0.19 $Y2=-0.24
cc_187 N_A_79_204#_c_107_n N_A_523_297#_M1017_d 0.00584656f $X=2.545 $Y=1.675
+ $X2=-0.19 $Y2=-0.24
cc_188 N_A_79_204#_M1006_s N_A_523_297#_c_677_n 0.00377586f $X=3.545 $Y=1.485
+ $X2=0 $Y2=0
cc_189 N_A_79_204#_c_105_n N_A_523_297#_c_677_n 0.0107845f $X=2.705 $Y=1.955
+ $X2=0 $Y2=0
cc_190 N_A_79_204#_c_114_p N_A_523_297#_c_677_n 0.0604959f $X=3.695 $Y=1.955
+ $X2=0 $Y2=0
cc_191 N_A_79_204#_c_114_p A_613_297# 0.00389435f $X=3.695 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_192 N_A_79_204#_c_97_n N_VGND_M1011_s 9.75292e-19 $X=2.507 $Y=1.045 $X2=0
+ $Y2=0
cc_193 N_A_79_204#_c_111_p N_VGND_M1011_s 0.00576059f $X=3.025 $Y=0.71 $X2=0
+ $Y2=0
cc_194 N_A_79_204#_c_189_p N_VGND_M1011_s 7.2107e-19 $X=2.62 $Y=0.71 $X2=0 $Y2=0
cc_195 N_A_79_204#_c_136_p N_VGND_M1012_s 0.00702892f $X=4.04 $Y=0.71 $X2=0
+ $Y2=0
cc_196 N_A_79_204#_c_122_p N_VGND_M1013_s 0.0164032f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_197 N_A_79_204#_c_111_p N_VGND_c_749_n 0.00330545f $X=3.025 $Y=0.71 $X2=0
+ $Y2=0
cc_198 N_A_79_204#_c_215_p N_VGND_c_749_n 0.0155765f $X=3.12 $Y=0.485 $X2=0
+ $Y2=0
cc_199 N_A_79_204#_c_136_p N_VGND_c_749_n 0.00272015f $X=4.04 $Y=0.71 $X2=0
+ $Y2=0
cc_200 N_A_79_204#_M1001_g N_VGND_c_752_n 0.00354245f $X=0.915 $Y=0.56 $X2=0
+ $Y2=0
cc_201 N_A_79_204#_M1004_g N_VGND_c_752_n 0.0035176f $X=1.395 $Y=0.56 $X2=0
+ $Y2=0
cc_202 N_A_79_204#_M1005_g N_VGND_c_753_n 0.00403223f $X=1.875 $Y=0.56 $X2=0
+ $Y2=0
cc_203 N_A_79_204#_M1011_g N_VGND_c_753_n 0.0119817f $X=2.42 $Y=0.56 $X2=0 $Y2=0
cc_204 N_A_79_204#_c_111_p N_VGND_c_753_n 0.0116493f $X=3.025 $Y=0.71 $X2=0
+ $Y2=0
cc_205 N_A_79_204#_c_189_p N_VGND_c_753_n 0.0119372f $X=2.62 $Y=0.71 $X2=0 $Y2=0
cc_206 N_A_79_204#_c_136_p N_VGND_c_754_n 0.00337739f $X=4.04 $Y=0.71 $X2=0
+ $Y2=0
cc_207 N_A_79_204#_c_122_p N_VGND_c_754_n 0.0033124f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_208 N_A_79_204#_c_121_p N_VGND_c_754_n 0.0244177f $X=4.235 $Y=0.38 $X2=0
+ $Y2=0
cc_209 N_A_79_204#_c_122_p N_VGND_c_755_n 0.0102742f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_210 N_A_79_204#_c_144_p N_VGND_c_755_n 0.020466f $X=5.875 $Y=0.36 $X2=0 $Y2=0
cc_211 N_A_79_204#_M1007_d N_VGND_c_757_n 0.00280564f $X=2.98 $Y=0.235 $X2=0
+ $Y2=0
cc_212 N_A_79_204#_M1023_d N_VGND_c_757_n 0.00373225f $X=4.035 $Y=0.235 $X2=0
+ $Y2=0
cc_213 N_A_79_204#_M1016_s N_VGND_c_757_n 0.00391417f $X=5.685 $Y=0.235 $X2=0
+ $Y2=0
cc_214 N_A_79_204#_M1001_g N_VGND_c_757_n 0.00423769f $X=0.915 $Y=0.56 $X2=0
+ $Y2=0
cc_215 N_A_79_204#_M1004_g N_VGND_c_757_n 0.0041977f $X=1.395 $Y=0.56 $X2=0
+ $Y2=0
cc_216 N_A_79_204#_M1005_g N_VGND_c_757_n 0.00434273f $X=1.875 $Y=0.56 $X2=0
+ $Y2=0
cc_217 N_A_79_204#_M1011_g N_VGND_c_757_n 0.00470696f $X=2.42 $Y=0.56 $X2=0
+ $Y2=0
cc_218 N_A_79_204#_c_111_p N_VGND_c_757_n 0.00639818f $X=3.025 $Y=0.71 $X2=0
+ $Y2=0
cc_219 N_A_79_204#_c_189_p N_VGND_c_757_n 0.00168439f $X=2.62 $Y=0.71 $X2=0
+ $Y2=0
cc_220 N_A_79_204#_c_215_p N_VGND_c_757_n 0.00930702f $X=3.12 $Y=0.485 $X2=0
+ $Y2=0
cc_221 N_A_79_204#_c_136_p N_VGND_c_757_n 0.0116351f $X=4.04 $Y=0.71 $X2=0 $Y2=0
cc_222 N_A_79_204#_c_122_p N_VGND_c_757_n 0.0247205f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_223 N_A_79_204#_c_121_p N_VGND_c_757_n 0.0144726f $X=4.235 $Y=0.38 $X2=0
+ $Y2=0
cc_224 N_A_79_204#_c_144_p N_VGND_c_757_n 0.0141362f $X=5.875 $Y=0.36 $X2=0
+ $Y2=0
cc_225 N_A_79_204#_M1001_g N_VGND_c_758_n 0.00799521f $X=0.915 $Y=0.56 $X2=0
+ $Y2=0
cc_226 N_A_79_204#_M1004_g N_VGND_c_758_n 5.06948e-19 $X=1.395 $Y=0.56 $X2=0
+ $Y2=0
cc_227 N_A_79_204#_M1001_g N_VGND_c_759_n 4.87918e-19 $X=0.915 $Y=0.56 $X2=0
+ $Y2=0
cc_228 N_A_79_204#_M1004_g N_VGND_c_759_n 0.00661042f $X=1.395 $Y=0.56 $X2=0
+ $Y2=0
cc_229 N_A_79_204#_M1005_g N_VGND_c_759_n 0.00689291f $X=1.875 $Y=0.56 $X2=0
+ $Y2=0
cc_230 N_A_79_204#_M1011_g N_VGND_c_759_n 5.05329e-19 $X=2.42 $Y=0.56 $X2=0
+ $Y2=0
cc_231 N_A_79_204#_c_136_p N_VGND_c_760_n 0.0244662f $X=4.04 $Y=0.71 $X2=0 $Y2=0
cc_232 N_A_79_204#_c_122_p N_VGND_c_761_n 0.0249683f $X=5.66 $Y=0.71 $X2=0 $Y2=0
cc_233 N_A_79_204#_c_144_p N_VGND_c_761_n 0.00463312f $X=5.875 $Y=0.36 $X2=0
+ $Y2=0
cc_234 N_A_79_204#_c_122_p A_1051_47# 0.00890637f $X=5.66 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_235 N_B1_M1007_g N_C1_c_341_n 0.0209223f $X=2.905 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_236 N_B1_c_256_n N_C1_c_341_n 8.86756e-19 $X=2.875 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_237 N_B1_c_253_n N_C1_c_345_n 0.0525852f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_238 N_B1_c_260_n N_C1_c_345_n 0.015641f $X=4.245 $Y=1.572 $X2=0 $Y2=0
cc_239 N_B1_c_256_n N_C1_c_345_n 6.98846e-19 $X=2.875 $Y=1.16 $X2=0 $Y2=0
cc_240 N_B1_c_254_n N_C1_c_346_n 0.0450471f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_241 N_B1_c_260_n N_C1_c_346_n 0.0178727f $X=4.245 $Y=1.572 $X2=0 $Y2=0
cc_242 N_B1_c_257_n N_C1_c_346_n 7.9991e-19 $X=4.41 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B1_c_254_n N_C1_c_342_n 0.0238768f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B1_c_255_n N_C1_c_342_n 0.0213053f $X=4.55 $Y=0.985 $X2=0 $Y2=0
cc_245 N_B1_c_257_n N_C1_c_342_n 3.511e-19 $X=4.41 $Y=1.16 $X2=0 $Y2=0
cc_246 N_B1_c_253_n C1 9.2392e-19 $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_247 N_B1_c_254_n C1 0.00182635f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B1_c_260_n C1 0.0578594f $X=4.245 $Y=1.572 $X2=0 $Y2=0
cc_249 N_B1_c_256_n C1 0.0255017f $X=2.875 $Y=1.16 $X2=0 $Y2=0
cc_250 N_B1_c_257_n C1 0.0217072f $X=4.41 $Y=1.16 $X2=0 $Y2=0
cc_251 N_B1_c_253_n N_C1_c_344_n 0.0242415f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B1_c_254_n N_C1_c_344_n 0.00210977f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B1_c_260_n N_C1_c_344_n 0.0100882f $X=4.245 $Y=1.572 $X2=0 $Y2=0
cc_254 N_B1_c_256_n N_C1_c_344_n 0.00293437f $X=2.875 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B1_c_257_n N_C1_c_344_n 0.00201166f $X=4.41 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B1_c_254_n N_A2_c_387_n 0.0381869f $X=4.455 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_257 B1 N_A2_c_387_n 0.00122212f $X=4.29 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_258 N_B1_c_257_n N_A2_c_387_n 0.0019696f $X=4.41 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_259 N_B1_c_255_n N_A2_M1002_g 0.0184281f $X=4.55 $Y=0.985 $X2=0 $Y2=0
cc_260 N_B1_c_254_n N_A2_c_391_n 0.00173038f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_261 B1 N_A2_c_391_n 0.00297653f $X=4.29 $Y=1.445 $X2=0 $Y2=0
cc_262 N_B1_c_257_n N_A2_c_391_n 0.0201759f $X=4.41 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B1_c_253_n N_VPWR_c_510_n 0.00570733f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B1_c_253_n N_VPWR_c_513_n 0.00429453f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B1_c_254_n N_VPWR_c_513_n 0.00429453f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B1_c_253_n N_VPWR_c_505_n 0.00739813f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B1_c_254_n N_VPWR_c_505_n 0.00649284f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_268 N_B1_c_254_n N_VPWR_c_518_n 9.27798e-19 $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_269 B1 N_A_523_297#_M1015_d 0.00284812f $X=4.29 $Y=1.445 $X2=0 $Y2=0
cc_270 N_B1_c_253_n N_A_523_297#_c_677_n 0.0114346f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B1_c_254_n N_A_523_297#_c_677_n 0.0138233f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B1_c_260_n N_A_523_297#_c_677_n 0.0104094f $X=4.245 $Y=1.572 $X2=0
+ $Y2=0
cc_273 B1 N_A_523_297#_c_677_n 0.00808046f $X=4.29 $Y=1.445 $X2=0 $Y2=0
cc_274 B1 N_A_523_297#_c_692_n 0.00197158f $X=4.29 $Y=1.445 $X2=0 $Y2=0
cc_275 N_B1_c_260_n A_613_297# 0.00200696f $X=4.245 $Y=1.572 $X2=-0.19 $Y2=-0.24
cc_276 N_B1_c_260_n A_805_297# 0.00299875f $X=4.245 $Y=1.572 $X2=-0.19 $Y2=-0.24
cc_277 B1 A_805_297# 0.00118775f $X=4.29 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_278 N_B1_M1007_g N_VGND_c_749_n 0.00422112f $X=2.905 $Y=0.56 $X2=0 $Y2=0
cc_279 N_B1_M1007_g N_VGND_c_753_n 0.00173477f $X=2.905 $Y=0.56 $X2=0 $Y2=0
cc_280 N_B1_c_255_n N_VGND_c_754_n 0.00422112f $X=4.55 $Y=0.985 $X2=0 $Y2=0
cc_281 N_B1_M1007_g N_VGND_c_757_n 0.00593073f $X=2.905 $Y=0.56 $X2=0 $Y2=0
cc_282 N_B1_c_255_n N_VGND_c_757_n 0.00643864f $X=4.55 $Y=0.985 $X2=0 $Y2=0
cc_283 N_B1_M1007_g N_VGND_c_760_n 5.36007e-19 $X=2.905 $Y=0.56 $X2=0 $Y2=0
cc_284 N_B1_c_255_n N_VGND_c_761_n 0.00343161f $X=4.55 $Y=0.985 $X2=0 $Y2=0
cc_285 N_C1_c_345_n N_VPWR_c_513_n 0.00429453f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_286 N_C1_c_346_n N_VPWR_c_513_n 0.00429453f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_287 N_C1_c_345_n N_VPWR_c_505_n 0.00618304f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_288 N_C1_c_346_n N_VPWR_c_505_n 0.0062771f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_289 N_C1_c_345_n N_A_523_297#_c_677_n 0.0146835f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_290 N_C1_c_346_n N_A_523_297#_c_677_n 0.0169151f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_291 N_C1_c_341_n N_VGND_c_749_n 0.00393972f $X=3.375 $Y=0.99 $X2=0 $Y2=0
cc_292 N_C1_c_342_n N_VGND_c_754_n 0.00422112f $X=3.96 $Y=0.99 $X2=0 $Y2=0
cc_293 N_C1_c_341_n N_VGND_c_757_n 0.00466358f $X=3.375 $Y=0.99 $X2=0 $Y2=0
cc_294 N_C1_c_342_n N_VGND_c_757_n 0.00653865f $X=3.96 $Y=0.99 $X2=0 $Y2=0
cc_295 N_C1_c_341_n N_VGND_c_760_n 0.00908582f $X=3.375 $Y=0.99 $X2=0 $Y2=0
cc_296 N_C1_c_342_n N_VGND_c_760_n 0.00550932f $X=3.96 $Y=0.99 $X2=0 $Y2=0
cc_297 N_A2_M1002_g N_A1_M1016_g 0.0426728f $X=5.18 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A2_c_387_n N_A1_c_463_n 0.0293762f $X=5.045 $Y=1.41 $X2=0 $Y2=0
cc_299 N_A2_c_391_n N_A1_c_463_n 0.00239464f $X=5.11 $Y=1.16 $X2=0 $Y2=0
cc_300 A2 N_A1_c_463_n 0.0141047f $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_301 N_A2_c_390_n N_A1_c_464_n 0.0355989f $X=6.595 $Y=1.41 $X2=0 $Y2=0
cc_302 A2 N_A1_c_464_n 0.0132131f $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_303 N_A2_c_416_p N_A1_c_464_n 0.00447766f $X=6.285 $Y=1.51 $X2=0 $Y2=0
cc_304 N_A2_c_389_n N_A1_M1014_g 0.0291905f $X=6.57 $Y=1.01 $X2=0 $Y2=0
cc_305 N_A2_c_387_n A1 0.00110216f $X=5.045 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A2_c_391_n A1 0.0200884f $X=5.11 $Y=1.16 $X2=0 $Y2=0
cc_307 N_A2_c_392_n A1 0.02175f $X=6.445 $Y=1.17 $X2=0 $Y2=0
cc_308 A2 A1 0.0257689f $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_309 N_A2_c_387_n N_A1_c_462_n 0.0248139f $X=5.045 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A2_c_390_n N_A1_c_462_n 0.0291905f $X=6.595 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A2_c_391_n N_A1_c_462_n 0.00112976f $X=5.11 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A2_c_392_n N_A1_c_462_n 0.0154437f $X=6.445 $Y=1.17 $X2=0 $Y2=0
cc_313 A2 N_A1_c_462_n 0.0111763f $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_314 N_A2_c_391_n N_VPWR_M1000_d 3.18056e-19 $X=5.11 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A2_c_428_p N_VPWR_M1000_d 0.001561f $X=5.325 $Y=1.605 $X2=0 $Y2=0
cc_316 A2 N_VPWR_M1000_d 0.00829608f $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_317 A2 N_VPWR_M1018_d 3.07655e-19 $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_318 N_A2_c_416_p N_VPWR_M1018_d 0.00428417f $X=6.285 $Y=1.51 $X2=0 $Y2=0
cc_319 N_A2_c_387_n N_VPWR_c_513_n 0.0032362f $X=5.045 $Y=1.41 $X2=0 $Y2=0
cc_320 N_A2_c_390_n N_VPWR_c_514_n 0.00465343f $X=6.595 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A2_c_387_n N_VPWR_c_505_n 0.00415547f $X=5.045 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A2_c_390_n N_VPWR_c_505_n 0.00629694f $X=6.595 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A2_c_387_n N_VPWR_c_518_n 0.0101529f $X=5.045 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A2_c_390_n N_VPWR_c_519_n 0.0078402f $X=6.595 $Y=1.41 $X2=0 $Y2=0
cc_325 A2 N_A_523_297#_M1008_s 0.00374184f $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_326 N_A2_c_387_n N_A_523_297#_c_696_n 0.0155072f $X=5.045 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A2_c_428_p N_A_523_297#_c_696_n 0.0238756f $X=5.325 $Y=1.605 $X2=0
+ $Y2=0
cc_328 A2 N_A_523_297#_c_696_n 0.0192901f $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_329 N_A2_c_387_n N_A_523_297#_c_699_n 5.24704e-19 $X=5.045 $Y=1.41 $X2=0
+ $Y2=0
cc_330 N_A2_c_390_n N_A_523_297#_c_700_n 0.011017f $X=6.595 $Y=1.41 $X2=0 $Y2=0
cc_331 N_A2_c_393_n N_A_523_297#_c_700_n 0.00405193f $X=6.66 $Y=1.16 $X2=0 $Y2=0
cc_332 A2 N_A_523_297#_c_700_n 0.00663989f $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_333 N_A2_c_416_p N_A_523_297#_c_700_n 0.0203906f $X=6.285 $Y=1.51 $X2=0 $Y2=0
cc_334 A2 N_A_523_297#_c_704_n 0.0191386f $X=6.125 $Y=1.445 $X2=0 $Y2=0
cc_335 N_A2_c_390_n N_A_523_297#_c_679_n 0.0209541f $X=6.595 $Y=1.41 $X2=0 $Y2=0
cc_336 N_A2_c_393_n N_A_523_297#_c_679_n 0.0152882f $X=6.66 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A2_c_416_p N_A_523_297#_c_679_n 0.0137613f $X=6.285 $Y=1.51 $X2=0 $Y2=0
cc_338 N_A2_c_389_n N_VGND_c_750_n 0.0171058f $X=6.57 $Y=1.01 $X2=0 $Y2=0
cc_339 N_A2_c_390_n N_VGND_c_750_n 0.00528052f $X=6.595 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A2_c_393_n N_VGND_c_750_n 0.0154635f $X=6.66 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A2_M1002_g N_VGND_c_755_n 0.00422112f $X=5.18 $Y=0.56 $X2=0 $Y2=0
cc_342 N_A2_c_389_n N_VGND_c_755_n 0.0046653f $X=6.57 $Y=1.01 $X2=0 $Y2=0
cc_343 N_A2_M1002_g N_VGND_c_757_n 0.00634927f $X=5.18 $Y=0.56 $X2=0 $Y2=0
cc_344 N_A2_c_389_n N_VGND_c_757_n 0.00802136f $X=6.57 $Y=1.01 $X2=0 $Y2=0
cc_345 N_A2_M1002_g N_VGND_c_761_n 0.00667888f $X=5.18 $Y=0.56 $X2=0 $Y2=0
cc_346 N_A1_c_463_n N_VPWR_c_511_n 0.00480127f $X=5.635 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A1_c_464_n N_VPWR_c_511_n 0.0032362f $X=6.115 $Y=1.41 $X2=0 $Y2=0
cc_348 N_A1_c_463_n N_VPWR_c_505_n 0.00679819f $X=5.635 $Y=1.41 $X2=0 $Y2=0
cc_349 N_A1_c_464_n N_VPWR_c_505_n 0.00384231f $X=6.115 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A1_c_463_n N_VPWR_c_518_n 0.00514469f $X=5.635 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A1_c_463_n N_VPWR_c_519_n 0.00108115f $X=5.635 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A1_c_464_n N_VPWR_c_519_n 0.00998776f $X=6.115 $Y=1.41 $X2=0 $Y2=0
cc_353 N_A1_c_463_n N_A_523_297#_c_696_n 0.0100405f $X=5.635 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A1_c_463_n N_A_523_297#_c_699_n 0.00733886f $X=5.635 $Y=1.41 $X2=0
+ $Y2=0
cc_355 N_A1_c_464_n N_A_523_297#_c_700_n 0.0153525f $X=6.115 $Y=1.41 $X2=0 $Y2=0
cc_356 N_A1_c_463_n N_A_523_297#_c_704_n 0.00517473f $X=5.635 $Y=1.41 $X2=0
+ $Y2=0
cc_357 N_A1_c_464_n N_A_523_297#_c_679_n 0.00114565f $X=6.115 $Y=1.41 $X2=0
+ $Y2=0
cc_358 N_A1_M1014_g N_VGND_c_750_n 0.00283791f $X=6.14 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A1_M1016_g N_VGND_c_755_n 0.00413555f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A1_M1014_g N_VGND_c_755_n 0.00585385f $X=6.14 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A1_M1016_g N_VGND_c_757_n 0.00600542f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A1_M1014_g N_VGND_c_757_n 0.0110535f $X=6.14 $Y=0.56 $X2=0 $Y2=0
cc_363 N_VPWR_c_505_n N_X_M1003_s 0.00638521f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_364 N_VPWR_c_505_n N_X_M1010_s 0.00621163f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_365 N_VPWR_M1003_d N_X_c_620_n 2.08577e-19 $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_366 N_VPWR_c_507_n N_X_c_620_n 0.00204919f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_367 N_VPWR_M1003_d N_X_c_615_n 0.00330363f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_368 N_VPWR_c_507_n N_X_c_615_n 0.0225608f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_369 N_VPWR_c_507_n N_X_c_622_n 0.0359873f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_370 N_VPWR_c_512_n N_X_c_622_n 0.0128338f $X=1.05 $Y=2.72 $X2=0 $Y2=0
cc_371 N_VPWR_c_505_n N_X_c_622_n 0.00704243f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_372 N_VPWR_M1009_d N_X_c_623_n 0.00354449f $X=1.065 $Y=1.485 $X2=0 $Y2=0
cc_373 N_VPWR_c_508_n N_X_c_623_n 0.0174312f $X=1.215 $Y=1.96 $X2=0 $Y2=0
cc_374 N_VPWR_c_509_n N_X_c_655_n 0.0131506f $X=2.01 $Y=2.72 $X2=0 $Y2=0
cc_375 N_VPWR_c_505_n N_X_c_655_n 0.00722976f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_376 N_VPWR_c_505_n N_A_523_297#_M1017_d 0.00217543f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_377 N_VPWR_c_505_n N_A_523_297#_M1015_d 0.0034615f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_505_n N_A_523_297#_M1008_s 0.00256642f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_505_n N_A_523_297#_M1021_s 0.00234791f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_510_n N_A_523_297#_c_677_n 0.0140426f $X=2.17 $Y=2 $X2=0 $Y2=0
cc_381 N_VPWR_c_513_n N_A_523_297#_c_677_n 0.116226f $X=5.07 $Y=2.72 $X2=0 $Y2=0
cc_382 N_VPWR_c_505_n N_A_523_297#_c_677_n 0.0717296f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_383 N_VPWR_M1000_d N_A_523_297#_c_696_n 0.00698442f $X=5.135 $Y=1.485 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_511_n N_A_523_297#_c_696_n 0.00329637f $X=6.14 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_513_n N_A_523_297#_c_696_n 0.00257431f $X=5.07 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_505_n N_A_523_297#_c_696_n 0.0117323f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_518_n N_A_523_297#_c_696_n 0.0244273f $X=5.285 $Y=2.36 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_511_n N_A_523_297#_c_699_n 0.0192787f $X=6.14 $Y=2.72 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_505_n N_A_523_297#_c_699_n 0.0114454f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_518_n N_A_523_297#_c_699_n 0.0126177f $X=5.285 $Y=2.36 $X2=0
+ $Y2=0
cc_391 N_VPWR_M1018_d N_A_523_297#_c_700_n 0.00386906f $X=6.205 $Y=1.485 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_511_n N_A_523_297#_c_700_n 0.00257431f $X=6.14 $Y=2.72 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_514_n N_A_523_297#_c_700_n 0.00165794f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_505_n N_A_523_297#_c_700_n 0.00843115f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_519_n N_A_523_297#_c_700_n 0.0199172f $X=6.355 $Y=2.36 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_514_n N_A_523_297#_c_678_n 0.0178099f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_505_n N_A_523_297#_c_678_n 0.00973825f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_513_n N_A_523_297#_c_692_n 0.0217227f $X=5.07 $Y=2.72 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_505_n N_A_523_297#_c_692_n 0.0125773f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_514_n N_A_523_297#_c_679_n 0.00184338f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_505_n N_A_523_297#_c_679_n 0.00334754f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_505_n A_613_297# 0.00240926f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_403 N_VPWR_c_505_n A_805_297# 0.00273049f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_404 N_X_c_612_n N_VGND_M1001_s 0.00655026f $X=1.085 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_405 N_X_c_627_n N_VGND_M1004_s 0.00420374f $X=2.045 $Y=0.745 $X2=0 $Y2=0
cc_406 N_X_c_612_n N_VGND_c_751_n 0.00270726f $X=1.085 $Y=0.755 $X2=0 $Y2=0
cc_407 N_X_c_614_n N_VGND_c_751_n 0.00517761f $X=0.212 $Y=0.875 $X2=0 $Y2=0
cc_408 N_X_c_612_n N_VGND_c_752_n 0.0033205f $X=1.085 $Y=0.755 $X2=0 $Y2=0
cc_409 N_X_c_662_p N_VGND_c_752_n 0.0127531f $X=1.18 $Y=0.42 $X2=0 $Y2=0
cc_410 N_X_c_627_n N_VGND_c_752_n 0.00266569f $X=2.045 $Y=0.745 $X2=0 $Y2=0
cc_411 N_X_c_627_n N_VGND_c_753_n 0.00349644f $X=2.045 $Y=0.745 $X2=0 $Y2=0
cc_412 N_X_c_634_n N_VGND_c_753_n 0.0252583f $X=2.14 $Y=0.42 $X2=0 $Y2=0
cc_413 N_X_M1001_d N_VGND_c_757_n 0.0031086f $X=0.99 $Y=0.235 $X2=0 $Y2=0
cc_414 N_X_M1005_d N_VGND_c_757_n 0.00770447f $X=1.95 $Y=0.235 $X2=0 $Y2=0
cc_415 N_X_c_612_n N_VGND_c_757_n 0.0115989f $X=1.085 $Y=0.755 $X2=0 $Y2=0
cc_416 N_X_c_662_p N_VGND_c_757_n 0.00722272f $X=1.18 $Y=0.42 $X2=0 $Y2=0
cc_417 N_X_c_627_n N_VGND_c_757_n 0.0119153f $X=2.045 $Y=0.745 $X2=0 $Y2=0
cc_418 N_X_c_634_n N_VGND_c_757_n 0.00683853f $X=2.14 $Y=0.42 $X2=0 $Y2=0
cc_419 N_X_c_614_n N_VGND_c_757_n 0.00767249f $X=0.212 $Y=0.875 $X2=0 $Y2=0
cc_420 N_X_c_612_n N_VGND_c_758_n 0.0250061f $X=1.085 $Y=0.755 $X2=0 $Y2=0
cc_421 N_X_c_662_p N_VGND_c_758_n 0.0129599f $X=1.18 $Y=0.42 $X2=0 $Y2=0
cc_422 N_X_c_627_n N_VGND_c_759_n 0.0202592f $X=2.045 $Y=0.745 $X2=0 $Y2=0
cc_423 N_X_c_634_n N_VGND_c_759_n 0.0116788f $X=2.14 $Y=0.42 $X2=0 $Y2=0
cc_424 N_A_523_297#_c_677_n A_613_297# 0.00377586f $X=4.57 $Y=2.337 $X2=-0.19
+ $Y2=1.305
cc_425 N_A_523_297#_c_677_n A_805_297# 0.00633152f $X=4.57 $Y=2.337 $X2=-0.19
+ $Y2=1.305
cc_426 N_VGND_c_757_n A_1051_47# 0.00318969f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
cc_427 N_VGND_c_757_n A_1243_47# 0.0119688f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
