* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VGND a_36_47# a_209_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_36_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VPWR a_209_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 X a_209_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VPWR A1 a_647_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_1115_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_647_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_935_47# A1 a_209_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_209_21# A1 a_1115_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_209_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_36_47# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_647_297# a_36_47# a_209_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VPWR A2 a_647_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_209_21# a_36_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_647_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 X a_209_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND A2 a_935_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_209_21# a_36_47# a_647_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND a_209_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 X a_209_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 VPWR a_209_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 X a_209_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
