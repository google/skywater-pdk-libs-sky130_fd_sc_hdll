* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__muxb16to1_1 D[15] D[14] D[13] D[12] D[11] D[10] D[9] D[8]
+ D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] S[15] S[14] S[13] S[12] S[11] S[10] S[9]
+ S[8] S[7] S[6] S[5] S[4] S[3] S[2] S[1] S[0] VGND VNB VPB VPWR Z
X0 VGND S[11] a_1361_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X1 VPWR D[8] a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VPWR S[1] a_533_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_109_911# S[8] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X4 VGND D[2] a_937_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_1840_265# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_1012_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X7 VGND D[4] a_1765_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_3218_333# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VGND D[10] a_937_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_2402_47# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND S[7] a_3017_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X12 VPWR S[13] a_2189_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VPWR D[4] a_1773_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VPWR D[10] a_945_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VPWR S[15] a_3017_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 Z S[7] a_3230_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X17 a_937_911# S[10] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X18 a_2390_333# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_1574_47# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_1765_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X21 a_1012_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_1765_911# S[12] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X23 VPWR S[11] a_1361_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 a_109_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X26 VGND S[13] a_2189_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X27 Z a_3017_937# a_3218_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X28 a_2593_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X29 VGND S[9] a_533_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X30 a_117_591# a_184_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X31 Z a_533_937# a_734_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X32 VGND S[15] a_3017_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X33 a_1562_591# D[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 VPWR D[2] a_945_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 VPWR S[5] a_2189_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X36 a_2668_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X37 Z S[13] a_2402_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X38 VPWR S[7] a_3017_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 VGND D[8] a_109_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X40 a_3230_937# D[15] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 Z a_2189_937# a_2390_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X42 a_2601_591# a_2668_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X43 VPWR S[3] a_1361_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 Z a_3017_47# a_3218_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X45 Z S[11] a_1574_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X46 a_117_297# a_184_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X47 Z a_533_47# a_734_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X48 a_184_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X49 VGND S[3] a_1361_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X50 a_1840_793# S[12] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X51 VGND D[14] a_2593_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X52 a_2593_911# S[14] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X53 VGND S[1] a_533_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X54 a_184_793# S[8] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X55 a_2402_937# D[13] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 a_2668_793# S[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 a_734_591# D[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X58 a_945_591# a_1012_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X59 a_2668_793# S[14] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 Z a_1361_937# a_1562_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X61 a_1562_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 a_1773_591# a_1840_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X63 Z a_2189_47# a_2390_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X64 VGND S[5] a_2189_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X65 a_746_937# D[9] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X66 a_2601_297# a_2668_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X67 a_1012_793# S[10] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X68 a_184_793# S[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X69 VGND D[12] a_1765_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X70 Z S[15] a_3230_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X71 Z S[5] a_2402_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X72 a_1574_937# D[11] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X73 VPWR D[14] a_2601_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X74 a_945_297# a_1012_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X75 VGND D[0] a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X76 Z a_1361_47# a_1562_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X77 a_937_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X78 VPWR S[9] a_533_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X79 a_3218_591# D[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X80 a_1773_297# a_1840_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X81 Z S[3] a_1574_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X82 a_2668_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X83 a_1840_793# S[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X84 Z S[1] a_746_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X85 VPWR D[12] a_1773_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X86 a_734_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X87 Z S[9] a_746_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X88 a_2390_591# D[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X89 VGND D[6] a_2593_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X90 a_1012_793# S[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X91 a_184_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X92 a_746_47# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X93 a_1840_265# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X94 a_3230_47# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X95 VPWR D[6] a_2601_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
