* File: sky130_fd_sc_hdll__diode_6.pxi.spice
* Created: Thu Aug 27 19:05:18 2020
* 
x_PM_SKY130_FD_SC_HDLL__DIODE_6%DIODE N_DIODE_D0_noxref_neg DIODE DIODE
+ N_DIODE_c_8_n PM_SKY130_FD_SC_HDLL__DIODE_6%DIODE
x_PM_SKY130_FD_SC_HDLL__DIODE_6%VGND VGND N_VGND_c_15_n N_VGND_c_16_n
+ PM_SKY130_FD_SC_HDLL__DIODE_6%VGND
x_PM_SKY130_FD_SC_HDLL__DIODE_6%VPWR VPWR N_VPWR_c_21_n N_VPWR_c_20_n
+ PM_SKY130_FD_SC_HDLL__DIODE_6%VPWR
cc_1 VNB N_DIODE_c_8_n 0.152104f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=0.37
cc_2 VNB N_VGND_c_15_n 0.0678606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_3 VNB N_VGND_c_16_n 0.161822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_4 VNB N_VPWR_c_20_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VPB N_DIODE_c_8_n 0.183015f $X=-0.19 $Y=1.305 $X2=2.415 $Y2=0.37
cc_6 VPB N_VPWR_c_21_n 0.0678606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_7 VPB N_VPWR_c_20_n 0.0641928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_8 N_DIODE_c_8_n N_VGND_c_15_n 0.181108f $X=2.415 $Y=0.37 $X2=0 $Y2=0
cc_9 N_DIODE_D0_noxref_neg N_VGND_c_16_n 0.023764f $X=0.135 $Y=0.195 $X2=0 $Y2=0
cc_10 N_DIODE_c_8_n N_VGND_c_16_n 0.099699f $X=2.415 $Y=0.37 $X2=0 $Y2=0
cc_11 N_DIODE_c_8_n N_VPWR_c_21_n 0.184527f $X=2.415 $Y=0.37 $X2=0 $Y2=0
cc_12 N_DIODE_c_8_n N_VPWR_c_20_n 0.099699f $X=2.415 $Y=0.37 $X2=0 $Y2=0
