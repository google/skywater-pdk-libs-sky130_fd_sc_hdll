* File: sky130_fd_sc_hdll__a21o_2.pxi.spice
* Created: Thu Aug 27 18:52:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21O_2%A_80_21# N_A_80_21#_M1006_d N_A_80_21#_M1004_s
+ N_A_80_21#_c_49_n N_A_80_21#_M1003_g N_A_80_21#_c_50_n N_A_80_21#_c_56_n
+ N_A_80_21#_M1002_g N_A_80_21#_c_51_n N_A_80_21#_c_52_n N_A_80_21#_M1005_g
+ N_A_80_21#_c_53_n N_A_80_21#_M1007_g N_A_80_21#_c_54_n N_A_80_21#_c_55_n
+ N_A_80_21#_c_62_p N_A_80_21#_c_102_p N_A_80_21#_c_59_n N_A_80_21#_c_78_p
+ N_A_80_21#_c_72_p N_A_80_21#_c_60_n PM_SKY130_FD_SC_HDLL__A21O_2%A_80_21#
x_PM_SKY130_FD_SC_HDLL__A21O_2%B1 N_B1_c_122_n N_B1_M1006_g N_B1_c_123_n
+ N_B1_M1004_g B1 PM_SKY130_FD_SC_HDLL__A21O_2%B1
x_PM_SKY130_FD_SC_HDLL__A21O_2%A1 N_A1_c_149_n N_A1_M1008_g N_A1_c_150_n
+ N_A1_M1001_g A1 A1 PM_SKY130_FD_SC_HDLL__A21O_2%A1
x_PM_SKY130_FD_SC_HDLL__A21O_2%A2 N_A2_c_185_n N_A2_M1009_g N_A2_c_186_n
+ N_A2_M1000_g A2 A2 PM_SKY130_FD_SC_HDLL__A21O_2%A2
x_PM_SKY130_FD_SC_HDLL__A21O_2%VPWR N_VPWR_M1002_s N_VPWR_M1005_s N_VPWR_M1001_d
+ N_VPWR_c_212_n N_VPWR_c_213_n N_VPWR_c_214_n N_VPWR_c_215_n N_VPWR_c_216_n
+ VPWR N_VPWR_c_217_n N_VPWR_c_218_n N_VPWR_c_211_n N_VPWR_c_220_n
+ PM_SKY130_FD_SC_HDLL__A21O_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A21O_2%X N_X_M1003_d N_X_M1002_d X N_X_c_261_n
+ PM_SKY130_FD_SC_HDLL__A21O_2%X
x_PM_SKY130_FD_SC_HDLL__A21O_2%A_444_297# N_A_444_297#_M1004_d
+ N_A_444_297#_M1000_d N_A_444_297#_c_281_n N_A_444_297#_c_290_n
+ N_A_444_297#_c_282_n N_A_444_297#_c_286_n N_A_444_297#_c_295_n
+ PM_SKY130_FD_SC_HDLL__A21O_2%A_444_297#
x_PM_SKY130_FD_SC_HDLL__A21O_2%VGND N_VGND_M1003_s N_VGND_M1007_s N_VGND_M1009_d
+ N_VGND_c_297_n N_VGND_c_298_n N_VGND_c_299_n N_VGND_c_300_n VGND
+ N_VGND_c_301_n N_VGND_c_302_n N_VGND_c_303_n N_VGND_c_304_n
+ PM_SKY130_FD_SC_HDLL__A21O_2%VGND
cc_1 VNB N_A_80_21#_c_49_n 0.0228695f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A_80_21#_c_50_n 0.0135094f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.31
cc_3 VNB N_A_80_21#_c_51_n 0.0185942f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=1.07
cc_4 VNB N_A_80_21#_c_52_n 0.0220188f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=1.41
cc_5 VNB N_A_80_21#_c_53_n 0.0212709f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_6 VNB N_A_80_21#_c_54_n 0.0114746f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.07
cc_7 VNB N_A_80_21#_c_55_n 0.00511977f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.16
cc_8 VNB N_B1_c_122_n 0.0217557f $X=-0.19 $Y=-0.24 $X2=2.02 $Y2=0.235
cc_9 VNB N_B1_c_123_n 0.029135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB B1 0.00744892f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_11 VNB N_A1_c_149_n 0.0177278f $X=-0.19 $Y=-0.24 $X2=2.02 $Y2=0.235
cc_12 VNB N_A1_c_150_n 0.0231799f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB A1 0.00426382f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_14 VNB N_A2_c_185_n 0.0201519f $X=-0.19 $Y=-0.24 $X2=2.02 $Y2=0.235
cc_15 VNB N_A2_c_186_n 0.0320172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB A2 0.0215441f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_17 VNB N_VPWR_c_211_n 0.155873f $X=-0.19 $Y=-0.24 $X2=2.155 $Y2=0.42
cc_18 VNB N_X_c_261_n 0.00160788f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.145
cc_19 VNB N_VGND_c_297_n 0.0110262f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.145
cc_20 VNB N_VGND_c_298_n 0.00472864f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_21 VNB N_VGND_c_299_n 0.0129243f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.985
cc_22 VNB N_VGND_c_300_n 0.0166106f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.07
cc_23 VNB N_VGND_c_301_n 0.025615f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_24 VNB N_VGND_c_302_n 0.0407742f $X=-0.19 $Y=-0.24 $X2=1.212 $Y2=1.69
cc_25 VNB N_VGND_c_303_n 0.01325f $X=-0.19 $Y=-0.24 $X2=2.145 $Y2=0.655
cc_26 VNB N_VGND_c_304_n 0.20296f $X=-0.19 $Y=-0.24 $X2=1.072 $Y2=1.16
cc_27 VPB N_A_80_21#_c_56_n 0.0305592f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_28 VPB N_A_80_21#_c_52_n 0.029534f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.41
cc_29 VPB N_A_80_21#_c_55_n 0.00253533f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.16
cc_30 VPB N_A_80_21#_c_59_n 0.0138064f $X=-0.19 $Y=1.305 $X2=1.675 $Y2=1.805
cc_31 VPB N_A_80_21#_c_60_n 0.00935252f $X=-0.19 $Y=1.305 $X2=1.84 $Y2=1.88
cc_32 VPB N_B1_c_123_n 0.0320907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB B1 0.00517668f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_34 VPB N_A1_c_150_n 0.0258916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB A1 0.00159181f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_36 VPB N_A2_c_186_n 0.0357032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB A2 0.00429335f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_38 VPB N_VPWR_c_212_n 0.0105879f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.145
cc_39 VPB N_VPWR_c_213_n 0.0379095f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_40 VPB N_VPWR_c_214_n 0.00561386f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.07
cc_41 VPB N_VPWR_c_215_n 0.0332141f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.985
cc_42 VPB N_VPWR_c_216_n 0.00632158f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=0.995
cc_43 VPB N_VPWR_c_217_n 0.0178083f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.07
cc_44 VPB N_VPWR_c_218_n 0.0206176f $X=-0.19 $Y=1.305 $X2=2.145 $Y2=0.42
cc_45 VPB N_VPWR_c_211_n 0.0504597f $X=-0.19 $Y=1.305 $X2=2.155 $Y2=0.42
cc_46 VPB N_VPWR_c_220_n 0.0130464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_X_c_261_n 0.00127832f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.145
cc_48 N_A_80_21#_c_55_n N_B1_c_122_n 0.00488357f $X=1.08 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_49 N_A_80_21#_c_62_p N_B1_c_122_n 0.0141619f $X=2.05 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_50 N_A_80_21#_c_52_n N_B1_c_123_n 0.00374157f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_51 N_A_80_21#_c_55_n N_B1_c_123_n 0.00888783f $X=1.08 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_80_21#_c_62_p N_B1_c_123_n 0.00130243f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_53 N_A_80_21#_c_60_n N_B1_c_123_n 0.0069822f $X=1.84 $Y=1.88 $X2=0 $Y2=0
cc_54 N_A_80_21#_c_52_n B1 0.00104495f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_55 N_A_80_21#_c_55_n B1 0.0186103f $X=1.08 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_80_21#_c_62_p B1 0.0268871f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_57 N_A_80_21#_c_60_n B1 0.00893004f $X=1.84 $Y=1.88 $X2=0 $Y2=0
cc_58 N_A_80_21#_c_62_p N_A1_c_149_n 6.14218e-19 $X=2.05 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_59 N_A_80_21#_c_72_p N_A1_c_149_n 0.0031074f $X=2.155 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_60 N_A_80_21#_M1006_d A1 0.00566932f $X=2.02 $Y=0.235 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_62_p A1 0.0144463f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_72_p A1 0.0222491f $X=2.155 $Y=0.42 $X2=0 $Y2=0
cc_63 N_A_80_21#_c_55_n N_VPWR_M1005_s 0.00516635f $X=1.08 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_59_n N_VPWR_M1005_s 9.21288e-19 $X=1.675 $Y=1.805 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_78_p N_VPWR_M1005_s 0.00519994f $X=1.43 $Y=1.805 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_56_n N_VPWR_c_213_n 0.00684339f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_80_21#_c_60_n N_VPWR_c_215_n 0.023629f $X=1.84 $Y=1.88 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_56_n N_VPWR_c_217_n 0.00635665f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_52_n N_VPWR_c_217_n 0.00448795f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_80_21#_M1004_s N_VPWR_c_211_n 0.00262606f $X=1.715 $Y=1.485 $X2=0
+ $Y2=0
cc_71 N_A_80_21#_c_56_n N_VPWR_c_211_n 0.0119178f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_52_n N_VPWR_c_211_n 0.00602407f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_59_n N_VPWR_c_211_n 0.00720548f $X=1.675 $Y=1.805 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_78_p N_VPWR_c_211_n 0.00388719f $X=1.43 $Y=1.805 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_60_n N_VPWR_c_211_n 0.0139798f $X=1.84 $Y=1.88 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_56_n N_VPWR_c_220_n 0.00101786f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_52_n N_VPWR_c_220_n 0.012565f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_59_n N_VPWR_c_220_n 0.00275096f $X=1.675 $Y=1.805 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_78_p N_VPWR_c_220_n 0.0163583f $X=1.43 $Y=1.805 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_60_n N_VPWR_c_220_n 0.0193958f $X=1.84 $Y=1.88 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_49_n N_X_c_261_n 0.025942f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_50_n N_X_c_261_n 0.00907092f $X=0.5 $Y=1.31 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_56_n N_X_c_261_n 0.031066f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_51_n N_X_c_261_n 0.0129612f $X=0.93 $Y=1.07 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_52_n N_X_c_261_n 0.0155122f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_53_n N_X_c_261_n 0.00983596f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_54_n N_X_c_261_n 0.00685943f $X=0.5 $Y=1.07 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_55_n N_X_c_261_n 0.0678249f $X=1.08 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_102_p N_X_c_261_n 0.0138428f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_78_p N_X_c_261_n 0.0187283f $X=1.43 $Y=1.805 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_55_n N_VGND_M1007_s 0.00107595f $X=1.08 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_62_p N_VGND_M1007_s 0.022301f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_102_p N_VGND_M1007_s 0.00452573f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_49_n N_VGND_c_298_n 0.00434782f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_49_n N_VGND_c_301_n 0.00579312f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_53_n N_VGND_c_301_n 0.00443627f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_102_p N_VGND_c_301_n 0.00447787f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_62_p N_VGND_c_302_n 0.00579931f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_72_p N_VGND_c_302_n 0.0121687f $X=2.155 $Y=0.42 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_53_n N_VGND_c_303_n 0.0091493f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_62_p N_VGND_c_303_n 0.014206f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_102_p N_VGND_c_303_n 0.0107715f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_80_21#_M1006_d N_VGND_c_304_n 0.0100715f $X=2.02 $Y=0.235 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_49_n N_VGND_c_304_n 0.0117373f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_53_n N_VGND_c_304_n 0.00816998f $X=1.055 $Y=0.995 $X2=0
+ $Y2=0
cc_106 N_A_80_21#_c_62_p N_VGND_c_304_n 0.011313f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_102_p N_VGND_c_304_n 0.00848677f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_72_p N_VGND_c_304_n 0.00720706f $X=2.155 $Y=0.42 $X2=0 $Y2=0
cc_109 N_B1_c_122_n N_A1_c_149_n 0.0143322f $X=1.945 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_110 N_B1_c_123_n N_A1_c_150_n 0.038581f $X=2.13 $Y=1.41 $X2=0 $Y2=0
cc_111 B1 N_A1_c_150_n 0.00277365f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_112 N_B1_c_122_n A1 0.00422125f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B1_c_123_n A1 0.00112461f $X=2.13 $Y=1.41 $X2=0 $Y2=0
cc_114 B1 A1 0.0276751f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_115 N_B1_c_123_n N_VPWR_c_215_n 0.00702461f $X=2.13 $Y=1.41 $X2=0 $Y2=0
cc_116 N_B1_c_123_n N_VPWR_c_211_n 0.0140657f $X=2.13 $Y=1.41 $X2=0 $Y2=0
cc_117 N_B1_c_123_n N_VPWR_c_220_n 0.00274938f $X=2.13 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B1_c_122_n N_VGND_c_302_n 0.00428022f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B1_c_122_n N_VGND_c_303_n 0.00813254f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B1_c_122_n N_VGND_c_304_n 0.00773499f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A1_c_149_n N_A2_c_185_n 0.0276193f $X=2.585 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_122 A1 N_A2_c_185_n 0.00738688f $X=2.465 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_123 N_A1_c_150_n N_A2_c_186_n 0.0548295f $X=2.61 $Y=1.41 $X2=0 $Y2=0
cc_124 A1 N_A2_c_186_n 0.00123506f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_125 N_A1_c_149_n A2 2.35582e-19 $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A1_c_150_n A2 9.83094e-19 $X=2.61 $Y=1.41 $X2=0 $Y2=0
cc_127 A1 A2 0.021279f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_128 N_A1_c_150_n N_VPWR_c_214_n 0.00337394f $X=2.61 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A1_c_150_n N_VPWR_c_215_n 0.00702461f $X=2.61 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A1_c_150_n N_VPWR_c_211_n 0.00713365f $X=2.61 $Y=1.41 $X2=0 $Y2=0
cc_131 A1 N_A_444_297#_c_281_n 0.0035028f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_132 N_A1_c_150_n N_A_444_297#_c_282_n 0.0172236f $X=2.61 $Y=1.41 $X2=0 $Y2=0
cc_133 A1 N_A_444_297#_c_282_n 0.00962215f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_134 N_A1_c_149_n N_VGND_c_300_n 0.00170451f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_135 A1 N_VGND_c_300_n 0.00771888f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_136 N_A1_c_149_n N_VGND_c_302_n 0.0037962f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_137 A1 N_VGND_c_302_n 0.0105675f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_138 N_A1_c_149_n N_VGND_c_304_n 0.00608811f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_139 A1 N_VGND_c_304_n 0.0108043f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_140 A1 A_532_47# 0.00713993f $X=2.465 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_141 N_A2_c_186_n N_VPWR_c_214_n 0.00336725f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A2_c_186_n N_VPWR_c_218_n 0.00700684f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A2_c_186_n N_VPWR_c_211_n 0.00802756f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A2_c_186_n N_A_444_297#_c_282_n 0.0192586f $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_145 A2 N_A_444_297#_c_282_n 0.00331088f $X=3.31 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A2_c_186_n N_A_444_297#_c_286_n 0.00255101f $X=3.125 $Y=1.41 $X2=0
+ $Y2=0
cc_147 A2 N_A_444_297#_c_286_n 0.0109464f $X=3.31 $Y=1.105 $X2=0 $Y2=0
cc_148 A2 N_VGND_M1009_d 0.00328988f $X=3.31 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A2_c_185_n N_VGND_c_300_n 0.0116645f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A2_c_186_n N_VGND_c_300_n 8.22261e-19 $X=3.125 $Y=1.41 $X2=0 $Y2=0
cc_151 A2 N_VGND_c_300_n 0.0252488f $X=3.31 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A2_c_185_n N_VGND_c_302_n 0.00505556f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A2_c_185_n N_VGND_c_304_n 0.00883429f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_154 A2 N_VGND_c_304_n 0.00158513f $X=3.31 $Y=1.105 $X2=0 $Y2=0
cc_155 N_VPWR_c_211_n N_X_M1002_d 0.00682945f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_c_217_n N_X_c_261_n 0.0174364f $X=1.055 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_211_n N_X_c_261_n 0.0104326f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_c_220_n N_X_c_261_n 0.0151867f $X=1.27 $Y=2.34 $X2=0 $Y2=0
cc_159 N_VPWR_c_211_n N_A_444_297#_M1004_d 0.00397303f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_160 N_VPWR_c_211_n N_A_444_297#_M1000_d 0.00277788f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_161 N_VPWR_c_215_n N_A_444_297#_c_290_n 0.0143924f $X=2.705 $Y=2.72 $X2=0
+ $Y2=0
cc_162 N_VPWR_c_211_n N_A_444_297#_c_290_n 0.00858812f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_163 N_VPWR_M1001_d N_A_444_297#_c_282_n 0.0107461f $X=2.7 $Y=1.485 $X2=0
+ $Y2=0
cc_164 N_VPWR_c_214_n N_A_444_297#_c_282_n 0.0164279f $X=2.87 $Y=2.34 $X2=0
+ $Y2=0
cc_165 N_VPWR_c_211_n N_A_444_297#_c_282_n 0.0148682f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_166 N_VPWR_c_218_n N_A_444_297#_c_295_n 0.0147725f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_167 N_VPWR_c_211_n N_A_444_297#_c_295_n 0.00839556f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_168 N_X_c_261_n N_VGND_c_301_n 0.017522f $X=0.74 $Y=0.42 $X2=0 $Y2=0
cc_169 N_X_c_261_n N_VGND_c_303_n 0.00740115f $X=0.74 $Y=0.42 $X2=0 $Y2=0
cc_170 N_X_M1003_d N_VGND_c_304_n 0.00887224f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_171 N_X_c_261_n N_VGND_c_304_n 0.0106155f $X=0.74 $Y=0.42 $X2=0 $Y2=0
cc_172 N_VGND_c_304_n A_532_47# 0.0132386f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
