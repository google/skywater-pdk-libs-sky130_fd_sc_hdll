* File: sky130_fd_sc_hdll__clkbuf_8.spice
* Created: Wed Sep  2 08:25:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkbuf_8.pex.spice"
.subckt sky130_fd_sc_hdll__clkbuf_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_A_118_297#_M1001_d N_A_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.1323 PD=0.75 PS=1.47 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.2
+ SB=75004.5 A=0.063 P=1.14 MULT=1
MM1002 N_A_118_297#_M1001_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0588 PD=0.75 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75004 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1002_s N_A_118_297#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0693 PD=0.7 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_118_297#_M1007_g N_X_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1007_d N_A_118_297#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_118_297#_M1009_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1009_d N_A_118_297#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.1
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_118_297#_M1014_g N_X_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.5
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1014_d N_A_118_297#_M1016_g N_X_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0798 PD=0.75 PS=0.8 NRD=0 NRS=14.28 M=1 R=2.8 SA=75004
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_118_297#_M1018_g N_X_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.0798 PD=1.38 PS=0.8 NRD=1.428 NRS=14.28 M=1 R=2.8 SA=75004.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_118_297#_M1004_d N_A_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1013 N_A_118_297#_M1004_d N_A_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90004 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1013_s N_A_118_297#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_118_297#_M1005_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.6
+ SB=90003.1 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1005_d N_A_118_297#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.1
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_118_297#_M1010_g N_X_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.6
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1010_d N_A_118_297#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.1
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_A_118_297#_M1015_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.5
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1015_d N_A_118_297#_M1017_g N_X_M1017_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90004
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1019_d N_A_118_297#_M1019_g N_X_M1017_s VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90004.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hdll__clkbuf_8.pxi.spice"
*
.ends
*
*
