# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.175000 1.075000 9.635000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.255000 0.995000 8.475000 1.445000 ;
        RECT 8.255000 1.445000 8.640000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.130000 0.995000 3.815000 1.325000 ;
    END
  END C
  PIN VGND
    ANTENNADIFFAREA  1.225400 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.490800 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.645000 0.350000 0.815000 0.660000 ;
        RECT 0.645000 0.660000 1.755000 0.925000 ;
        RECT 0.745000 1.440000 1.570000 1.455000 ;
        RECT 0.745000 1.455000 1.855000 2.045000 ;
        RECT 0.745000 2.045000 0.915000 2.465000 ;
        RECT 1.205000 0.925000 1.570000 1.440000 ;
        RECT 1.585000 0.350000 1.755000 0.660000 ;
        RECT 1.685000 2.045000 1.855000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.175000  0.085000  0.345000 0.545000 ;
      RECT  0.275000  2.135000  0.445000 2.635000 ;
      RECT  0.985000  0.085000  1.365000 0.465000 ;
      RECT  1.135000  2.215000  1.465000 2.635000 ;
      RECT  2.020000  0.965000  2.245000 1.325000 ;
      RECT  2.055000  0.085000  2.225000 0.525000 ;
      RECT  2.075000  0.695000  2.565000 0.865000 ;
      RECT  2.075000  0.865000  2.245000 0.965000 ;
      RECT  2.075000  1.325000  2.245000 1.875000 ;
      RECT  2.075000  1.875000  2.795000 2.045000 ;
      RECT  2.075000  2.215000  2.405000 2.635000 ;
      RECT  2.395000  0.255000  4.060000 0.425000 ;
      RECT  2.395000  0.425000  2.565000 0.695000 ;
      RECT  2.570000  1.535000  4.155000 1.705000 ;
      RECT  2.575000  2.045000  2.795000 2.235000 ;
      RECT  2.575000  2.235000  4.215000 2.405000 ;
      RECT  2.790000  0.595000  2.960000 1.535000 ;
      RECT  3.140000  1.895000  4.545000 2.065000 ;
      RECT  3.240000  0.655000  4.450000 0.825000 ;
      RECT  3.660000  0.425000  4.060000 0.455000 ;
      RECT  3.985000  0.995000  4.405000 1.325000 ;
      RECT  3.985000  1.325000  4.155000 1.535000 ;
      RECT  4.230000  0.255000  5.130000 0.425000 ;
      RECT  4.230000  0.425000  4.450000 0.655000 ;
      RECT  4.375000  1.525000  4.905000 1.695000 ;
      RECT  4.375000  1.695000  4.545000 1.895000 ;
      RECT  4.480000  2.235000  4.885000 2.405000 ;
      RECT  4.620000  0.595000  4.790000 1.375000 ;
      RECT  4.620000  1.375000  4.905000 1.525000 ;
      RECT  4.715000  1.895000  5.990000 2.065000 ;
      RECT  4.715000  2.065000  4.885000 2.235000 ;
      RECT  4.960000  0.425000  5.130000 1.035000 ;
      RECT  4.960000  1.035000  5.215000 1.040000 ;
      RECT  4.960000  1.040000  5.230000 1.045000 ;
      RECT  4.960000  1.045000  5.240000 1.050000 ;
      RECT  4.960000  1.050000  5.245000 1.205000 ;
      RECT  5.055000  2.235000  5.385000 2.635000 ;
      RECT  5.075000  1.205000  5.245000 1.895000 ;
      RECT  5.300000  0.085000  5.470000 0.885000 ;
      RECT  5.475000  1.445000  5.990000 1.715000 ;
      RECT  5.700000  0.415000  5.990000 1.445000 ;
      RECT  5.820000  2.065000  5.990000 2.275000 ;
      RECT  5.820000  2.275000  9.115000 2.445000 ;
      RECT  6.165000  0.265000  6.580000 0.485000 ;
      RECT  6.165000  0.485000  6.385000 0.595000 ;
      RECT  6.165000  0.595000  6.335000 2.105000 ;
      RECT  6.525000  0.720000  6.970000 0.825000 ;
      RECT  6.525000  0.825000  6.775000 0.890000 ;
      RECT  6.525000  0.890000  6.695000 2.275000 ;
      RECT  6.555000  0.655000  6.970000 0.720000 ;
      RECT  6.800000  0.320000  6.970000 0.655000 ;
      RECT  6.915000  1.445000  7.745000 1.615000 ;
      RECT  6.915000  1.615000  7.330000 2.045000 ;
      RECT  6.930000  0.995000  7.355000 1.270000 ;
      RECT  7.140000  0.630000  7.355000 0.995000 ;
      RECT  7.575000  0.255000  8.770000 0.425000 ;
      RECT  7.575000  0.425000  7.745000 1.445000 ;
      RECT  7.915000  0.595000  8.085000 1.935000 ;
      RECT  7.915000  1.935000 10.425000 2.105000 ;
      RECT  8.255000  0.425000  8.770000 0.465000 ;
      RECT  8.645000  0.730000  8.850000 0.945000 ;
      RECT  8.645000  0.945000  8.955000 1.275000 ;
      RECT  9.105000  1.495000  9.975000 1.705000 ;
      RECT  9.145000  0.295000  9.435000 0.735000 ;
      RECT  9.145000  0.735000  9.975000 0.750000 ;
      RECT  9.185000  0.750000  9.975000 0.905000 ;
      RECT  9.615000  2.275000  9.945000 2.635000 ;
      RECT  9.695000  0.085000  9.865000 0.565000 ;
      RECT  9.805000  0.905000  9.975000 0.995000 ;
      RECT  9.805000  0.995000 10.035000 1.325000 ;
      RECT  9.805000  1.325000  9.975000 1.495000 ;
      RECT  9.890000  1.875000 10.425000 1.935000 ;
      RECT 10.165000  0.255000 10.425000 0.585000 ;
      RECT 10.165000  2.105000 10.425000 2.465000 ;
      RECT 10.255000  0.585000 10.425000 1.875000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.735000  1.445000  4.905000 1.615000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.705000  0.765000  5.875000 0.935000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.215000  0.425000  6.385000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.185000  0.765000  7.355000 0.935000 ;
      RECT  7.185000  1.445000  7.355000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.665000  0.765000  8.835000 0.935000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.175000  0.425000  9.345000 0.595000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.460000 7.415000 1.600000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
      RECT 5.645000 0.735000 5.985000 0.780000 ;
      RECT 5.645000 0.780000 8.895000 0.920000 ;
      RECT 5.645000 0.920000 5.985000 0.965000 ;
      RECT 6.155000 0.395000 6.445000 0.440000 ;
      RECT 6.155000 0.440000 9.405000 0.580000 ;
      RECT 6.155000 0.580000 6.445000 0.625000 ;
      RECT 7.125000 0.735000 7.415000 0.780000 ;
      RECT 7.125000 0.920000 7.415000 0.965000 ;
      RECT 7.125000 1.415000 7.415000 1.460000 ;
      RECT 7.125000 1.600000 7.415000 1.645000 ;
      RECT 8.605000 0.735000 8.895000 0.780000 ;
      RECT 8.605000 0.920000 8.895000 0.965000 ;
      RECT 9.115000 0.395000 9.405000 0.440000 ;
      RECT 9.115000 0.580000 9.405000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor3_4
END LIBRARY
