* File: sky130_fd_sc_hdll__nor3b_1.pex.spice
* Created: Thu Aug 27 19:16:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR3B_1%A_91_199# 1 2 7 9 10 12 13 19 20 21 25 27
r56 24 27 4.85669 $w=3.14e-07 $l=2.65236e-07 $layer=LI1_cond $X=2.59 $Y=0.825
+ $X2=2.465 $Y2=0.615
r57 24 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.59 $Y=0.825
+ $X2=2.59 $Y2=1.785
r58 21 23 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=0.885 $Y=1.87
+ $X2=2.465 $Y2=1.87
r59 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=1.87
+ $X2=2.59 $Y2=1.785
r60 20 23 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.505 $Y=1.87
+ $X2=2.465 $Y2=1.87
r61 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.8 $Y=1.785
+ $X2=0.885 $Y2=1.87
r62 18 19 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.8 $Y=1.245 $X2=0.8
+ $Y2=1.785
r63 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r64 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.715 $Y=1.16
+ $X2=0.8 $Y2=1.245
r65 13 15 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.715 $Y=1.16
+ $X2=0.59 $Y2=1.16
r66 10 16 38.8967 $w=3.59e-07 $l=2.18746e-07 $layer=POLY_cond $X=0.78 $Y=0.995
+ $X2=0.655 $Y2=1.16
r67 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.78 $Y=0.995
+ $X2=0.78 $Y2=0.56
r68 7 16 45.5371 $w=3.59e-07 $l=2.95804e-07 $layer=POLY_cond $X=0.755 $Y=1.41
+ $X2=0.655 $Y2=1.16
r69 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.755 $Y=1.41
+ $X2=0.755 $Y2=1.985
r70 2 23 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.65 $X2=2.465 $Y2=1.87
r71 1 27 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=2.33
+ $Y=0.465 $X2=2.465 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_1%B 1 3 4 6 7
r30 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2 $Y=1.16
+ $X2=1.2 $Y2=1.16
r31 4 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.25 $Y=0.995
+ $X2=1.225 $Y2=1.16
r32 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.25 $Y=0.995 $X2=1.25
+ $Y2=0.56
r33 1 10 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.225 $Y=1.41
+ $X2=1.225 $Y2=1.16
r34 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.225 $Y=1.41
+ $X2=1.225 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_1%A 1 3 4 6 7 13
r30 7 13 2.31499 $w=6.18e-07 $l=1.2e-07 $layer=LI1_cond $X=1.73 $Y=1.305
+ $X2=1.61 $Y2=1.305
r31 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.16 $X2=1.73 $Y2=1.16
r32 4 10 48.651 $w=2.87e-07 $l=2.76134e-07 $layer=POLY_cond $X=1.695 $Y=1.41
+ $X2=1.75 $Y2=1.16
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.695 $Y=1.41
+ $X2=1.695 $Y2=1.985
r34 1 10 38.6443 $w=2.87e-07 $l=2.0106e-07 $layer=POLY_cond $X=1.67 $Y=0.995
+ $X2=1.75 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.67 $Y=0.995 $X2=1.67
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_1%C_N 2 3 5 8 9 12 14
r33 12 15 37.7413 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.16
+ $X2=2.28 $Y2=1.325
r34 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.16
+ $X2=2.28 $Y2=0.995
r35 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r36 8 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.255 $Y=0.675
+ $X2=2.255 $Y2=0.995
r37 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.23 $Y=1.575
+ $X2=2.23 $Y2=1.86
r38 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.23 $Y=1.475 $X2=2.23
+ $Y2=1.575
r39 2 15 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.23 $Y=1.475 $X2=2.23
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_1%Y 1 2 3 10 14 18 22 23
r34 27 35 0.650043 $w=4.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.315 $Y=1.675
+ $X2=0.315 $Y2=1.65
r35 23 27 5.17174 $w=4.6e-07 $l=1.95e-07 $layer=LI1_cond $X=0.315 $Y=1.87
+ $X2=0.315 $Y2=1.675
r36 22 35 3.1202 $w=4.58e-07 $l=1.2e-07 $layer=LI1_cond $X=0.315 $Y=1.53
+ $X2=0.315 $Y2=1.65
r37 21 22 26.7323 $w=2.78e-07 $l=6.2e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.445
r38 20 21 7.80118 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.345 $Y2=0.825
r39 18 20 8.05053 $w=5.18e-07 $l=3.5e-07 $layer=LI1_cond $X=0.345 $Y=0.39
+ $X2=0.345 $Y2=0.74
r40 12 14 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.46 $Y=0.655
+ $X2=1.46 $Y2=0.495
r41 11 20 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.74
+ $X2=0.345 $Y2=0.74
r42 10 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.375 $Y=0.74
+ $X2=1.46 $Y2=0.655
r43 10 11 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.375 $Y=0.74
+ $X2=0.605 $Y2=0.74
r44 3 35 300 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=2 $X=0.335
+ $Y=1.485 $X2=0.46 $Y2=1.65
r45 2 14 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.325
+ $Y=0.235 $X2=1.46 $Y2=0.495
r46 1 18 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.315
+ $Y=0.235 $X2=0.44 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_1%VPWR 1 6 9 10 11 21 22
r27 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r28 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r29 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r30 14 18 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r31 11 19 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r32 11 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r33 9 18 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.715 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 9 10 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.715 $Y=2.72
+ $X2=1.905 $Y2=2.72
r35 8 21 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.095 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 8 10 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.095 $Y=2.72
+ $X2=1.905 $Y2=2.72
r37 4 10 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=2.635
+ $X2=1.905 $Y2=2.72
r38 4 6 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=1.905 $Y=2.635
+ $X2=1.905 $Y2=2.21
r39 1 6 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=1.785
+ $Y=1.485 $X2=1.93 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_1%VGND 1 2 9 13 16 17 19 20 21 31 32
r39 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r40 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r41 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r42 25 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r43 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r44 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r45 19 28 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.715 $Y=0 $X2=1.61
+ $Y2=0
r46 19 20 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.715 $Y=0 $X2=1.905
+ $Y2=0
r47 18 31 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.53
+ $Y2=0
r48 18 20 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=1.905
+ $Y2=0
r49 16 24 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.69
+ $Y2=0
r50 16 17 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.965
+ $Y2=0
r51 15 28 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.61
+ $Y2=0
r52 15 17 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=0.965
+ $Y2=0
r53 11 20 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=0.085
+ $X2=1.905 $Y2=0
r54 11 13 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=1.905 $Y=0.085
+ $X2=1.905 $Y2=0.39
r55 7 17 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=0.085
+ $X2=0.965 $Y2=0
r56 7 9 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.965 $Y=0.085
+ $X2=0.965 $Y2=0.39
r57 2 13 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.745
+ $Y=0.235 $X2=1.93 $Y2=0.39
r58 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.855
+ $Y=0.235 $X2=0.99 $Y2=0.39
.ends

