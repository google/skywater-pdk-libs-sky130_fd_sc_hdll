* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1612_47# a_1188_47# a_1403_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1403_21# a_1188_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 a_865_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1188_47# a_27_47# a_1317_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X5 a_1317_47# a_1403_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_1403_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 Q a_1403_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR RESET_B a_699_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X9 a_1188_47# a_211_363# a_1388_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X10 Q a_1403_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VGND a_27_47# a_211_363# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR RESET_B a_1403_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X13 a_699_413# a_811_289# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X14 a_689_47# a_811_289# a_865_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_811_289# a_27_47# a_1188_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X16 a_583_47# a_211_363# a_689_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VPWR D a_468_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X18 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_468_47# a_27_47# a_583_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X20 VPWR a_1403_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VGND RESET_B a_1612_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 Q a_1403_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR a_27_47# a_211_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X24 a_1388_413# a_1403_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X25 a_811_289# a_211_363# a_1188_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X26 VGND a_583_47# a_811_289# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 VGND a_1403_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_583_47# a_27_47# a_699_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X29 VGND D a_468_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_468_47# a_211_363# a_583_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X31 VPWR a_583_47# a_811_289# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X32 Q a_1403_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 VGND a_1403_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
