* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_525_413# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X1 a_79_21# a_243_47# a_525_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_241_297# A2_N a_243_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X4 VGND A1_N a_243_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR A1_N a_241_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X6 a_243_47# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_79_21# B2 a_611_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_611_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR B1 a_525_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X11 VGND a_243_47# a_79_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
