# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__ebufn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__ebufn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.765000 0.775000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.516600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.765000 1.300000 1.275000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.445000 4.460000 1.625000 ;
        RECT 1.985000 1.625000 3.995000 1.765000 ;
        RECT 3.545000 0.635000 4.460000 0.855000 ;
        RECT 3.595000 1.765000 3.995000 2.125000 ;
        RECT 4.230000 0.855000 4.460000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.900000 0.595000 ;
      RECT 0.515000  1.845000 1.000000 2.635000 ;
      RECT 1.070000  0.255000 1.830000 0.595000 ;
      RECT 1.220000  1.445000 1.815000 1.765000 ;
      RECT 1.220000  1.765000 1.510000 2.465000 ;
      RECT 1.550000  0.595000 1.830000 1.025000 ;
      RECT 1.550000  1.025000 3.215000 1.275000 ;
      RECT 1.550000  1.275000 1.815000 1.445000 ;
      RECT 1.700000  1.935000 3.375000 2.105000 ;
      RECT 1.700000  2.105000 1.910000 2.465000 ;
      RECT 2.000000  0.255000 2.320000 0.655000 ;
      RECT 2.000000  0.655000 3.375000 0.855000 ;
      RECT 2.080000  2.275000 2.460000 2.635000 ;
      RECT 2.490000  0.085000 2.870000 0.485000 ;
      RECT 2.680000  2.105000 3.375000 2.295000 ;
      RECT 2.680000  2.295000 4.425000 2.465000 ;
      RECT 3.090000  0.275000 4.400000 0.465000 ;
      RECT 3.090000  0.465000 3.375000 0.655000 ;
      RECT 3.495000  1.025000 3.955000 1.275000 ;
      RECT 4.165000  1.795000 4.425000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.150000  1.060000 0.320000 1.230000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.680000  1.060000 3.850000 1.230000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 1.030000 0.380000 1.120000 ;
      RECT 0.085000 1.120000 3.910000 1.260000 ;
      RECT 3.570000 1.030000 3.910000 1.120000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_2
END LIBRARY
