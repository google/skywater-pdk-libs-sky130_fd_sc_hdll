* File: sky130_fd_sc_hdll__o22a_4.spice
* Created: Thu Aug 27 19:21:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o22a_4.pex.spice"
.subckt sky130_fd_sc_hdll__o22a_4  VNB VPB B1 B2 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_X_M1007_d N_A_96_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.182 PD=0.97 PS=1.86 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1007_d N_A_96_21#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1014 N_X_M1014_d N_A_96_21#_M1014_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1015 N_X_M1014_d N_A_96_21#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_A_524_47#_M1009_d N_B1_M1009_g N_A_96_21#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1010 N_A_96_21#_M1009_s N_B2_M1010_g N_A_524_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1016 N_A_96_21#_M1016_d N_B2_M1016_g N_A_524_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1019 N_A_524_47#_M1019_d N_B1_M1019_g N_A_96_21#_M1016_d VNB NSHORT L=0.15
+ W=0.65 AD=0.13 AS=0.104 PD=1.05 PS=0.97 NRD=7.38 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A1_M1000_g N_A_524_47#_M1019_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.13 PD=0.92 PS=1.05 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75002.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1000_d N_A2_M1012_g N_A_524_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_A2_M1020_g N_A_524_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1020_d N_A1_M1004_g N_A_524_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_96_21#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90006 A=0.18 P=2.36 MULT=1
MM1005 N_X_M1001_d N_A_96_21#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90005.5 A=0.18 P=2.36 MULT=1
MM1018 N_X_M1018_d N_A_96_21#_M1018_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90005 A=0.18 P=2.36 MULT=1
MM1022 N_X_M1018_d N_A_96_21#_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.405 PD=1.29 PS=1.81 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90004.6 A=0.18 P=2.36 MULT=1
MM1013 N_A_614_297#_M1013_d N_B1_M1013_g N_VPWR_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.405 PD=1.29 PS=1.81 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90003.6 A=0.18 P=2.36 MULT=1
MM1003 N_A_614_297#_M1013_d N_B2_M1003_g N_A_96_21#_M1003_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1006 N_A_614_297#_M1006_d N_B2_M1006_g N_A_96_21#_M1003_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1023 N_A_614_297#_M1006_d N_B1_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.185 PD=1.29 PS=1.37 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1002 N_A_1006_297#_M1002_d N_A1_M1002_g N_VPWR_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.185 PD=1.29 PS=1.37 NRD=0.9653 NRS=16.7253 M=1 R=5.55556
+ SA=90004.6 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1017 N_A_1006_297#_M1002_d N_A2_M1017_g N_A_96_21#_M1017_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1021 N_A_1006_297#_M1021_d N_A2_M1021_g N_A_96_21#_M1017_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.5 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1011 N_A_1006_297#_M1021_d N_A1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.295 PD=1.29 PS=2.59 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90006
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=11.6844 P=17.77
pX25_noxref noxref_14 A2 A2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o22a_4.pxi.spice"
*
.ends
*
*
