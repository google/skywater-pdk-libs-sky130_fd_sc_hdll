* File: sky130_fd_sc_hdll__or4bb_4.pxi.spice
* Created: Wed Sep  2 08:50:12 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%C_N N_C_N_c_112_n N_C_N_c_113_n N_C_N_M1014_g
+ N_C_N_M1008_g C_N C_N N_C_N_c_109_n N_C_N_c_110_n N_C_N_c_111_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_4%C_N
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%D_N N_D_N_c_144_n N_D_N_M1017_g N_D_N_c_145_n
+ N_D_N_M1004_g D_N PM_SKY130_FD_SC_HDLL__OR4BB_4%D_N
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%A_224_297# N_A_224_297#_M1004_d
+ N_A_224_297#_M1017_d N_A_224_297#_c_181_n N_A_224_297#_M1001_g
+ N_A_224_297#_c_175_n N_A_224_297#_M1011_g N_A_224_297#_c_176_n
+ N_A_224_297#_c_177_n N_A_224_297#_c_184_n N_A_224_297#_c_185_n
+ N_A_224_297#_c_178_n N_A_224_297#_c_179_n N_A_224_297#_c_180_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_4%A_224_297#
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%A_27_410# N_A_27_410#_M1008_s
+ N_A_27_410#_M1014_s N_A_27_410#_c_240_n N_A_27_410#_M1010_g
+ N_A_27_410#_c_241_n N_A_27_410#_M1012_g N_A_27_410#_c_242_n
+ N_A_27_410#_c_247_n N_A_27_410#_c_248_n N_A_27_410#_c_249_n
+ N_A_27_410#_c_250_n N_A_27_410#_c_251_n N_A_27_410#_c_243_n
+ N_A_27_410#_c_244_n N_A_27_410#_c_253_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_4%A_27_410#
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%B N_B_c_321_n N_B_M1009_g N_B_c_322_n
+ N_B_M1005_g B B N_B_c_323_n PM_SKY130_FD_SC_HDLL__OR4BB_4%B
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%A N_A_c_352_n N_A_M1002_g N_A_c_353_n
+ N_A_M1003_g N_A_c_356_n N_A_c_354_n A A PM_SKY130_FD_SC_HDLL__OR4BB_4%A
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%A_335_297# N_A_335_297#_M1011_d
+ N_A_335_297#_M1005_d N_A_335_297#_M1001_s N_A_335_297#_c_390_n
+ N_A_335_297#_M1006_g N_A_335_297#_c_398_n N_A_335_297#_M1000_g
+ N_A_335_297#_c_391_n N_A_335_297#_M1013_g N_A_335_297#_c_399_n
+ N_A_335_297#_M1007_g N_A_335_297#_c_392_n N_A_335_297#_M1015_g
+ N_A_335_297#_c_400_n N_A_335_297#_M1016_g N_A_335_297#_c_401_n
+ N_A_335_297#_M1018_g N_A_335_297#_c_393_n N_A_335_297#_M1019_g
+ N_A_335_297#_c_402_n N_A_335_297#_c_394_n N_A_335_297#_c_419_n
+ N_A_335_297#_c_432_n N_A_335_297#_c_420_n N_A_335_297#_c_523_p
+ N_A_335_297#_c_442_n N_A_335_297#_c_395_n N_A_335_297#_c_396_n
+ N_A_335_297#_c_471_p N_A_335_297#_c_438_n N_A_335_297#_c_397_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_4%A_335_297#
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%VPWR N_VPWR_M1014_d N_VPWR_M1003_d
+ N_VPWR_M1007_s N_VPWR_M1018_s N_VPWR_c_539_n N_VPWR_c_540_n N_VPWR_c_541_n
+ N_VPWR_c_542_n N_VPWR_c_543_n N_VPWR_c_544_n N_VPWR_c_545_n N_VPWR_c_546_n
+ N_VPWR_c_547_n VPWR N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n
+ N_VPWR_c_538_n PM_SKY130_FD_SC_HDLL__OR4BB_4%VPWR
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%X N_X_M1006_d N_X_M1015_d N_X_M1000_d
+ N_X_M1016_d N_X_c_626_n N_X_c_670_n N_X_c_635_n N_X_c_627_n N_X_c_620_n
+ N_X_c_621_n N_X_c_653_n N_X_c_674_n N_X_c_628_n N_X_c_622_n N_X_c_623_n
+ N_X_c_629_n X N_X_c_625_n PM_SKY130_FD_SC_HDLL__OR4BB_4%X
x_PM_SKY130_FD_SC_HDLL__OR4BB_4%VGND N_VGND_M1008_d N_VGND_M1011_s
+ N_VGND_M1012_d N_VGND_M1002_d N_VGND_M1013_s N_VGND_M1019_s N_VGND_c_697_n
+ N_VGND_c_698_n N_VGND_c_699_n N_VGND_c_700_n N_VGND_c_701_n N_VGND_c_702_n
+ N_VGND_c_703_n N_VGND_c_704_n N_VGND_c_705_n N_VGND_c_706_n N_VGND_c_707_n
+ N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n VGND
+ N_VGND_c_712_n N_VGND_c_713_n N_VGND_c_714_n N_VGND_c_715_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_4%VGND
cc_1 VNB N_C_N_c_109_n 0.0256354f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_2 VNB N_C_N_c_110_n 0.00772584f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_3 VNB N_C_N_c_111_n 0.0212836f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.995
cc_4 VNB N_D_N_c_144_n 0.0281042f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_5 VNB N_D_N_c_145_n 0.0193872f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.26
cc_6 VNB D_N 0.00218634f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.675
cc_7 VNB N_A_224_297#_c_175_n 0.0201398f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_8 VNB N_A_224_297#_c_176_n 0.0254549f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.16
cc_9 VNB N_A_224_297#_c_177_n 0.0110628f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_10 VNB N_A_224_297#_c_178_n 0.0111709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_224_297#_c_179_n 0.00325774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_224_297#_c_180_n 0.0028325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_410#_c_240_n 0.0240813f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.675
cc_14 VNB N_A_27_410#_c_241_n 0.0174761f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_15 VNB N_A_27_410#_c_242_n 0.0213305f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_16 VNB N_A_27_410#_c_243_n 0.00111747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_410#_c_244_n 0.0183099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_c_321_n 0.0222503f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_19 VNB N_B_c_322_n 0.01695f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.26
cc_20 VNB N_B_c_323_n 0.00347568f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.16
cc_21 VNB N_A_c_352_n 0.0177141f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_22 VNB N_A_c_353_n 0.0245697f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.26
cc_23 VNB N_A_c_354_n 0.00110761f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_24 VNB N_A_335_297#_c_390_n 0.0170949f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_25 VNB N_A_335_297#_c_391_n 0.0167552f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.995
cc_26 VNB N_A_335_297#_c_392_n 0.0171975f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.53
cc_27 VNB N_A_335_297#_c_393_n 0.0200652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_335_297#_c_394_n 0.00288951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_335_297#_c_395_n 0.0016277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_335_297#_c_396_n 0.00466338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_335_297#_c_397_n 0.0717345f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_538_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_620_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_621_n 0.00175721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_622_n 6.97233e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_623_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB X 0.0187238f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_625_n 0.00760418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_697_n 0.0151513f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_698_n 0.0111532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_699_n 0.00218082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_700_n 0.00259443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_701_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_702_n 0.0108398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_703_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_704_n 0.0226239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_705_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_706_n 0.0212426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_707_n 0.00631534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_708_n 0.0161956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_709_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_710_n 0.0177951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_711_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_712_n 0.0171208f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_713_n 0.019291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_714_n 0.00609289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_715_n 0.321037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VPB N_C_N_c_112_n 0.0336446f $X=-0.19 $Y=1.285 $X2=0.495 $Y2=1.875
cc_59 VPB N_C_N_c_113_n 0.0283638f $X=-0.19 $Y=1.285 $X2=0.495 $Y2=1.975
cc_60 VPB N_C_N_c_109_n 0.00623853f $X=-0.19 $Y=1.285 $X2=0.52 $Y2=1.16
cc_61 VPB N_C_N_c_110_n 0.00263638f $X=-0.19 $Y=1.285 $X2=0.52 $Y2=1.16
cc_62 VPB N_D_N_c_144_n 0.0316212f $X=-0.19 $Y=1.285 $X2=0.495 $Y2=1.325
cc_63 VPB D_N 6.63091e-19 $X=-0.19 $Y=1.285 $X2=0.555 $Y2=0.675
cc_64 VPB N_A_224_297#_c_181_n 0.0194802f $X=-0.19 $Y=1.285 $X2=0.555 $Y2=0.675
cc_65 VPB N_A_224_297#_c_176_n 0.012942f $X=-0.19 $Y=1.285 $X2=0.535 $Y2=1.16
cc_66 VPB N_A_224_297#_c_177_n 0.00700747f $X=-0.19 $Y=1.285 $X2=0.52 $Y2=1.16
cc_67 VPB N_A_224_297#_c_184_n 0.00974573f $X=-0.19 $Y=1.285 $X2=0.52 $Y2=1.16
cc_68 VPB N_A_224_297#_c_185_n 0.00431421f $X=-0.19 $Y=1.285 $X2=0.63 $Y2=1.53
cc_69 VPB N_A_224_297#_c_179_n 0.00187624f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_70 VPB N_A_27_410#_c_240_n 0.0293863f $X=-0.19 $Y=1.285 $X2=0.555 $Y2=0.675
cc_71 VPB N_A_27_410#_c_242_n 0.0287885f $X=-0.19 $Y=1.285 $X2=0.52 $Y2=1.16
cc_72 VPB N_A_27_410#_c_247_n 0.0146752f $X=-0.19 $Y=1.285 $X2=0.535 $Y2=1.325
cc_73 VPB N_A_27_410#_c_248_n 0.00874217f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_74 VPB N_A_27_410#_c_249_n 0.00665675f $X=-0.19 $Y=1.285 $X2=0.63 $Y2=1.53
cc_75 VPB N_A_27_410#_c_250_n 0.00759776f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_76 VPB N_A_27_410#_c_251_n 0.00398727f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_77 VPB N_A_27_410#_c_243_n 0.00100873f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_78 VPB N_A_27_410#_c_253_n 0.0107579f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_79 VPB N_B_c_321_n 0.0272744f $X=-0.19 $Y=1.285 $X2=0.495 $Y2=1.325
cc_80 VPB N_B_c_323_n 0.00255428f $X=-0.19 $Y=1.285 $X2=0.535 $Y2=1.16
cc_81 VPB N_A_c_353_n 0.0280012f $X=-0.19 $Y=1.285 $X2=0.495 $Y2=2.26
cc_82 VPB N_A_c_356_n 0.00297959f $X=-0.19 $Y=1.285 $X2=0.555 $Y2=0.675
cc_83 VPB N_A_c_354_n 0.00102254f $X=-0.19 $Y=1.285 $X2=0.605 $Y2=1.105
cc_84 VPB N_A_335_297#_c_398_n 0.0171379f $X=-0.19 $Y=1.285 $X2=0.535 $Y2=1.16
cc_85 VPB N_A_335_297#_c_399_n 0.0159747f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_86 VPB N_A_335_297#_c_400_n 0.0159552f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_87 VPB N_A_335_297#_c_401_n 0.0191382f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_88 VPB N_A_335_297#_c_402_n 0.00299875f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_89 VPB N_A_335_297#_c_394_n 0.00123572f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_90 VPB N_A_335_297#_c_397_n 0.0509526f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_539_n 0.00718943f $X=-0.19 $Y=1.285 $X2=0.52 $Y2=1.16
cc_92 VPB N_VPWR_c_540_n 0.00519418f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_541_n 0.00516582f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_542_n 0.0112901f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_543_n 0.00518f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_544_n 0.0712566f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_545_n 0.0047828f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_546_n 0.0213107f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_547_n 0.0047828f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_548_n 0.014554f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_549_n 0.0195604f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_550_n 0.00593536f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_538_n 0.0554153f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_104 VPB N_X_c_626_n 0.0019666f $X=-0.19 $Y=1.285 $X2=0.535 $Y2=1.16
cc_105 VPB N_X_c_627_n 0.00206401f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_106 VPB N_X_c_628_n 0.00817154f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_107 VPB N_X_c_629_n 0.00161374f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_108 VPB X 0.00823301f $X=-0.19 $Y=1.285 $X2=0 $Y2=0
cc_109 N_C_N_c_112_n N_D_N_c_144_n 0.0219419f $X=0.495 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_110 N_C_N_c_113_n N_D_N_c_144_n 0.00196013f $X=0.495 $Y=1.975 $X2=-0.19
+ $Y2=-0.24
cc_111 N_C_N_c_109_n N_D_N_c_144_n 0.017826f $X=0.52 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_112 N_C_N_c_110_n N_D_N_c_144_n 0.00984276f $X=0.52 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_113 N_C_N_c_111_n N_D_N_c_145_n 0.00921668f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_114 N_C_N_c_109_n D_N 2.94462e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_115 N_C_N_c_110_n D_N 0.0264894f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_116 N_C_N_c_112_n N_A_224_297#_c_184_n 2.80344e-19 $X=0.495 $Y=1.875 $X2=0
+ $Y2=0
cc_117 N_C_N_c_110_n N_A_224_297#_c_184_n 0.00929331f $X=0.52 $Y=1.16 $X2=0
+ $Y2=0
cc_118 N_C_N_c_112_n N_A_27_410#_c_242_n 0.0153708f $X=0.495 $Y=1.875 $X2=0
+ $Y2=0
cc_119 N_C_N_c_109_n N_A_27_410#_c_242_n 0.0078918f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_120 N_C_N_c_110_n N_A_27_410#_c_242_n 0.0532478f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_121 N_C_N_c_111_n N_A_27_410#_c_242_n 0.00504599f $X=0.535 $Y=0.995 $X2=0
+ $Y2=0
cc_122 N_C_N_c_113_n N_A_27_410#_c_247_n 0.00475322f $X=0.495 $Y=1.975 $X2=0
+ $Y2=0
cc_123 N_C_N_c_113_n N_A_27_410#_c_248_n 0.0170384f $X=0.495 $Y=1.975 $X2=0
+ $Y2=0
cc_124 N_C_N_c_109_n N_A_27_410#_c_248_n 8.16996e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_125 N_C_N_c_110_n N_A_27_410#_c_248_n 0.0269325f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_126 N_C_N_c_113_n N_A_27_410#_c_249_n 0.00245287f $X=0.495 $Y=1.975 $X2=0
+ $Y2=0
cc_127 N_C_N_c_109_n N_A_27_410#_c_244_n 0.00104536f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_128 N_C_N_c_111_n N_A_27_410#_c_244_n 0.00216055f $X=0.535 $Y=0.995 $X2=0
+ $Y2=0
cc_129 N_C_N_c_110_n N_VPWR_M1014_d 0.00455141f $X=0.52 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_130 N_C_N_c_113_n N_VPWR_c_539_n 0.0122493f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_131 N_C_N_c_113_n N_VPWR_c_548_n 0.00306699f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_132 N_C_N_c_113_n N_VPWR_c_538_n 0.00454334f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_133 N_C_N_c_110_n N_VGND_c_697_n 0.0108718f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_134 N_C_N_c_111_n N_VGND_c_697_n 0.00455093f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_135 N_C_N_c_111_n N_VGND_c_704_n 0.00510437f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_136 N_C_N_c_111_n N_VGND_c_715_n 0.00512902f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_137 N_D_N_c_144_n N_A_224_297#_c_176_n 0.0150381f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_138 D_N N_A_224_297#_c_176_n 9.72671e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_139 N_D_N_c_144_n N_A_224_297#_c_184_n 0.00876768f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_140 D_N N_A_224_297#_c_184_n 0.0153006f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_141 N_D_N_c_144_n N_A_224_297#_c_185_n 0.00558433f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_D_N_c_144_n N_A_224_297#_c_178_n 0.00272654f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_143 N_D_N_c_145_n N_A_224_297#_c_178_n 3.54632e-19 $X=1.05 $Y=0.995 $X2=0
+ $Y2=0
cc_144 D_N N_A_224_297#_c_178_n 0.012483f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_145 N_D_N_c_144_n N_A_224_297#_c_179_n 0.00101579f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_146 D_N N_A_224_297#_c_179_n 0.0272275f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_147 N_D_N_c_145_n N_A_224_297#_c_180_n 0.0042717f $X=1.05 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_D_N_c_144_n N_A_27_410#_c_248_n 0.0141438f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_149 D_N N_A_27_410#_c_248_n 0.00117737f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_150 N_D_N_c_144_n N_A_335_297#_c_402_n 3.45722e-19 $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_D_N_c_144_n N_VPWR_c_544_n 6.50559e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_152 N_D_N_c_145_n N_VGND_c_697_n 0.004325f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_153 N_D_N_c_145_n N_VGND_c_698_n 0.00311391f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_154 N_D_N_c_145_n N_VGND_c_706_n 0.00510437f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_155 N_D_N_c_145_n N_VGND_c_715_n 0.00512902f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_224_297#_c_181_n N_A_27_410#_c_240_n 0.0409425f $X=2.035 $Y=1.41
+ $X2=0 $Y2=0
cc_157 N_A_224_297#_c_177_n N_A_27_410#_c_240_n 0.0236026f $X=2.035 $Y=1.202
+ $X2=0 $Y2=0
cc_158 N_A_224_297#_c_175_n N_A_27_410#_c_241_n 0.0183508f $X=2.04 $Y=0.995
+ $X2=0 $Y2=0
cc_159 N_A_224_297#_M1017_d N_A_27_410#_c_248_n 0.00222919f $X=1.12 $Y=1.485
+ $X2=0 $Y2=0
cc_160 N_A_224_297#_c_184_n N_A_27_410#_c_248_n 0.022478f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_161 N_A_224_297#_c_181_n N_A_27_410#_c_249_n 0.00269387f $X=2.035 $Y=1.41
+ $X2=0 $Y2=0
cc_162 N_A_224_297#_c_181_n N_A_27_410#_c_250_n 0.0132574f $X=2.035 $Y=1.41
+ $X2=0 $Y2=0
cc_163 N_A_224_297#_c_184_n N_A_27_410#_c_250_n 0.00739005f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_164 N_A_224_297#_c_181_n N_A_27_410#_c_243_n 0.00510813f $X=2.035 $Y=1.41
+ $X2=0 $Y2=0
cc_165 N_A_224_297#_c_177_n N_A_27_410#_c_243_n 5.43086e-19 $X=2.035 $Y=1.202
+ $X2=0 $Y2=0
cc_166 N_A_224_297#_c_184_n N_A_335_297#_M1001_s 0.00244104f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_167 N_A_224_297#_c_185_n N_A_335_297#_M1001_s 9.10467e-19 $X=1.6 $Y=1.56
+ $X2=0 $Y2=0
cc_168 N_A_224_297#_c_181_n N_A_335_297#_c_402_n 0.0104787f $X=2.035 $Y=1.41
+ $X2=0 $Y2=0
cc_169 N_A_224_297#_c_176_n N_A_335_297#_c_402_n 0.00352492f $X=1.935 $Y=1.16
+ $X2=0 $Y2=0
cc_170 N_A_224_297#_c_184_n N_A_335_297#_c_402_n 0.0057931f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_171 N_A_224_297#_c_179_n N_A_335_297#_c_402_n 0.00260172f $X=1.71 $Y=1.16
+ $X2=0 $Y2=0
cc_172 N_A_224_297#_c_181_n N_A_335_297#_c_394_n 0.0199805f $X=2.035 $Y=1.41
+ $X2=0 $Y2=0
cc_173 N_A_224_297#_c_175_n N_A_335_297#_c_394_n 0.00492528f $X=2.04 $Y=0.995
+ $X2=0 $Y2=0
cc_174 N_A_224_297#_c_177_n N_A_335_297#_c_394_n 0.0128708f $X=2.035 $Y=1.202
+ $X2=0 $Y2=0
cc_175 N_A_224_297#_c_184_n N_A_335_297#_c_394_n 0.00791794f $X=1.505 $Y=1.645
+ $X2=0 $Y2=0
cc_176 N_A_224_297#_c_185_n N_A_335_297#_c_394_n 0.0100327f $X=1.6 $Y=1.56 $X2=0
+ $Y2=0
cc_177 N_A_224_297#_c_179_n N_A_335_297#_c_394_n 0.017853f $X=1.71 $Y=1.16 $X2=0
+ $Y2=0
cc_178 N_A_224_297#_c_180_n N_A_335_297#_c_394_n 0.00723177f $X=1.65 $Y=0.995
+ $X2=0 $Y2=0
cc_179 N_A_224_297#_c_175_n N_A_335_297#_c_419_n 0.00558723f $X=2.04 $Y=0.995
+ $X2=0 $Y2=0
cc_180 N_A_224_297#_c_175_n N_A_335_297#_c_420_n 0.00786296f $X=2.04 $Y=0.995
+ $X2=0 $Y2=0
cc_181 N_A_224_297#_c_178_n N_A_335_297#_c_420_n 0.00841259f $X=1.26 $Y=0.66
+ $X2=0 $Y2=0
cc_182 N_A_224_297#_c_181_n N_VPWR_c_544_n 0.00429453f $X=2.035 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_224_297#_c_181_n N_VPWR_c_538_n 0.00760487f $X=2.035 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_224_297#_c_178_n N_VGND_M1011_s 0.00280084f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_185 N_A_224_297#_c_180_n N_VGND_M1011_s 6.86606e-19 $X=1.65 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_224_297#_c_178_n N_VGND_c_697_n 0.00936362f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_187 N_A_224_297#_c_175_n N_VGND_c_698_n 0.00341589f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_224_297#_c_176_n N_VGND_c_698_n 0.0048595f $X=1.935 $Y=1.16 $X2=0
+ $Y2=0
cc_189 N_A_224_297#_c_178_n N_VGND_c_698_n 0.00836504f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_190 N_A_224_297#_c_179_n N_VGND_c_698_n 0.00340568f $X=1.71 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_A_224_297#_c_175_n N_VGND_c_699_n 7.4352e-19 $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_224_297#_c_178_n N_VGND_c_706_n 0.0100997f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_193 N_A_224_297#_c_175_n N_VGND_c_708_n 0.00501458f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_224_297#_c_175_n N_VGND_c_715_n 0.00957001f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_224_297#_c_178_n N_VGND_c_715_n 0.0138693f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_196 N_A_27_410#_c_240_n N_B_c_321_n 0.0736643f $X=2.565 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_197 N_A_27_410#_c_250_n N_B_c_321_n 5.49195e-19 $X=2.395 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_198 N_A_27_410#_c_243_n N_B_c_321_n 0.00130107f $X=2.48 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_199 N_A_27_410#_c_241_n N_B_c_322_n 0.0215187f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_27_410#_c_240_n N_B_c_323_n 0.00985564f $X=2.565 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_27_410#_c_250_n N_B_c_323_n 0.00445377f $X=2.395 $Y=2.38 $X2=0 $Y2=0
cc_202 N_A_27_410#_c_243_n N_B_c_323_n 0.0659017f $X=2.48 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_27_410#_c_250_n N_A_335_297#_M1001_s 0.00509651f $X=2.395 $Y=2.38
+ $X2=0 $Y2=0
cc_204 N_A_27_410#_c_240_n N_A_335_297#_c_402_n 5.77294e-19 $X=2.565 $Y=1.41
+ $X2=0 $Y2=0
cc_205 N_A_27_410#_c_248_n N_A_335_297#_c_402_n 0.00897715f $X=1.225 $Y=1.985
+ $X2=0 $Y2=0
cc_206 N_A_27_410#_c_249_n N_A_335_297#_c_402_n 0.0038017f $X=1.31 $Y=2.295
+ $X2=0 $Y2=0
cc_207 N_A_27_410#_c_250_n N_A_335_297#_c_402_n 0.0344881f $X=2.395 $Y=2.38
+ $X2=0 $Y2=0
cc_208 N_A_27_410#_c_243_n N_A_335_297#_c_402_n 0.0137192f $X=2.48 $Y=1.16 $X2=0
+ $Y2=0
cc_209 N_A_27_410#_c_240_n N_A_335_297#_c_394_n 0.00370199f $X=2.565 $Y=1.41
+ $X2=0 $Y2=0
cc_210 N_A_27_410#_c_241_n N_A_335_297#_c_394_n 0.00327649f $X=2.59 $Y=0.995
+ $X2=0 $Y2=0
cc_211 N_A_27_410#_c_248_n N_A_335_297#_c_394_n 0.00163234f $X=1.225 $Y=1.985
+ $X2=0 $Y2=0
cc_212 N_A_27_410#_c_243_n N_A_335_297#_c_394_n 0.0703486f $X=2.48 $Y=1.16 $X2=0
+ $Y2=0
cc_213 N_A_27_410#_c_241_n N_A_335_297#_c_432_n 0.0144855f $X=2.59 $Y=0.995
+ $X2=0 $Y2=0
cc_214 N_A_27_410#_c_240_n N_A_335_297#_c_420_n 0.00262417f $X=2.565 $Y=1.41
+ $X2=0 $Y2=0
cc_215 N_A_27_410#_c_243_n N_A_335_297#_c_420_n 0.0109703f $X=2.48 $Y=1.16 $X2=0
+ $Y2=0
cc_216 N_A_27_410#_c_248_n N_VPWR_M1014_d 0.00618252f $X=1.225 $Y=1.985
+ $X2=-0.19 $Y2=-0.24
cc_217 N_A_27_410#_c_247_n N_VPWR_c_539_n 0.0165151f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_218 N_A_27_410#_c_248_n N_VPWR_c_539_n 0.0243391f $X=1.225 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_A_27_410#_c_249_n N_VPWR_c_539_n 0.00276283f $X=1.31 $Y=2.295 $X2=0
+ $Y2=0
cc_220 N_A_27_410#_c_251_n N_VPWR_c_539_n 0.00957921f $X=1.395 $Y=2.38 $X2=0
+ $Y2=0
cc_221 N_A_27_410#_c_240_n N_VPWR_c_544_n 0.00565831f $X=2.565 $Y=1.41 $X2=0
+ $Y2=0
cc_222 N_A_27_410#_c_248_n N_VPWR_c_544_n 0.00582587f $X=1.225 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_27_410#_c_250_n N_VPWR_c_544_n 0.0697892f $X=2.395 $Y=2.38 $X2=0
+ $Y2=0
cc_224 N_A_27_410#_c_251_n N_VPWR_c_544_n 0.0120191f $X=1.395 $Y=2.38 $X2=0
+ $Y2=0
cc_225 N_A_27_410#_c_247_n N_VPWR_c_548_n 0.0163643f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_226 N_A_27_410#_c_248_n N_VPWR_c_548_n 0.00229383f $X=1.225 $Y=1.985 $X2=0
+ $Y2=0
cc_227 N_A_27_410#_c_240_n N_VPWR_c_538_n 0.00962783f $X=2.565 $Y=1.41 $X2=0
+ $Y2=0
cc_228 N_A_27_410#_c_247_n N_VPWR_c_538_n 0.00948926f $X=0.26 $Y=2.29 $X2=0
+ $Y2=0
cc_229 N_A_27_410#_c_248_n N_VPWR_c_538_n 0.0151126f $X=1.225 $Y=1.985 $X2=0
+ $Y2=0
cc_230 N_A_27_410#_c_250_n N_VPWR_c_538_n 0.0425445f $X=2.395 $Y=2.38 $X2=0
+ $Y2=0
cc_231 N_A_27_410#_c_251_n N_VPWR_c_538_n 0.00651555f $X=1.395 $Y=2.38 $X2=0
+ $Y2=0
cc_232 N_A_27_410#_c_250_n A_425_297# 0.00910103f $X=2.395 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_233 N_A_27_410#_c_243_n A_425_297# 0.00767598f $X=2.48 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_234 N_A_27_410#_c_244_n N_VGND_c_697_n 0.0185179f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_235 N_A_27_410#_c_241_n N_VGND_c_699_n 0.0105789f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_27_410#_c_244_n N_VGND_c_704_n 0.00926968f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_237 N_A_27_410#_c_241_n N_VGND_c_708_n 0.00199015f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_27_410#_c_241_n N_VGND_c_715_n 0.00298198f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A_27_410#_c_244_n N_VGND_c_715_n 0.0102233f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_240 N_B_c_322_n N_A_c_352_n 0.0249353f $X=3.06 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_241 N_B_c_321_n N_A_c_353_n 0.0748761f $X=3.035 $Y=1.41 $X2=0 $Y2=0
cc_242 N_B_c_323_n N_A_c_353_n 0.0019253f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B_c_321_n N_A_c_356_n 7.30212e-19 $X=3.035 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B_c_323_n N_A_c_356_n 0.0122483f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_245 N_B_c_321_n N_A_c_354_n 0.00118842f $X=3.035 $Y=1.41 $X2=0 $Y2=0
cc_246 N_B_c_323_n N_A_c_354_n 0.0184035f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_247 N_B_c_321_n N_A_335_297#_c_432_n 6.47027e-19 $X=3.035 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B_c_322_n N_A_335_297#_c_432_n 0.01167f $X=3.06 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B_c_323_n N_A_335_297#_c_432_n 0.020783f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_250 N_B_c_321_n N_A_335_297#_c_438_n 2.69871e-19 $X=3.035 $Y=1.41 $X2=0 $Y2=0
cc_251 N_B_c_321_n N_VPWR_c_544_n 0.00450951f $X=3.035 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B_c_323_n N_VPWR_c_544_n 0.0113003f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_253 N_B_c_321_n N_VPWR_c_538_n 0.00622433f $X=3.035 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_323_n N_VPWR_c_538_n 0.0100722f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B_c_323_n A_531_297# 0.00983665f $X=3.01 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_256 N_B_c_322_n N_VGND_c_699_n 0.00175252f $X=3.06 $Y=0.995 $X2=0 $Y2=0
cc_257 N_B_c_322_n N_VGND_c_712_n 0.00428022f $X=3.06 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B_c_322_n N_VGND_c_715_n 0.00585784f $X=3.06 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_c_352_n N_A_335_297#_c_390_n 0.0175202f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_c_353_n N_A_335_297#_c_398_n 0.0232871f $X=3.505 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_c_356_n N_A_335_297#_c_398_n 0.00237135f $X=3.565 $Y=1.4 $X2=0 $Y2=0
cc_262 N_A_c_352_n N_A_335_297#_c_442_n 0.012805f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A_c_353_n N_A_335_297#_c_442_n 0.00261534f $X=3.505 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_c_356_n N_A_335_297#_c_442_n 0.00215831f $X=3.565 $Y=1.4 $X2=0 $Y2=0
cc_265 N_A_c_354_n N_A_335_297#_c_442_n 0.0141192f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_c_352_n N_A_335_297#_c_395_n 0.00322035f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_c_353_n N_A_335_297#_c_395_n 5.08531e-19 $X=3.505 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_c_354_n N_A_335_297#_c_395_n 0.00579357f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_c_353_n N_A_335_297#_c_396_n 0.00124764f $X=3.505 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A_c_354_n N_A_335_297#_c_396_n 0.0139493f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_c_356_n N_A_335_297#_c_438_n 0.00124265f $X=3.565 $Y=1.4 $X2=0 $Y2=0
cc_272 N_A_c_353_n N_A_335_297#_c_397_n 0.0196968f $X=3.505 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A_c_354_n N_A_335_297#_c_397_n 0.00224534f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_c_356_n N_VPWR_M1003_d 0.00237148f $X=3.565 $Y=1.4 $X2=0 $Y2=0
cc_275 N_A_c_353_n N_VPWR_c_540_n 0.0113068f $X=3.505 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A_c_356_n N_VPWR_c_540_n 0.00110888f $X=3.565 $Y=1.4 $X2=0 $Y2=0
cc_277 N_A_c_353_n N_VPWR_c_544_n 0.00702461f $X=3.505 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_c_353_n N_VPWR_c_538_n 0.01287f $X=3.505 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A_c_356_n A_625_297# 0.00279786f $X=3.565 $Y=1.4 $X2=-0.19 $Y2=-0.24
cc_280 N_A_c_356_n N_X_c_626_n 0.00354304f $X=3.565 $Y=1.4 $X2=0 $Y2=0
cc_281 N_A_c_352_n N_VGND_c_700_n 0.00474653f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A_c_352_n N_VGND_c_712_n 0.00428022f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A_c_352_n N_VGND_c_715_n 0.00622134f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A_335_297#_c_398_n N_VPWR_c_540_n 0.0100747f $X=4.075 $Y=1.41 $X2=0
+ $Y2=0
cc_285 N_A_335_297#_c_396_n N_VPWR_c_540_n 0.00249053f $X=4.015 $Y=1.16 $X2=0
+ $Y2=0
cc_286 N_A_335_297#_c_399_n N_VPWR_c_541_n 0.00300743f $X=4.545 $Y=1.41 $X2=0
+ $Y2=0
cc_287 N_A_335_297#_c_400_n N_VPWR_c_541_n 0.00300743f $X=5.015 $Y=1.41 $X2=0
+ $Y2=0
cc_288 N_A_335_297#_c_401_n N_VPWR_c_543_n 0.00479105f $X=5.485 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_335_297#_c_398_n N_VPWR_c_546_n 0.00702461f $X=4.075 $Y=1.41 $X2=0
+ $Y2=0
cc_290 N_A_335_297#_c_399_n N_VPWR_c_546_n 0.00702461f $X=4.545 $Y=1.41 $X2=0
+ $Y2=0
cc_291 N_A_335_297#_c_400_n N_VPWR_c_549_n 0.00702461f $X=5.015 $Y=1.41 $X2=0
+ $Y2=0
cc_292 N_A_335_297#_c_401_n N_VPWR_c_549_n 0.00702461f $X=5.485 $Y=1.41 $X2=0
+ $Y2=0
cc_293 N_A_335_297#_M1001_s N_VPWR_c_538_n 0.00218346f $X=1.675 $Y=1.485 $X2=0
+ $Y2=0
cc_294 N_A_335_297#_c_398_n N_VPWR_c_538_n 0.012878f $X=4.075 $Y=1.41 $X2=0
+ $Y2=0
cc_295 N_A_335_297#_c_399_n N_VPWR_c_538_n 0.0124092f $X=4.545 $Y=1.41 $X2=0
+ $Y2=0
cc_296 N_A_335_297#_c_400_n N_VPWR_c_538_n 0.0124092f $X=5.015 $Y=1.41 $X2=0
+ $Y2=0
cc_297 N_A_335_297#_c_401_n N_VPWR_c_538_n 0.0133206f $X=5.485 $Y=1.41 $X2=0
+ $Y2=0
cc_298 N_A_335_297#_c_402_n A_425_297# 0.00194751f $X=2.035 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_335_297#_c_394_n A_425_297# 0.00405738f $X=2.13 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_300 N_A_335_297#_c_398_n N_X_c_626_n 4.56612e-19 $X=4.075 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A_335_297#_c_471_p N_X_c_626_n 0.0172229f $X=5.28 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_335_297#_c_397_n N_X_c_626_n 0.00674235f $X=5.485 $Y=1.202 $X2=0
+ $Y2=0
cc_303 N_A_335_297#_c_390_n N_X_c_635_n 0.00488834f $X=4.05 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A_335_297#_c_391_n N_X_c_635_n 0.00766092f $X=4.52 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A_335_297#_c_392_n N_X_c_635_n 5.47877e-19 $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A_335_297#_c_442_n N_X_c_635_n 0.00476601f $X=3.845 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A_335_297#_c_399_n N_X_c_627_n 0.0158555f $X=4.545 $Y=1.41 $X2=0 $Y2=0
cc_308 N_A_335_297#_c_400_n N_X_c_627_n 0.0159162f $X=5.015 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_335_297#_c_471_p N_X_c_627_n 0.0406907f $X=5.28 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A_335_297#_c_397_n N_X_c_627_n 0.00881912f $X=5.485 $Y=1.202 $X2=0
+ $Y2=0
cc_311 N_A_335_297#_c_391_n N_X_c_620_n 0.00901745f $X=4.52 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_335_297#_c_392_n N_X_c_620_n 0.00895898f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A_335_297#_c_471_p N_X_c_620_n 0.0392656f $X=5.28 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_335_297#_c_397_n N_X_c_620_n 0.00345541f $X=5.485 $Y=1.202 $X2=0
+ $Y2=0
cc_315 N_A_335_297#_c_390_n N_X_c_621_n 0.00154411f $X=4.05 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A_335_297#_c_391_n N_X_c_621_n 0.00270583f $X=4.52 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A_335_297#_c_442_n N_X_c_621_n 0.00741575f $X=3.845 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_335_297#_c_395_n N_X_c_621_n 0.00537347f $X=3.93 $Y=1.075 $X2=0 $Y2=0
cc_319 N_A_335_297#_c_471_p N_X_c_621_n 0.0199589f $X=5.28 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_335_297#_c_397_n N_X_c_621_n 0.0033272f $X=5.485 $Y=1.202 $X2=0 $Y2=0
cc_321 N_A_335_297#_c_391_n N_X_c_653_n 5.24597e-19 $X=4.52 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A_335_297#_c_392_n N_X_c_653_n 0.00651696f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A_335_297#_c_401_n N_X_c_628_n 0.0184873f $X=5.485 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A_335_297#_c_471_p N_X_c_628_n 0.00405064f $X=5.28 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_335_297#_c_397_n N_X_c_628_n 9.44246e-19 $X=5.485 $Y=1.202 $X2=0
+ $Y2=0
cc_326 N_A_335_297#_c_393_n N_X_c_622_n 0.0137132f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_335_297#_c_471_p N_X_c_622_n 0.00208021f $X=5.28 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_335_297#_c_392_n N_X_c_623_n 0.00119564f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A_335_297#_c_471_p N_X_c_623_n 0.0304076f $X=5.28 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A_335_297#_c_397_n N_X_c_623_n 0.00486271f $X=5.485 $Y=1.202 $X2=0
+ $Y2=0
cc_331 N_A_335_297#_c_471_p N_X_c_629_n 0.0172229f $X=5.28 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A_335_297#_c_397_n N_X_c_629_n 0.0065364f $X=5.485 $Y=1.202 $X2=0 $Y2=0
cc_333 N_A_335_297#_c_401_n X 0.00181588f $X=5.485 $Y=1.41 $X2=0 $Y2=0
cc_334 N_A_335_297#_c_393_n X 0.0204329f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A_335_297#_c_471_p X 0.0131388f $X=5.28 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_335_297#_c_432_n N_VGND_M1012_d 0.0075965f $X=3.185 $Y=0.74 $X2=0
+ $Y2=0
cc_337 N_A_335_297#_c_442_n N_VGND_M1002_d 0.00924952f $X=3.845 $Y=0.74 $X2=0
+ $Y2=0
cc_338 N_A_335_297#_c_395_n N_VGND_M1002_d 7.52091e-19 $X=3.93 $Y=1.075 $X2=0
+ $Y2=0
cc_339 N_A_335_297#_c_419_n N_VGND_c_699_n 0.013438f $X=2.33 $Y=0.49 $X2=0 $Y2=0
cc_340 N_A_335_297#_c_432_n N_VGND_c_699_n 0.0214497f $X=3.185 $Y=0.74 $X2=0
+ $Y2=0
cc_341 N_A_335_297#_c_390_n N_VGND_c_700_n 0.00814668f $X=4.05 $Y=0.995 $X2=0
+ $Y2=0
cc_342 N_A_335_297#_c_391_n N_VGND_c_700_n 0.00115121f $X=4.52 $Y=0.995 $X2=0
+ $Y2=0
cc_343 N_A_335_297#_c_442_n N_VGND_c_700_n 0.0251303f $X=3.845 $Y=0.74 $X2=0
+ $Y2=0
cc_344 N_A_335_297#_c_391_n N_VGND_c_701_n 0.00379224f $X=4.52 $Y=0.995 $X2=0
+ $Y2=0
cc_345 N_A_335_297#_c_392_n N_VGND_c_701_n 0.00276126f $X=4.99 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_A_335_297#_c_393_n N_VGND_c_703_n 0.00438629f $X=5.51 $Y=0.995 $X2=0
+ $Y2=0
cc_347 N_A_335_297#_c_419_n N_VGND_c_708_n 0.00852533f $X=2.33 $Y=0.49 $X2=0
+ $Y2=0
cc_348 N_A_335_297#_c_420_n N_VGND_c_708_n 0.00535673f $X=2.415 $Y=0.74 $X2=0
+ $Y2=0
cc_349 N_A_335_297#_c_390_n N_VGND_c_710_n 0.00485605f $X=4.05 $Y=0.995 $X2=0
+ $Y2=0
cc_350 N_A_335_297#_c_391_n N_VGND_c_710_n 0.00423334f $X=4.52 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_335_297#_c_442_n N_VGND_c_710_n 3.30713e-19 $X=3.845 $Y=0.74 $X2=0
+ $Y2=0
cc_352 N_A_335_297#_c_432_n N_VGND_c_712_n 0.0029785f $X=3.185 $Y=0.74 $X2=0
+ $Y2=0
cc_353 N_A_335_297#_c_523_p N_VGND_c_712_n 0.00846569f $X=3.27 $Y=0.49 $X2=0
+ $Y2=0
cc_354 N_A_335_297#_c_442_n N_VGND_c_712_n 0.00337235f $X=3.845 $Y=0.74 $X2=0
+ $Y2=0
cc_355 N_A_335_297#_c_392_n N_VGND_c_713_n 0.00423334f $X=4.99 $Y=0.995 $X2=0
+ $Y2=0
cc_356 N_A_335_297#_c_393_n N_VGND_c_713_n 0.00437852f $X=5.51 $Y=0.995 $X2=0
+ $Y2=0
cc_357 N_A_335_297#_M1011_d N_VGND_c_715_n 0.00417844f $X=2.115 $Y=0.235 $X2=0
+ $Y2=0
cc_358 N_A_335_297#_M1005_d N_VGND_c_715_n 0.00256656f $X=3.135 $Y=0.235 $X2=0
+ $Y2=0
cc_359 N_A_335_297#_c_390_n N_VGND_c_715_n 0.00802939f $X=4.05 $Y=0.995 $X2=0
+ $Y2=0
cc_360 N_A_335_297#_c_391_n N_VGND_c_715_n 0.00613677f $X=4.52 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A_335_297#_c_392_n N_VGND_c_715_n 0.00608558f $X=4.99 $Y=0.995 $X2=0
+ $Y2=0
cc_362 N_A_335_297#_c_393_n N_VGND_c_715_n 0.00708323f $X=5.51 $Y=0.995 $X2=0
+ $Y2=0
cc_363 N_A_335_297#_c_419_n N_VGND_c_715_n 0.00618681f $X=2.33 $Y=0.49 $X2=0
+ $Y2=0
cc_364 N_A_335_297#_c_432_n N_VGND_c_715_n 0.00691826f $X=3.185 $Y=0.74 $X2=0
+ $Y2=0
cc_365 N_A_335_297#_c_420_n N_VGND_c_715_n 0.00992647f $X=2.415 $Y=0.74 $X2=0
+ $Y2=0
cc_366 N_A_335_297#_c_523_p N_VGND_c_715_n 0.00625722f $X=3.27 $Y=0.49 $X2=0
+ $Y2=0
cc_367 N_A_335_297#_c_442_n N_VGND_c_715_n 0.00873958f $X=3.845 $Y=0.74 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_538_n A_425_297# 0.00281072f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_369 N_VPWR_c_538_n A_531_297# 0.00899181f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_370 N_VPWR_c_538_n A_625_297# 0.0117429f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_371 N_VPWR_c_538_n N_X_M1000_d 0.00370124f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_372 N_VPWR_c_538_n N_X_M1016_d 0.00370124f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_373 N_VPWR_c_546_n N_X_c_670_n 0.0149311f $X=4.655 $Y=2.72 $X2=0 $Y2=0
cc_374 N_VPWR_c_538_n N_X_c_670_n 0.00955092f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_375 N_VPWR_M1007_s N_X_c_627_n 0.00187091f $X=4.635 $Y=1.485 $X2=0 $Y2=0
cc_376 N_VPWR_c_541_n N_X_c_627_n 0.0143191f $X=4.78 $Y=1.96 $X2=0 $Y2=0
cc_377 N_VPWR_c_549_n N_X_c_674_n 0.0149311f $X=5.595 $Y=2.72 $X2=0 $Y2=0
cc_378 N_VPWR_c_538_n N_X_c_674_n 0.00955092f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_379 N_VPWR_M1018_s N_X_c_628_n 0.00304346f $X=5.575 $Y=1.485 $X2=0 $Y2=0
cc_380 N_VPWR_c_543_n N_X_c_628_n 0.0191143f $X=5.72 $Y=1.96 $X2=0 $Y2=0
cc_381 N_X_c_620_n N_VGND_M1013_s 0.00251047f $X=5.035 $Y=0.815 $X2=0 $Y2=0
cc_382 N_X_c_625_n N_VGND_M1019_s 0.00326313f $X=5.74 $Y=0.905 $X2=0 $Y2=0
cc_383 N_X_c_635_n N_VGND_c_700_n 0.0140037f $X=4.31 $Y=0.485 $X2=0 $Y2=0
cc_384 N_X_c_635_n N_VGND_c_701_n 0.0177813f $X=4.31 $Y=0.485 $X2=0 $Y2=0
cc_385 N_X_c_620_n N_VGND_c_701_n 0.0127273f $X=5.035 $Y=0.815 $X2=0 $Y2=0
cc_386 N_X_c_625_n N_VGND_c_702_n 8.14798e-19 $X=5.74 $Y=0.905 $X2=0 $Y2=0
cc_387 N_X_c_625_n N_VGND_c_703_n 0.0140097f $X=5.74 $Y=0.905 $X2=0 $Y2=0
cc_388 N_X_c_635_n N_VGND_c_710_n 0.0153475f $X=4.31 $Y=0.485 $X2=0 $Y2=0
cc_389 N_X_c_620_n N_VGND_c_710_n 0.00266636f $X=5.035 $Y=0.815 $X2=0 $Y2=0
cc_390 N_X_c_620_n N_VGND_c_713_n 0.00198695f $X=5.035 $Y=0.815 $X2=0 $Y2=0
cc_391 N_X_c_653_n N_VGND_c_713_n 0.0231806f $X=5.25 $Y=0.39 $X2=0 $Y2=0
cc_392 N_X_c_622_n N_VGND_c_713_n 0.00247541f $X=5.625 $Y=0.815 $X2=0 $Y2=0
cc_393 N_X_M1006_d N_VGND_c_715_n 0.00607585f $X=4.125 $Y=0.235 $X2=0 $Y2=0
cc_394 N_X_M1015_d N_VGND_c_715_n 0.00304143f $X=5.065 $Y=0.235 $X2=0 $Y2=0
cc_395 N_X_c_635_n N_VGND_c_715_n 0.00940698f $X=4.31 $Y=0.485 $X2=0 $Y2=0
cc_396 N_X_c_620_n N_VGND_c_715_n 0.00972452f $X=5.035 $Y=0.815 $X2=0 $Y2=0
cc_397 N_X_c_653_n N_VGND_c_715_n 0.0143352f $X=5.25 $Y=0.39 $X2=0 $Y2=0
cc_398 N_X_c_622_n N_VGND_c_715_n 0.00471693f $X=5.625 $Y=0.815 $X2=0 $Y2=0
cc_399 N_X_c_625_n N_VGND_c_715_n 0.0024595f $X=5.74 $Y=0.905 $X2=0 $Y2=0
