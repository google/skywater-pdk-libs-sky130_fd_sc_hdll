# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o22ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o22ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 1.565000 1.275000 ;
        RECT 1.250000 1.275000 1.565000 1.445000 ;
        RECT 1.250000 1.445000 4.030000 1.615000 ;
        RECT 3.625000 1.075000 4.030000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.835000 1.075000 3.445000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745000 0.995000 5.490000 1.445000 ;
        RECT 4.745000 1.445000 7.735000 1.615000 ;
        RECT 7.465000 0.995000 7.735000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.660000 1.075000 7.160000 1.275000 ;
    END
  END B2
  PIN VGND
    ANTENNADIFFAREA  0.799500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  1.490000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.959500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 1.785000 4.370000 1.955000 ;
        RECT 1.955000 1.955000 2.295000 2.125000 ;
        RECT 2.985000 1.955000 3.235000 2.125000 ;
        RECT 4.200000 1.445000 4.575000 1.615000 ;
        RECT 4.200000 1.615000 4.370000 1.785000 ;
        RECT 4.355000 0.645000 8.170000 0.820000 ;
        RECT 4.355000 0.820000 4.575000 1.445000 ;
        RECT 5.855000 1.785000 8.170000 1.955000 ;
        RECT 5.855000 1.955000 6.105000 2.125000 ;
        RECT 6.795000 1.955000 7.045000 2.125000 ;
        RECT 7.905000 0.820000 8.170000 1.785000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.125000  0.255000 0.455000 0.725000 ;
      RECT 0.125000  0.725000 1.395000 0.735000 ;
      RECT 0.125000  0.735000 4.185000 0.905000 ;
      RECT 0.165000  1.445000 0.415000 2.635000 ;
      RECT 0.635000  1.445000 0.885000 1.785000 ;
      RECT 0.635000  1.785000 1.785000 1.955000 ;
      RECT 0.635000  1.955000 0.885000 2.465000 ;
      RECT 0.675000  0.085000 0.845000 0.555000 ;
      RECT 1.015000  0.255000 1.395000 0.725000 ;
      RECT 1.105000  2.125000 1.355000 2.635000 ;
      RECT 1.575000  1.955000 1.785000 2.295000 ;
      RECT 1.575000  2.295000 3.745000 2.465000 ;
      RECT 1.615000  0.085000 1.785000 0.555000 ;
      RECT 1.955000  0.255000 2.335000 0.725000 ;
      RECT 1.955000  0.725000 3.275000 0.735000 ;
      RECT 2.515000  2.125000 2.765000 2.295000 ;
      RECT 2.555000  0.085000 2.725000 0.555000 ;
      RECT 2.895000  0.255000 3.275000 0.725000 ;
      RECT 3.455000  2.125000 3.745000 2.295000 ;
      RECT 3.495000  0.085000 3.665000 0.555000 ;
      RECT 3.835000  0.255000 8.045000 0.475000 ;
      RECT 3.835000  0.475000 4.185000 0.735000 ;
      RECT 3.965000  2.125000 4.185000 2.635000 ;
      RECT 4.355000  2.125000 4.710000 2.465000 ;
      RECT 4.540000  1.785000 5.635000 1.955000 ;
      RECT 4.540000  1.955000 4.710000 2.125000 ;
      RECT 4.925000  2.125000 5.165000 2.635000 ;
      RECT 5.385000  1.955000 5.635000 2.295000 ;
      RECT 5.385000  2.295000 7.515000 2.465000 ;
      RECT 6.325000  2.125000 6.575000 2.295000 ;
      RECT 7.265000  2.135000 7.515000 2.295000 ;
      RECT 7.735000  2.125000 8.015000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22ai_4
END LIBRARY
