* File: sky130_fd_sc_hdll__a32o_4.pex.spice
* Created: Thu Aug 27 18:56:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A32O_4%A_79_21# 1 2 3 4 13 15 16 18 19 21 22 24 25
+ 27 28 30 31 33 34 36 37 46 47 48 49 54 56 58 63 67 69 70 71 80
c179 80 0 1.75139e-19 $X=1.905 $Y=1.202
c180 46 0 1.04313e-19 $X=2.06 $Y=1.495
r181 80 81 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r182 77 78 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r183 76 77 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.41 $Y2=1.202
r184 75 76 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r185 72 73 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r186 70 71 4.00505 $w=1.78e-07 $l=6.5e-08 $layer=LI1_cond $X=6.445 $Y=1.995
+ $X2=6.51 $Y2=1.995
r187 65 67 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.865 $Y=0.72
+ $X2=6.565 $Y2=0.72
r188 61 63 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.61 $Y=2 $X2=7.55
+ $Y2=2
r189 61 71 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.61 $Y=2 $X2=6.51
+ $Y2=2
r190 58 70 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.95 $Y=1.99
+ $X2=6.445 $Y2=1.99
r191 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.865 $Y=1.905
+ $X2=5.95 $Y2=1.99
r192 55 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.865 $Y=1.665
+ $X2=5.865 $Y2=1.58
r193 55 56 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.865 $Y=1.665
+ $X2=5.865 $Y2=1.905
r194 54 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.865 $Y=1.495
+ $X2=5.865 $Y2=1.58
r195 53 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.865 $Y=0.805
+ $X2=5.865 $Y2=0.72
r196 53 54 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.865 $Y=0.805
+ $X2=5.865 $Y2=1.495
r197 49 65 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.78 $Y=0.72
+ $X2=5.865 $Y2=0.72
r198 49 51 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.78 $Y=0.72
+ $X2=5.01 $Y2=0.72
r199 47 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.78 $Y=1.58
+ $X2=5.865 $Y2=1.58
r200 47 48 235.519 $w=1.68e-07 $l=3.61e-06 $layer=LI1_cond $X=5.78 $Y=1.58
+ $X2=2.17 $Y2=1.58
r201 46 48 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.06 $Y=1.495
+ $X2=2.17 $Y2=1.58
r202 45 46 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=2.06 $Y=1.325
+ $X2=2.06 $Y2=1.495
r203 44 80 53.1237 $w=3.72e-07 $l=4.1e-07 $layer=POLY_cond $X=1.495 $Y=1.202
+ $X2=1.905 $Y2=1.202
r204 44 78 7.77419 $w=3.72e-07 $l=6e-08 $layer=POLY_cond $X=1.495 $Y=1.202
+ $X2=1.435 $Y2=1.202
r205 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=1.16 $X2=1.495 $Y2=1.16
r206 40 75 30.4489 $w=3.72e-07 $l=2.35e-07 $layer=POLY_cond $X=0.705 $Y=1.202
+ $X2=0.94 $Y2=1.202
r207 40 73 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=0.705 $Y=1.202
+ $X2=0.495 $Y2=1.202
r208 39 43 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.705 $Y=1.16
+ $X2=1.495 $Y2=1.16
r209 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.705
+ $Y=1.16 $X2=0.705 $Y2=1.16
r210 37 45 7.17723 $w=3.3e-07 $l=2.13014e-07 $layer=LI1_cond $X=1.95 $Y=1.16
+ $X2=2.06 $Y2=1.325
r211 37 43 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.95 $Y=1.16
+ $X2=1.495 $Y2=1.16
r212 34 81 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r213 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r214 31 80 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r215 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r216 28 78 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r217 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r218 25 77 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r219 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r220 22 76 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r221 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r222 19 75 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r223 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r224 16 73 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r225 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r226 13 72 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r227 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r228 4 63 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=7.405
+ $Y=1.485 $X2=7.55 $Y2=2
r229 3 61 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=6.465
+ $Y=1.485 $X2=6.61 $Y2=2
r230 2 67 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.43
+ $Y=0.235 $X2=6.565 $Y2=0.72
r231 1 51 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.235 $X2=5.01 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%A3 1 3 4 6 7 9 10 12 13 14 20 25 29
c50 14 0 1.75139e-19 $X=2.915 $Y=1.105
r51 22 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.965
+ $Y=1.16 $X2=2.965 $Y2=1.16
r52 20 22 16.0222 $w=3.61e-07 $l=1.2e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=2.965 $Y2=1.202
r53 19 20 3.33795 $w=3.61e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r54 18 19 59.4155 $w=3.61e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.82 $Y2=1.202
r55 17 18 3.33795 $w=3.61e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r56 14 29 1.83343 $w=2.18e-07 $l=3.5e-08 $layer=LI1_cond $X=3 $Y=1.185 $X2=2.965
+ $Y2=1.185
r57 13 29 22.2631 $w=2.18e-07 $l=4.25e-07 $layer=LI1_cond $X=2.54 $Y=1.185
+ $X2=2.965 $Y2=1.185
r58 13 25 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=2.54 $Y=1.185
+ $X2=2.535 $Y2=1.185
r59 10 20 19.0337 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r60 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r61 7 19 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r62 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995 $X2=2.82
+ $Y2=0.56
r63 4 18 19.0337 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r64 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r65 1 17 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r66 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995 $X2=2.35
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%A2 1 3 4 6 7 9 10 12 13 23 28
r46 23 24 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.33 $Y2=1.202
r47 21 23 14.9407 $w=3.71e-07 $l=1.15e-07 $layer=POLY_cond $X=4.19 $Y=1.202
+ $X2=4.305 $Y2=1.202
r48 19 21 42.8733 $w=3.71e-07 $l=3.3e-07 $layer=POLY_cond $X=3.86 $Y=1.202
+ $X2=4.19 $Y2=1.202
r49 18 19 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=3.835 $Y=1.202
+ $X2=3.86 $Y2=1.202
r50 17 28 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=3.8 $Y=1.2
+ $X2=4.115 $Y2=1.2
r51 16 18 4.54717 $w=3.71e-07 $l=3.5e-08 $layer=POLY_cond $X=3.8 $Y=1.202
+ $X2=3.835 $Y2=1.202
r52 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.8
+ $Y=1.16 $X2=3.8 $Y2=1.16
r53 13 28 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.12 $Y=1.2 $X2=4.115
+ $Y2=1.2
r54 13 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.19
+ $Y=1.16 $X2=4.19 $Y2=1.16
r55 10 24 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.33 $Y=0.995
+ $X2=4.33 $Y2=1.202
r56 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.33 $Y=0.995
+ $X2=4.33 $Y2=0.56
r57 7 23 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r58 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r59 4 19 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=1.202
r60 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995 $X2=3.86
+ $Y2=0.56
r61 1 18 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.202
r62 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%A1 3 5 7 10 12 14 15 16 25 32 36
c48 25 0 9.29584e-20 $X=5.245 $Y=1.212
r49 27 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.36
+ $Y=1.16 $X2=5.36 $Y2=1.16
r50 25 27 16.1604 $w=3.43e-07 $l=1.15e-07 $layer=POLY_cond $X=5.245 $Y=1.212
+ $X2=5.36 $Y2=1.212
r51 24 25 3.51312 $w=3.43e-07 $l=2.5e-08 $layer=POLY_cond $X=5.22 $Y=1.212
+ $X2=5.245 $Y2=1.212
r52 23 32 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.02 $Y=1.2
+ $X2=4.855 $Y2=1.2
r53 22 24 28.105 $w=3.43e-07 $l=2e-07 $layer=POLY_cond $X=5.02 $Y=1.212 $X2=5.22
+ $Y2=1.212
r54 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.02
+ $Y=1.16 $X2=5.02 $Y2=1.16
r55 20 22 34.4286 $w=3.43e-07 $l=2.45e-07 $layer=POLY_cond $X=4.775 $Y=1.212
+ $X2=5.02 $Y2=1.212
r56 19 20 3.51312 $w=3.43e-07 $l=2.5e-08 $layer=POLY_cond $X=4.75 $Y=1.212
+ $X2=4.775 $Y2=1.212
r57 16 36 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=5.305 $Y=1.2 $X2=5.345
+ $Y2=1.2
r58 16 23 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=5.305 $Y=1.2
+ $X2=5.02 $Y2=1.2
r59 15 32 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=4.835 $Y=1.2
+ $X2=4.855 $Y2=1.2
r60 12 25 17.8339 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.212
r61 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r62 8 24 22.1447 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=5.22 $Y=1.015
+ $X2=5.22 $Y2=1.212
r63 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.22 $Y=1.015
+ $X2=5.22 $Y2=0.56
r64 5 20 17.8339 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.212
r65 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r66 1 19 22.1447 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=1.212
r67 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%B1 3 5 7 10 12 14 15 17 31 36 39 44
c53 31 0 1.76016e-19 $X=6.825 $Y=1.217
c54 3 0 9.29584e-20 $X=6.355 $Y=0.56
r55 36 39 0.0217469 $w=5.48e-07 $l=1e-09 $layer=LI1_cond $X=6.534 $Y=1.35
+ $X2=6.535 $Y2=1.35
r56 31 32 2.83529 $w=3.4e-07 $l=2e-08 $layer=POLY_cond $X=6.825 $Y=1.217
+ $X2=6.845 $Y2=1.217
r57 30 44 5.76292 $w=5.48e-07 $l=2.65e-07 $layer=LI1_cond $X=6.73 $Y=1.35
+ $X2=6.995 $Y2=1.35
r58 29 31 13.4676 $w=3.4e-07 $l=9.5e-08 $layer=POLY_cond $X=6.73 $Y=1.217
+ $X2=6.825 $Y2=1.217
r59 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.73
+ $Y=1.16 $X2=6.73 $Y2=1.16
r60 27 29 50.3265 $w=3.4e-07 $l=3.55e-07 $layer=POLY_cond $X=6.375 $Y=1.217
+ $X2=6.73 $Y2=1.217
r61 26 27 2.83529 $w=3.4e-07 $l=2e-08 $layer=POLY_cond $X=6.355 $Y=1.217
+ $X2=6.375 $Y2=1.217
r62 25 36 4.21889 $w=5.48e-07 $l=1.94e-07 $layer=LI1_cond $X=6.34 $Y=1.35
+ $X2=6.534 $Y2=1.35
r63 24 26 2.12647 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=6.34 $Y=1.217
+ $X2=6.355 $Y2=1.217
r64 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.34
+ $Y=1.16 $X2=6.34 $Y2=1.16
r65 17 44 1.19608 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=7.05 $Y=1.35
+ $X2=6.995 $Y2=1.35
r66 15 30 2.28342 $w=5.48e-07 $l=1.05e-07 $layer=LI1_cond $X=6.625 $Y=1.35
+ $X2=6.73 $Y2=1.35
r67 15 39 1.95722 $w=5.48e-07 $l=9e-08 $layer=LI1_cond $X=6.625 $Y=1.35
+ $X2=6.535 $Y2=1.35
r68 12 32 17.6285 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.845 $Y=1.41
+ $X2=6.845 $Y2=1.217
r69 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.845 $Y=1.41
+ $X2=6.845 $Y2=1.985
r70 8 31 21.9347 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.825 $Y=1.025
+ $X2=6.825 $Y2=1.217
r71 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.825 $Y=1.025
+ $X2=6.825 $Y2=0.56
r72 5 27 17.6285 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.375 $Y=1.41
+ $X2=6.375 $Y2=1.217
r73 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.375 $Y=1.41
+ $X2=6.375 $Y2=1.985
r74 1 26 21.9347 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.355 $Y=1.025
+ $X2=6.355 $Y2=1.217
r75 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.355 $Y=1.025
+ $X2=6.355 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%B2 3 5 7 10 12 14 15 20 21 22 27 30 36
c45 30 0 1.54818e-19 $X=7.537 $Y=1.295
c46 21 0 2.11977e-20 $X=7.525 $Y=1.53
r47 34 36 14.6675 $w=2.18e-07 $l=2.8e-07 $layer=LI1_cond $X=7.635 $Y=1.185
+ $X2=7.915 $Y2=1.185
r48 22 36 4.71454 $w=2.18e-07 $l=9e-08 $layer=LI1_cond $X=8.005 $Y=1.185
+ $X2=7.915 $Y2=1.185
r49 22 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.005
+ $Y=1.16 $X2=8.005 $Y2=1.16
r50 21 30 13.366 $w=1.93e-07 $l=2.35e-07 $layer=LI1_cond $X=7.537 $Y=1.53
+ $X2=7.537 $Y2=1.295
r51 20 30 3.62192 $w=1.95e-07 $l=1.1e-07 $layer=LI1_cond $X=7.537 $Y=1.185
+ $X2=7.537 $Y2=1.295
r52 20 34 3.2268 $w=2.2e-07 $l=9.8e-08 $layer=LI1_cond $X=7.537 $Y=1.185
+ $X2=7.635 $Y2=1.185
r53 18 19 3.44286 $w=3.5e-07 $l=2.5e-08 $layer=POLY_cond $X=7.76 $Y=1.217
+ $X2=7.785 $Y2=1.217
r54 17 18 61.2829 $w=3.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.315 $Y=1.217
+ $X2=7.76 $Y2=1.217
r55 16 17 3.44286 $w=3.5e-07 $l=2.5e-08 $layer=POLY_cond $X=7.29 $Y=1.217
+ $X2=7.315 $Y2=1.217
r56 15 27 25.7087 $w=2.8e-07 $l=1.2e-07 $layer=POLY_cond $X=7.885 $Y=1.165
+ $X2=8.005 $Y2=1.165
r57 15 19 15.8382 $w=3.5e-07 $l=1.23288e-07 $layer=POLY_cond $X=7.885 $Y=1.165
+ $X2=7.785 $Y2=1.217
r58 12 19 18.307 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.785 $Y=1.41
+ $X2=7.785 $Y2=1.217
r59 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.785 $Y=1.41
+ $X2=7.785 $Y2=1.985
r60 8 18 22.6286 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.76 $Y=1.025
+ $X2=7.76 $Y2=1.217
r61 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.76 $Y=1.025
+ $X2=7.76 $Y2=0.56
r62 5 17 18.307 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.315 $Y=1.41
+ $X2=7.315 $Y2=1.217
r63 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.315 $Y=1.41
+ $X2=7.315 $Y2=1.985
r64 1 16 22.6286 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.29 $Y=1.025
+ $X2=7.29 $Y2=1.217
r65 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.29 $Y=1.025
+ $X2=7.29 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%VPWR 1 2 3 4 5 6 19 21 25 29 31 33 35 37 42
+ 47 57 58 64 67 70 77 84
c131 3 0 1.04313e-19 $X=1.995 $Y=1.485
c132 1 0 1.47114e-19 $X=0.135 $Y=1.485
r133 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r134 84 87 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=4.985 $Y=2.34
+ $X2=4.985 $Y2=2.72
r135 81 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r136 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r137 77 80 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=4.045 $Y=2.34
+ $X2=4.045 $Y2=2.72
r138 74 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r139 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r140 70 73 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.055 $Y=2.34
+ $X2=3.055 $Y2=2.72
r141 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r142 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 57 58 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r144 55 58 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=8.05 $Y2=2.72
r145 55 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r146 54 57 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=8.05 $Y2=2.72
r147 54 55 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r148 52 87 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=2.72
+ $X2=4.985 $Y2=2.72
r149 52 54 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.175 $Y=2.72
+ $X2=5.29 $Y2=2.72
r150 51 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r151 51 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r152 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r153 48 67 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.305 $Y=2.72
+ $X2=2.115 $Y2=2.72
r154 48 50 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.305 $Y=2.72
+ $X2=2.53 $Y2=2.72
r155 47 73 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.055 $Y2=2.72
r156 47 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.53 $Y2=2.72
r157 46 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r158 46 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r159 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r160 43 64 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.175 $Y2=2.72
r161 43 45 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.61 $Y2=2.72
r162 42 67 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.925 $Y=2.72
+ $X2=2.115 $Y2=2.72
r163 42 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.925 $Y=2.72
+ $X2=1.61 $Y2=2.72
r164 41 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r165 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r166 38 61 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r167 38 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r168 37 64 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=1.175 $Y2=2.72
r169 37 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=0.69 $Y2=2.72
r170 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r171 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r172 34 80 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.235 $Y=2.72
+ $X2=4.045 $Y2=2.72
r173 33 87 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.985 $Y2=2.72
r174 33 34 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.235 $Y2=2.72
r175 32 73 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.055 $Y2=2.72
r176 31 80 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=4.045 $Y2=2.72
r177 31 32 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=3.245 $Y2=2.72
r178 27 67 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=2.635
+ $X2=2.115 $Y2=2.72
r179 27 29 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.115 $Y=2.635
+ $X2=2.115 $Y2=2
r180 23 64 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=2.635
+ $X2=1.175 $Y2=2.72
r181 23 25 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=1.175 $Y=2.635
+ $X2=1.175 $Y2=2
r182 19 61 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r183 19 21 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2
r184 6 84 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.34
r185 5 77 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.34
r186 4 70 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2.34
r187 3 29 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r188 2 25 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r189 1 21 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%X 1 2 3 4 13 15 19 23 25 27 31 35 37 38 39
+ 40 41 47 48 50
c70 50 0 1.47114e-19 $X=0.235 $Y=0.85
r71 47 50 2.35727 $w=2.18e-07 $l=4.5e-08 $layer=LI1_cond $X=0.23 $Y=0.805
+ $X2=0.23 $Y2=0.85
r72 41 48 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=1.58 $X2=0.23
+ $Y2=1.495
r73 41 48 1.30959 $w=2.18e-07 $l=2.5e-08 $layer=LI1_cond $X=0.23 $Y=1.47
+ $X2=0.23 $Y2=1.495
r74 40 41 14.6675 $w=2.18e-07 $l=2.8e-07 $layer=LI1_cond $X=0.23 $Y=1.19
+ $X2=0.23 $Y2=1.47
r75 39 47 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=0.72 $X2=0.23
+ $Y2=0.805
r76 39 40 16.7628 $w=2.18e-07 $l=3.2e-07 $layer=LI1_cond $X=0.23 $Y=0.87
+ $X2=0.23 $Y2=1.19
r77 39 50 1.04768 $w=2.18e-07 $l=2e-08 $layer=LI1_cond $X=0.23 $Y=0.87 $X2=0.23
+ $Y2=0.85
r78 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.96
r79 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.67 $Y=0.635
+ $X2=1.67 $Y2=0.42
r80 28 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=1.58
+ $X2=0.73 $Y2=1.58
r81 27 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.585 $Y=1.58
+ $X2=1.67 $Y2=1.665
r82 27 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=1.58
+ $X2=0.815 $Y2=1.58
r83 26 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.72
+ $X2=0.73 $Y2=0.72
r84 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.585 $Y=0.72
+ $X2=1.67 $Y2=0.635
r85 25 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0.72
+ $X2=0.815 $Y2=0.72
r86 21 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.58
r87 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.96
r88 17 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.635
+ $X2=0.73 $Y2=0.72
r89 17 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.73 $Y=0.635
+ $X2=0.73 $Y2=0.42
r90 16 41 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.34 $Y=1.58 $X2=0.23
+ $Y2=1.58
r91 15 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.645 $Y=1.58
+ $X2=0.73 $Y2=1.58
r92 15 16 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.645 $Y=1.58
+ $X2=0.34 $Y2=1.58
r93 14 39 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.34 $Y=0.72 $X2=0.23
+ $Y2=0.72
r94 13 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.645 $Y=0.72
+ $X2=0.73 $Y2=0.72
r95 13 14 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.645 $Y=0.72
+ $X2=0.34 $Y2=0.72
r96 4 35 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.96
r97 3 23 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
r98 2 31 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.42
r99 1 19 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%A_493_297# 1 2 3 4 5 6 21 23 24 27 29 33 35
+ 38 39 40 45 47 49 50
r91 45 52 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.06 $Y=2.255
+ $X2=8.06 $Y2=2.34
r92 45 47 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.06 $Y=2.255
+ $X2=8.06 $Y2=1.92
r93 42 44 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.14 $Y=2.34
+ $X2=7.08 $Y2=2.34
r94 40 42 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.565 $Y=2.34
+ $X2=6.14 $Y2=2.34
r95 39 52 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.935 $Y=2.34
+ $X2=8.06 $Y2=2.34
r96 39 44 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=7.935 $Y=2.34
+ $X2=7.08 $Y2=2.34
r97 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.48 $Y=2.255
+ $X2=5.565 $Y2=2.34
r98 37 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.48 $Y=2.085
+ $X2=5.48 $Y2=2.255
r99 36 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=2 $X2=4.54
+ $Y2=2
r100 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.395 $Y=2
+ $X2=5.48 $Y2=2.085
r101 35 36 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.395 $Y=2
+ $X2=4.625 $Y2=2
r102 31 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.085
+ $X2=4.54 $Y2=2
r103 31 33 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.54 $Y=2.085
+ $X2=4.54 $Y2=2.3
r104 30 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=2 $X2=3.6
+ $Y2=2
r105 29 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=2 $X2=4.54
+ $Y2=2
r106 29 30 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.455 $Y=2
+ $X2=3.685 $Y2=2
r107 25 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.085 $X2=3.6
+ $Y2=2
r108 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.6 $Y=2.085
+ $X2=3.6 $Y2=2.3
r109 23 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=2 $X2=3.6
+ $Y2=2
r110 23 24 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.515 $Y=2
+ $X2=2.695 $Y2=2
r111 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.61 $Y=2.085
+ $X2=2.695 $Y2=2
r112 19 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.61 $Y=2.085
+ $X2=2.61 $Y2=2.3
r113 6 52 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.485 $X2=8.02 $Y2=2.34
r114 6 47 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.485 $X2=8.02 $Y2=1.92
r115 5 44 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.935
+ $Y=1.485 $X2=7.08 $Y2=2.34
r116 4 42 600 $w=1.7e-07 $l=1.19134e-06 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=6.14 $Y2=2.34
r117 3 33 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=2.3
r118 2 27 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.485 $X2=3.6 $Y2=2.3
r119 1 21 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%VGND 1 2 3 4 5 16 18 20 22 27 32 37 47 48
+ 55 62 69 76
r113 76 79 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=7.525 $Y=0
+ $X2=7.525 $Y2=0.38
r114 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r115 69 72 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.055 $Y=0
+ $X2=3.055 $Y2=0.38
r116 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r117 62 65 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=2.115 $Y2=0.38
r118 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r119 55 58 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.175 $Y=0
+ $X2=1.175 $Y2=0.38
r120 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r121 48 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=7.59
+ $Y2=0
r122 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r123 45 76 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.715 $Y=0 $X2=7.525
+ $Y2=0
r124 45 47 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=8.05 $Y2=0
r125 44 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r126 43 44 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r127 41 44 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=7.13
+ $Y2=0
r128 41 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r129 40 43 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=7.13
+ $Y2=0
r130 40 41 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r131 38 69 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.055
+ $Y2=0
r132 38 40 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.245 $Y=0
+ $X2=3.45 $Y2=0
r133 37 76 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.525
+ $Y2=0
r134 37 43 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=7.13 $Y2=0
r135 36 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r136 36 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r137 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r138 33 62 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.115
+ $Y2=0
r139 33 35 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.53 $Y2=0
r140 32 69 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=3.055
+ $Y2=0
r141 32 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=2.53 $Y2=0
r142 31 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r143 31 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r144 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r145 28 55 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.175
+ $Y2=0
r146 28 30 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r147 27 62 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=2.115
+ $Y2=0
r148 27 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.925 $Y=0
+ $X2=1.61 $Y2=0
r149 26 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r150 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r151 23 51 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r152 23 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r153 22 55 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.175
+ $Y2=0
r154 22 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.69
+ $Y2=0
r155 20 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r156 20 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r157 16 51 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r158 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r159 5 79 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.235 $X2=7.55 $Y2=0.38
r160 4 72 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.38
r161 3 65 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r162 2 58 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.38
r163 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%A_485_47# 1 2 9 11 13
r25 11 13 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.695 $Y=0.74
+ $X2=4.07 $Y2=0.74
r26 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.61 $Y=0.655
+ $X2=2.695 $Y2=0.74
r27 7 9 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.61 $Y=0.655
+ $X2=2.61 $Y2=0.42
r28 2 13 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.74
r29 1 9 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%A_695_47# 1 2 3 16
r20 14 16 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.54 $Y=0.38
+ $X2=5.48 $Y2=0.38
r21 11 14 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.6 $Y=0.38 $X2=4.54
+ $Y2=0.38
r22 3 16 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.235 $X2=5.48 $Y2=0.38
r23 2 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.405
+ $Y=0.235 $X2=4.54 $Y2=0.38
r24 1 11 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.475
+ $Y=0.235 $X2=3.6 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_4%A_1194_47# 1 2 3 10 14 15 16 17 20
r33 18 20 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.02 $Y=0.645
+ $X2=8.02 $Y2=0.42
r34 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.935 $Y=0.73
+ $X2=8.02 $Y2=0.645
r35 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.935 $Y=0.73
+ $X2=7.165 $Y2=0.73
r36 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.08 $Y=0.645
+ $X2=7.165 $Y2=0.73
r37 14 23 3.40825 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.08 $Y=0.465
+ $X2=7.08 $Y2=0.36
r38 14 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.08 $Y=0.465
+ $X2=7.08 $Y2=0.645
r39 10 23 3.40825 $w=1.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=6.995 $Y=0.38
+ $X2=7.08 $Y2=0.36
r40 10 12 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=6.995 $Y=0.38
+ $X2=6.095 $Y2=0.38
r41 3 20 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=7.835
+ $Y=0.235 $X2=8.02 $Y2=0.42
r42 2 23 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.235 $X2=7.08 $Y2=0.42
r43 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.97
+ $Y=0.235 $X2=6.095 $Y2=0.38
.ends

