# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.075000 5.390000 1.275000 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA  0.617500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  1.825000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.576000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.635000 2.840000 0.905000 ;
        RECT 1.505000 1.445000 4.720000 1.665000 ;
        RECT 1.505000 1.665000 1.885000 2.465000 ;
        RECT 2.445000 1.665000 2.840000 2.465000 ;
        RECT 2.575000 0.905000 2.840000 1.445000 ;
        RECT 3.400000 1.665000 3.780000 2.465000 ;
        RECT 4.340000 1.665000 4.720000 2.465000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.715000 ;
      RECT 0.090000  0.715000 0.830000 0.905000 ;
      RECT 0.090000  1.445000 0.830000 1.665000 ;
      RECT 0.090000  1.665000 0.425000 2.465000 ;
      RECT 0.645000  0.085000 0.840000 0.545000 ;
      RECT 0.645000  1.835000 1.335000 2.635000 ;
      RECT 0.660000  0.905000 0.830000 1.075000 ;
      RECT 0.660000  1.075000 2.355000 1.275000 ;
      RECT 0.660000  1.275000 0.830000 1.445000 ;
      RECT 1.020000  1.445000 1.335000 1.835000 ;
      RECT 1.085000  0.255000 3.310000 0.465000 ;
      RECT 1.085000  0.465000 1.335000 0.905000 ;
      RECT 2.105000  1.835000 2.275000 2.635000 ;
      RECT 3.060000  0.465000 3.310000 0.715000 ;
      RECT 3.060000  0.715000 5.300000 0.905000 ;
      RECT 3.060000  1.835000 3.230000 2.635000 ;
      RECT 3.530000  0.085000 3.700000 0.545000 ;
      RECT 3.870000  0.255000 4.250000 0.715000 ;
      RECT 4.000000  1.835000 4.170000 2.635000 ;
      RECT 4.470000  0.085000 4.710000 0.545000 ;
      RECT 4.970000  0.255000 5.300000 0.715000 ;
      RECT 4.970000  1.495000 5.300000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2b_4
END LIBRARY
