* File: sky130_fd_sc_hdll__dlygate4sd2_1.pxi.spice
* Created: Wed Sep  2 08:30:22 2020
* 
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%A N_A_M1007_g N_A_M1005_g A A N_A_c_67_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%A
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%A_27_47# N_A_27_47#_M1005_s
+ N_A_27_47#_M1007_s N_A_27_47#_M1000_g N_A_27_47#_M1004_g N_A_27_47#_c_105_n
+ N_A_27_47#_c_99_n N_A_27_47#_c_100_n N_A_27_47#_c_101_n N_A_27_47#_c_106_n
+ N_A_27_47#_c_107_n N_A_27_47#_c_102_n N_A_27_47#_c_109_n N_A_27_47#_c_103_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%A_213_47# N_A_213_47#_M1000_d
+ N_A_213_47#_M1004_d N_A_213_47#_c_170_n N_A_213_47#_M1006_g
+ N_A_213_47#_c_177_n N_A_213_47#_M1002_g N_A_213_47#_c_171_n
+ N_A_213_47#_c_172_n N_A_213_47#_c_173_n N_A_213_47#_c_174_n
+ N_A_213_47#_c_175_n N_A_213_47#_c_180_n N_A_213_47#_c_176_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%A_213_47#
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%A_319_93# N_A_319_93#_M1006_s
+ N_A_319_93#_M1002_s N_A_319_93#_M1003_g N_A_319_93#_c_234_n
+ N_A_319_93#_M1001_g N_A_319_93#_c_247_n N_A_319_93#_c_235_n
+ N_A_319_93#_c_240_n N_A_319_93#_c_241_n N_A_319_93#_c_236_n
+ N_A_319_93#_c_243_n N_A_319_93#_c_237_n N_A_319_93#_c_238_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%A_319_93#
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%VPWR N_VPWR_M1007_d N_VPWR_M1002_d
+ N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_304_n VPWR
+ N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_300_n N_VPWR_c_308_n VPWR
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%VPWR
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%X N_X_M1001_d N_X_M1003_d X X X X X X
+ N_X_c_343_n X X PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%X
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%VGND N_VGND_M1005_d N_VGND_M1006_d
+ N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n VGND
+ N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n N_VGND_c_372_n VGND
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD2_1%VGND
cc_1 VNB N_A_M1005_g 0.0356862f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A 0.0125899f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_3 VNB N_A_c_67_n 0.0340348f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_27_47#_M1000_g 0.0341113f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_5 VNB N_A_27_47#_c_99_n 0.0186036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_100_n 0.00873805f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.53
cc_7 VNB N_A_27_47#_c_101_n 0.00988907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_102_n 0.00477608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_103_n 0.0242552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_213_47#_c_170_n 0.0415875f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_11 VNB N_A_213_47#_c_171_n 0.0097609f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_213_47#_c_172_n 4.49131e-19 $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_13 VNB N_A_213_47#_c_173_n 0.00459684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_213_47#_c_174_n 0.0453397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_213_47#_c_175_n 0.00575742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_213_47#_c_176_n 0.00131467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_319_93#_c_234_n 0.0216281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_319_93#_c_235_n 0.00521148f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_19 VNB N_A_319_93#_c_236_n 0.00651269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_319_93#_c_237_n 0.00154131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_319_93#_c_238_n 0.0330023f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_300_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB X 0.00638732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_343_n 0.0159232f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.53
cc_25 VNB X 0.0230432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_365_n 0.00493236f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_27 VNB N_VGND_c_366_n 0.00609109f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_28 VNB N_VGND_c_367_n 0.0351647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_368_n 0.00785847f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.16
cc_30 VNB N_VGND_c_369_n 0.0176957f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.16
cc_31 VNB N_VGND_c_370_n 0.0198931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_371_n 0.194223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_372_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_A_M1007_g 0.0644496f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=2.275
cc_35 VPB A 0.0179822f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_36 VPB N_A_c_67_n 0.00852761f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_37 VPB N_A_27_47#_M1004_g 0.0564089f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_38 VPB N_A_27_47#_c_105_n 0.0188411f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.16
cc_39 VPB N_A_27_47#_c_106_n 0.00971013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_107_n 0.012476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_102_n 6.81118e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_109_n 0.00337745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_103_n 0.00631651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_213_47#_c_177_n 0.0701267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_213_47#_c_172_n 0.0183355f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_46 VPB N_A_213_47#_c_174_n 0.0171648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_213_47#_c_180_n 0.00597064f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_319_93#_M1003_g 0.026562f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_49 VPB N_A_319_93#_c_240_n 0.0013599f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.16
cc_50 VPB N_A_319_93#_c_241_n 0.00317192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_319_93#_c_236_n 2.35122e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_319_93#_c_243_n 0.00283065f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.53
cc_53 VPB N_A_319_93#_c_238_n 0.0081194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_301_n 0.00493236f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_55 VPB N_VPWR_c_302_n 0.00586751f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_56 VPB N_VPWR_c_303_n 0.0365727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_304_n 0.00709097f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.16
cc_58 VPB N_VPWR_c_305_n 0.0176016f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.16
cc_59 VPB N_VPWR_c_306_n 0.0213696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_300_n 0.060682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_308_n 0.00406576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB X 0.0308524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB X 0.00895973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB X 0.00629578f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 N_A_M1005_g N_A_27_47#_M1000_g 0.0237725f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_66 N_A_M1007_g N_A_27_47#_M1004_g 0.0409596f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_67 A N_A_27_47#_M1004_g 8.58794e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_M1007_g N_A_27_47#_c_105_n 0.0037728f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_69 N_A_M1005_g N_A_27_47#_c_99_n 0.00709694f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_M1005_g N_A_27_47#_c_100_n 0.0137054f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_71 A N_A_27_47#_c_100_n 0.017067f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_72 N_A_c_67_n N_A_27_47#_c_100_n 0.00168708f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_73 A N_A_27_47#_c_101_n 0.0252593f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_c_67_n N_A_27_47#_c_101_n 0.00511105f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_M1007_g N_A_27_47#_c_106_n 0.0178074f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_76 A N_A_27_47#_c_106_n 0.017423f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_77 A N_A_27_47#_c_107_n 0.0271506f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A_c_67_n N_A_27_47#_c_107_n 8.59854e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_M1005_g N_A_27_47#_c_102_n 0.00363534f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_80 A N_A_27_47#_c_102_n 0.0232483f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A_c_67_n N_A_27_47#_c_102_n 8.544e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_M1007_g N_A_27_47#_c_109_n 0.00439862f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_83 A N_A_27_47#_c_109_n 0.0238071f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_84 A N_A_27_47#_c_103_n 8.94748e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_85 N_A_c_67_n N_A_27_47#_c_103_n 0.0213608f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_M1007_g N_VPWR_c_301_n 0.00304969f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_87 N_A_M1007_g N_VPWR_c_305_n 0.00523784f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_88 N_A_M1007_g N_VPWR_c_300_n 0.0077765f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_89 N_A_M1005_g N_VGND_c_365_n 0.00303707f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_90 N_A_M1005_g N_VGND_c_369_n 0.00436487f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_M1005_g N_VGND_c_371_n 0.00690659f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_27_47#_M1000_g N_A_213_47#_c_171_n 0.0111711f $X=0.975 $Y=0.445 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_c_102_n N_A_213_47#_c_171_n 0.0198042f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_c_103_n N_A_213_47#_c_171_n 5.89871e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_M1004_g N_A_213_47#_c_172_n 0.0195497f $X=0.975 $Y=2.275 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_c_106_n N_A_213_47#_c_172_n 0.0113209f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_c_102_n N_A_213_47#_c_172_n 0.00371586f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_c_109_n N_A_213_47#_c_172_n 0.0212546f $X=0.86 $Y=1.785 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_103_n N_A_213_47#_c_172_n 3.67773e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_102_n N_A_213_47#_c_174_n 2.17863e-19 $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_103_n N_A_213_47#_c_174_n 0.0110765f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_M1000_g N_A_213_47#_c_175_n 0.00679988f $X=0.975 $Y=0.445
+ $X2=0 $Y2=0
cc_103 N_A_27_47#_c_102_n N_A_213_47#_c_175_n 0.00294768f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_103_n N_A_213_47#_c_175_n 7.21452e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_M1004_g N_A_213_47#_c_180_n 0.00862725f $X=0.975 $Y=2.275
+ $X2=0 $Y2=0
cc_106 N_A_27_47#_c_102_n N_A_213_47#_c_176_n 0.0168575f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_103_n N_A_213_47#_c_176_n 0.0016685f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_M1004_g N_VPWR_c_301_n 0.00389952f $X=0.975 $Y=2.275 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_c_106_n N_VPWR_c_301_n 0.0151692f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_M1004_g N_VPWR_c_303_n 0.0052151f $X=0.975 $Y=2.275 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_c_106_n N_VPWR_c_303_n 0.0021103f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_c_105_n N_VPWR_c_305_n 0.0199397f $X=0.26 $Y=2.21 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_106_n N_VPWR_c_305_n 0.0031219f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_M1007_s N_VPWR_c_300_n 0.00242594f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_M1004_g N_VPWR_c_300_n 0.00905583f $X=0.975 $Y=2.275 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_105_n N_VPWR_c_300_n 0.0112839f $X=0.26 $Y=2.21 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_106_n N_VPWR_c_300_n 0.00921336f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_M1000_g N_VGND_c_365_n 0.00389952f $X=0.975 $Y=0.445 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_c_100_n N_VGND_c_365_n 0.0115001f $X=0.775 $Y=0.8 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_102_n N_VGND_c_365_n 0.00342769f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_M1000_g N_VGND_c_367_n 0.0052151f $X=0.975 $Y=0.445 $X2=0
+ $Y2=0
cc_122 N_A_27_47#_c_102_n N_VGND_c_367_n 0.0021103f $X=0.86 $Y=1.325 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_99_n N_VGND_c_369_n 0.0198425f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_100_n N_VGND_c_369_n 0.00312415f $X=0.775 $Y=0.8 $X2=0 $Y2=0
cc_125 N_A_27_47#_M1005_s N_VGND_c_371_n 0.00281655f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_M1000_g N_VGND_c_371_n 0.00905583f $X=0.975 $Y=0.445 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_c_99_n N_VGND_c_371_n 0.010877f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_100_n N_VGND_c_371_n 0.00573429f $X=0.775 $Y=0.8 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_102_n N_VGND_c_371_n 0.00355539f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_130 N_A_213_47#_c_177_n N_A_319_93#_M1003_g 0.0213988f $X=1.975 $Y=1.325
+ $X2=0 $Y2=0
cc_131 N_A_213_47#_c_170_n N_A_319_93#_c_234_n 0.0137479f $X=1.975 $Y=0.995
+ $X2=0 $Y2=0
cc_132 N_A_213_47#_c_172_n N_A_319_93#_c_247_n 0.0228797f $X=1.335 $Y=2.175
+ $X2=0 $Y2=0
cc_133 N_A_213_47#_c_170_n N_A_319_93#_c_235_n 0.013511f $X=1.975 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_A_213_47#_c_173_n N_A_319_93#_c_235_n 0.0178643f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_213_47#_c_174_n N_A_319_93#_c_235_n 0.00108706f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_213_47#_c_177_n N_A_319_93#_c_240_n 0.0200447f $X=1.975 $Y=1.325
+ $X2=0 $Y2=0
cc_137 N_A_213_47#_c_173_n N_A_319_93#_c_240_n 0.0114744f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_213_47#_c_174_n N_A_319_93#_c_240_n 9.55192e-19 $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_213_47#_c_172_n N_A_319_93#_c_241_n 0.012958f $X=1.335 $Y=2.175 $X2=0
+ $Y2=0
cc_140 N_A_213_47#_c_173_n N_A_319_93#_c_241_n 0.0117302f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A_213_47#_c_174_n N_A_319_93#_c_241_n 0.00509069f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_142 N_A_213_47#_c_170_n N_A_319_93#_c_236_n 0.0018158f $X=1.975 $Y=0.995
+ $X2=0 $Y2=0
cc_143 N_A_213_47#_c_173_n N_A_319_93#_c_236_n 0.0107502f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_144 N_A_213_47#_c_174_n N_A_319_93#_c_236_n 0.00118125f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_213_47#_c_177_n N_A_319_93#_c_243_n 0.00492289f $X=1.975 $Y=1.325
+ $X2=0 $Y2=0
cc_146 N_A_213_47#_c_170_n N_A_319_93#_c_237_n 3.3286e-19 $X=1.975 $Y=0.995
+ $X2=0 $Y2=0
cc_147 N_A_213_47#_c_171_n N_A_319_93#_c_237_n 0.0246532f $X=1.335 $Y=1.075
+ $X2=0 $Y2=0
cc_148 N_A_213_47#_c_173_n N_A_319_93#_c_237_n 0.0173672f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_213_47#_c_174_n N_A_319_93#_c_237_n 0.00562337f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_150 N_A_213_47#_c_175_n N_A_319_93#_c_237_n 0.00251361f $X=1.335 $Y=0.4 $X2=0
+ $Y2=0
cc_151 N_A_213_47#_c_173_n N_A_319_93#_c_238_n 9.30121e-19 $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_213_47#_c_174_n N_A_319_93#_c_238_n 0.0120031f $X=1.93 $Y=1.16 $X2=0
+ $Y2=0
cc_153 N_A_213_47#_c_180_n N_VPWR_c_301_n 0.0222152f $X=1.335 $Y=2.32 $X2=0
+ $Y2=0
cc_154 N_A_213_47#_c_177_n N_VPWR_c_302_n 0.0173349f $X=1.975 $Y=1.325 $X2=0
+ $Y2=0
cc_155 N_A_213_47#_c_177_n N_VPWR_c_303_n 0.00702461f $X=1.975 $Y=1.325 $X2=0
+ $Y2=0
cc_156 N_A_213_47#_c_180_n N_VPWR_c_303_n 0.026749f $X=1.335 $Y=2.32 $X2=0 $Y2=0
cc_157 N_A_213_47#_M1004_d N_VPWR_c_300_n 0.00209344f $X=1.065 $Y=2.065 $X2=0
+ $Y2=0
cc_158 N_A_213_47#_c_177_n N_VPWR_c_300_n 0.0145798f $X=1.975 $Y=1.325 $X2=0
+ $Y2=0
cc_159 N_A_213_47#_c_180_n N_VPWR_c_300_n 0.0159536f $X=1.335 $Y=2.32 $X2=0
+ $Y2=0
cc_160 N_A_213_47#_c_175_n N_VGND_c_365_n 0.0222152f $X=1.335 $Y=0.4 $X2=0 $Y2=0
cc_161 N_A_213_47#_c_170_n N_VGND_c_366_n 0.0124367f $X=1.975 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A_213_47#_c_170_n N_VGND_c_367_n 0.00527047f $X=1.975 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_213_47#_c_175_n N_VGND_c_367_n 0.0267806f $X=1.335 $Y=0.4 $X2=0 $Y2=0
cc_164 N_A_213_47#_M1000_d N_VGND_c_371_n 0.00209344f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_165 N_A_213_47#_c_170_n N_VGND_c_371_n 0.00902847f $X=1.975 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_213_47#_c_175_n N_VGND_c_371_n 0.0159581f $X=1.335 $Y=0.4 $X2=0 $Y2=0
cc_167 N_A_319_93#_c_240_n N_VPWR_M1002_d 0.0146765f $X=2.4 $Y=1.66 $X2=0 $Y2=0
cc_168 N_A_319_93#_c_243_n N_VPWR_M1002_d 0.00179207f $X=2.505 $Y=1.575 $X2=0
+ $Y2=0
cc_169 N_A_319_93#_M1003_g N_VPWR_c_302_n 0.00994494f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_319_93#_c_240_n N_VPWR_c_302_n 0.030862f $X=2.4 $Y=1.66 $X2=0 $Y2=0
cc_171 N_A_319_93#_c_238_n N_VPWR_c_302_n 3.81644e-19 $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_172 N_A_319_93#_c_247_n N_VPWR_c_303_n 0.00407287f $X=1.73 $Y=1.915 $X2=0
+ $Y2=0
cc_173 N_A_319_93#_M1003_g N_VPWR_c_306_n 0.00688798f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_319_93#_M1003_g N_VPWR_c_300_n 0.0138459f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_319_93#_c_247_n N_VPWR_c_300_n 0.00659363f $X=1.73 $Y=1.915 $X2=0
+ $Y2=0
cc_176 N_A_319_93#_c_234_n X 0.00501504f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_319_93#_M1003_g X 0.0155768f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_319_93#_c_234_n N_X_c_343_n 0.00820457f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_319_93#_M1003_g X 0.00382735f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_319_93#_c_234_n X 0.0115734f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_319_93#_c_236_n X 0.0321163f $X=2.505 $Y=1.325 $X2=0 $Y2=0
cc_182 N_A_319_93#_c_243_n X 0.00982184f $X=2.505 $Y=1.575 $X2=0 $Y2=0
cc_183 N_A_319_93#_M1003_g X 0.00231137f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_319_93#_c_240_n X 0.0135325f $X=2.4 $Y=1.66 $X2=0 $Y2=0
cc_185 N_A_319_93#_c_235_n N_VGND_M1006_d 0.00374668f $X=2.4 $Y=0.82 $X2=0 $Y2=0
cc_186 N_A_319_93#_c_236_n N_VGND_M1006_d 0.00353182f $X=2.505 $Y=1.325 $X2=0
+ $Y2=0
cc_187 N_A_319_93#_c_234_n N_VGND_c_366_n 0.00699004f $X=2.735 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_319_93#_c_235_n N_VGND_c_366_n 0.0198976f $X=2.4 $Y=0.82 $X2=0 $Y2=0
cc_189 N_A_319_93#_c_236_n N_VGND_c_366_n 0.0133517f $X=2.505 $Y=1.325 $X2=0
+ $Y2=0
cc_190 N_A_319_93#_c_238_n N_VGND_c_366_n 6.79215e-19 $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_A_319_93#_c_235_n N_VGND_c_367_n 0.00344355f $X=2.4 $Y=0.82 $X2=0 $Y2=0
cc_192 N_A_319_93#_c_237_n N_VGND_c_367_n 0.00546027f $X=1.72 $Y=0.675 $X2=0
+ $Y2=0
cc_193 N_A_319_93#_c_234_n N_VGND_c_370_n 0.00541359f $X=2.735 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_319_93#_c_236_n N_VGND_c_370_n 8.01519e-19 $X=2.505 $Y=1.325 $X2=0
+ $Y2=0
cc_195 N_A_319_93#_c_234_n N_VGND_c_371_n 0.011327f $X=2.735 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_319_93#_c_235_n N_VGND_c_371_n 0.00807282f $X=2.4 $Y=0.82 $X2=0 $Y2=0
cc_197 N_A_319_93#_c_236_n N_VGND_c_371_n 0.0022347f $X=2.505 $Y=1.325 $X2=0
+ $Y2=0
cc_198 N_A_319_93#_c_237_n N_VGND_c_371_n 0.00718111f $X=1.72 $Y=0.675 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_300_n N_X_M1003_d 0.00238012f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_200 N_VPWR_c_302_n X 0.0306504f $X=2.33 $Y=2 $X2=0 $Y2=0
cc_201 N_VPWR_c_306_n X 0.0210604f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_202 N_VPWR_c_300_n X 0.0125182f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_203 N_X_c_343_n N_VGND_c_366_n 0.0197349f $X=2.945 $Y=0.38 $X2=0 $Y2=0
cc_204 N_X_c_343_n N_VGND_c_370_n 0.0210139f $X=2.945 $Y=0.38 $X2=0 $Y2=0
cc_205 N_X_M1001_d N_VGND_c_371_n 0.00209319f $X=2.81 $Y=0.235 $X2=0 $Y2=0
cc_206 N_X_c_343_n N_VGND_c_371_n 0.0124133f $X=2.945 $Y=0.38 $X2=0 $Y2=0
