* File: sky130_fd_sc_hdll__o211ai_4.spice
* Created: Thu Aug 27 19:18:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o211ai_4.pex.spice"
.subckt sky130_fd_sc_hdll__o211ai_4  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM0_noxref N_VGND_M0_noxref_d N_A1_M0_noxref_g N_noxref_10_M0_noxref_s VNB
+ NSHORT L=0.15 W=0.65 AD=0.10725 AS=0.17225 PD=0.98 PS=1.83 NRD=9.228 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75007.6 A=0.0975 P=1.6 MULT=1
MM1_noxref N_noxref_10_M1_noxref_d N_A1_M1_noxref_g N_VGND_M0_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.1235 AS=0.10725 PD=1.03 PS=0.98 NRD=9.228 NRS=0 M=1
+ R=4.33333 SA=75000.7 SB=75007.1 A=0.0975 P=1.6 MULT=1
MM2_noxref N_VGND_M2_noxref_d N_A1_M2_noxref_g N_noxref_10_M1_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.1235 PD=0.93 PS=1.03 NRD=0 NRS=9.228 M=1
+ R=4.33333 SA=75001.2 SB=75006.6 A=0.0975 P=1.6 MULT=1
MM3_noxref N_noxref_10_M3_noxref_d N_A2_M3_noxref_g N_VGND_M2_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.10725 AS=0.091 PD=0.98 PS=0.93 NRD=9.228 NRS=0 M=1
+ R=4.33333 SA=75001.6 SB=75006.2 A=0.0975 P=1.6 MULT=1
MM4_noxref N_VGND_M4_noxref_d N_A2_M4_noxref_g N_noxref_10_M3_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=9.228 NRS=0 M=1
+ R=4.33333 SA=75002.1 SB=75005.7 A=0.0975 P=1.6 MULT=1
MM5_noxref N_noxref_10_M5_noxref_d N_A2_M5_noxref_g N_VGND_M4_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.1235 AS=0.10725 PD=1.03 PS=0.98 NRD=9.228 NRS=0 M=1
+ R=4.33333 SA=75002.6 SB=75005.2 A=0.0975 P=1.6 MULT=1
MM6_noxref N_VGND_M6_noxref_d N_A2_M6_noxref_g N_noxref_10_M5_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.1105 AS=0.1235 PD=0.99 PS=1.03 NRD=0 NRS=9.228 M=1
+ R=4.33333 SA=75003.1 SB=75004.7 A=0.0975 P=1.6 MULT=1
MM7_noxref N_noxref_10_M7_noxref_d N_A1_M7_noxref_g N_VGND_M6_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.10075 AS=0.1105 PD=0.96 PS=0.99 NRD=1.836 NRS=11.076
+ M=1 R=4.33333 SA=75003.6 SB=75004.2 A=0.0975 P=1.6 MULT=1
MM8_noxref N_noxref_12_M8_noxref_d N_B1_M8_noxref_g N_noxref_10_M7_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.10725 AS=0.10075 PD=0.98 PS=0.96 NRD=9.228 NRS=3.684
+ M=1 R=4.33333 SA=75004.1 SB=75003.7 A=0.0975 P=1.6 MULT=1
MM9_noxref N_noxref_10_M9_noxref_d N_B1_M9_noxref_g N_noxref_12_M8_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.1235 AS=0.10725 PD=1.03 PS=0.98 NRD=9.228 NRS=0 M=1
+ R=4.33333 SA=75004.5 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM10_noxref noxref_13 N_B1_M10_noxref_g N_noxref_10_M9_noxref_d VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.1235 PD=0.92 PS=1.03 NRD=14.76 NRS=9.228 M=1
+ R=4.33333 SA=75005.1 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM11_noxref N_Y_M11_noxref_d N_C1_M11_noxref_g noxref_13 VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=14.76 M=1 R=4.33333
+ SA=75005.5 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM12_noxref N_noxref_12_M12_noxref_d N_C1_M12_noxref_g N_Y_M11_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1
+ R=4.33333 SA=75006 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM13_noxref N_Y_M13_noxref_d N_C1_M13_noxref_g N_noxref_12_M12_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1
+ R=4.33333 SA=75006.4 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM14_noxref noxref_14 N_C1_M14_noxref_g N_Y_M13_noxref_d VNB NSHORT L=0.15
+ W=0.65 AD=0.1235 AS=0.12025 PD=1.03 PS=1.02 NRD=24.912 NRS=8.304 M=1 R=4.33333
+ SA=75007 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM15_noxref N_noxref_10_M15_noxref_d N_B1_M15_noxref_g noxref_14 VNB NSHORT
+ L=0.15 W=0.65 AD=0.25675 AS=0.1235 PD=2.09 PS=1.03 NRD=0 NRS=24.912 M=1
+ R=4.33333 SA=75007.5 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1011 N_A_118_297#_M1011_d N_A1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90007.8 A=0.18 P=2.36 MULT=1
MM1014 N_A_118_297#_M1011_d N_A1_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90007.3 A=0.18 P=2.36 MULT=1
MM1017 N_A_118_297#_M1017_d N_A1_M1017_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90006.8 A=0.18 P=2.36 MULT=1
MM1002 N_Y_M1002_d N_A2_M1002_g N_A_118_297#_M1017_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.6
+ SB=90006.3 A=0.18 P=2.36 MULT=1
MM1021 N_Y_M1002_d N_A2_M1021_g N_A_118_297#_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.1
+ SB=90005.9 A=0.18 P=2.36 MULT=1
MM1027 N_Y_M1027_d N_A2_M1027_g N_A_118_297#_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.6
+ SB=90005.4 A=0.18 P=2.36 MULT=1
MM1029 N_Y_M1027_d N_A2_M1029_g N_A_118_297#_M1029_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.1
+ SB=90004.9 A=0.18 P=2.36 MULT=1
MM1024 N_A_118_297#_M1029_s N_A1_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.17 PD=1.3 PS=1.34 NRD=1.9503 NRS=5.8903 M=1 R=5.55556 SA=90003.5
+ SB=90004.4 A=0.18 P=2.36 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_VPWR_M1024_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.17 PD=1.3 PS=1.34 NRD=1.9503 NRS=5.8903 M=1 R=5.55556 SA=90004.1
+ SB=90003.9 A=0.18 P=2.36 MULT=1
MM1009 N_Y_M1006_d N_B1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90004.5
+ SB=90003.4 A=0.18 P=2.36 MULT=1
MM1012 N_Y_M1012_d N_B1_M1012_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.15 PD=1.29 PS=1.3 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90005 SB=90002.9
+ A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_C1_M1001_g N_Y_M1012_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.5
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1001_d N_C1_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006 SB=90002
+ A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1023_d N_C1_M1023_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006.4
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1031 N_VPWR_M1023_d N_C1_M1031_g N_Y_M1031_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006.9
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1025 N_Y_M1031_s N_B1_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.685 PD=1.29 PS=3.37 NRD=0.9653 NRS=78.7803 M=1 R=5.55556 SA=90007.4
+ SB=90000.6 A=0.18 P=2.36 MULT=1
DX32_noxref VNB VPB NWDIODE A=14.6376 P=21.45
pX33_noxref noxref_15 A2 A2 PROBETYPE=1
pX34_noxref noxref_16 B1 B1 PROBETYPE=1
pX35_noxref noxref_17 C1 C1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o211ai_4.pxi.spice"
*
.ends
*
*
