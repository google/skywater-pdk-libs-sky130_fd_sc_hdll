* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
X0 VPWR A a_1187_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_797_297# a_27_297# a_331_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_797_297# B a_1187_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 Y a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_331_297# a_27_297# a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_27_297# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND a_27_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y a_207_47# a_331_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR A a_1187_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 Y a_207_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND a_27_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_1187_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VGND D_N a_207_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 Y a_207_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_27_297# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_331_297# a_27_297# a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 a_1187_297# B a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_331_297# a_207_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 Y a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Y a_207_47# a_331_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 a_797_297# B a_1187_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 VGND a_207_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_1187_297# B a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_797_297# a_27_297# a_331_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 VGND a_207_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_1187_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 VPWR D_N a_207_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 a_331_297# a_207_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
