* File: sky130_fd_sc_hdll__or2b_4.pxi.spice
* Created: Thu Aug 27 19:23:58 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR2B_4%B_N N_B_N_c_79_n N_B_N_c_80_n N_B_N_M1001_g
+ N_B_N_M1000_g B_N B_N B_N N_B_N_c_78_n PM_SKY130_FD_SC_HDLL__OR2B_4%B_N
x_PM_SKY130_FD_SC_HDLL__OR2B_4%A_27_53# N_A_27_53#_M1000_s N_A_27_53#_M1001_d
+ N_A_27_53#_c_102_n N_A_27_53#_M1004_g N_A_27_53#_c_109_n N_A_27_53#_M1005_g
+ N_A_27_53#_c_103_n N_A_27_53#_c_104_n N_A_27_53#_c_105_n N_A_27_53#_c_106_n
+ N_A_27_53#_c_107_n N_A_27_53#_c_108_n N_A_27_53#_c_113_n
+ PM_SKY130_FD_SC_HDLL__OR2B_4%A_27_53#
x_PM_SKY130_FD_SC_HDLL__OR2B_4%A N_A_c_163_n N_A_M1003_g N_A_c_164_n N_A_M1007_g
+ A A PM_SKY130_FD_SC_HDLL__OR2B_4%A
x_PM_SKY130_FD_SC_HDLL__OR2B_4%A_229_297# N_A_229_297#_M1004_d
+ N_A_229_297#_M1005_s N_A_229_297#_c_194_n N_A_229_297#_M1008_g
+ N_A_229_297#_c_201_n N_A_229_297#_M1002_g N_A_229_297#_c_195_n
+ N_A_229_297#_M1009_g N_A_229_297#_c_202_n N_A_229_297#_M1006_g
+ N_A_229_297#_c_196_n N_A_229_297#_M1010_g N_A_229_297#_c_203_n
+ N_A_229_297#_M1011_g N_A_229_297#_c_204_n N_A_229_297#_M1012_g
+ N_A_229_297#_c_197_n N_A_229_297#_M1013_g N_A_229_297#_c_205_n
+ N_A_229_297#_c_198_n N_A_229_297#_c_219_n N_A_229_297#_c_207_n
+ N_A_229_297#_c_238_n N_A_229_297#_c_208_n N_A_229_297#_c_273_p
+ N_A_229_297#_c_209_n N_A_229_297#_c_199_n N_A_229_297#_c_200_n
+ PM_SKY130_FD_SC_HDLL__OR2B_4%A_229_297#
x_PM_SKY130_FD_SC_HDLL__OR2B_4%VPWR N_VPWR_M1001_s N_VPWR_M1007_d N_VPWR_M1006_d
+ N_VPWR_M1012_d N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n
+ N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n
+ VPWR N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_320_n N_VPWR_c_333_n
+ PM_SKY130_FD_SC_HDLL__OR2B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__OR2B_4%X N_X_M1008_d N_X_M1010_d N_X_M1002_s N_X_M1011_s
+ N_X_c_390_n N_X_c_428_n N_X_c_393_n N_X_c_381_n N_X_c_382_n N_X_c_405_n
+ N_X_c_430_n N_X_c_386_n N_X_c_383_n N_X_c_411_n N_X_c_387_n N_X_c_384_n X X
+ PM_SKY130_FD_SC_HDLL__OR2B_4%X
x_PM_SKY130_FD_SC_HDLL__OR2B_4%VGND N_VGND_M1000_d N_VGND_M1003_d N_VGND_M1009_s
+ N_VGND_M1013_s N_VGND_c_456_n N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n
+ N_VGND_c_460_n N_VGND_c_461_n N_VGND_c_462_n N_VGND_c_463_n N_VGND_c_464_n
+ VGND N_VGND_c_465_n N_VGND_c_466_n N_VGND_c_467_n N_VGND_c_468_n
+ PM_SKY130_FD_SC_HDLL__OR2B_4%VGND
cc_1 VNB N_B_N_M1000_g 0.0401066f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_2 VNB B_N 0.00936139f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_B_N_c_78_n 0.0412036f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_27_53#_c_102_n 0.019479f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_5 VNB N_A_27_53#_c_103_n 0.034905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_53#_c_104_n 0.0136875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_53#_c_105_n 0.0205152f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_8 VNB N_A_27_53#_c_106_n 0.00290113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_53#_c_107_n 0.00967243f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_10 VNB N_A_27_53#_c_108_n 0.0129276f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_11 VNB N_A_c_163_n 0.0173697f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_12 VNB N_A_c_164_n 0.0272921f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_13 VNB A 0.00812636f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_14 VNB N_A_229_297#_c_194_n 0.0176527f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_15 VNB N_A_229_297#_c_195_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_229_297#_c_196_n 0.0172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_229_297#_c_197_n 0.02013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_229_297#_c_198_n 0.00216527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_229_297#_c_199_n 0.00306421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_229_297#_c_200_n 0.0759666f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_320_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_381_n 0.00247032f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.16
cc_23 VNB N_X_c_382_n 0.00336485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_383_n 0.013209f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_384_n 0.00262156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.0241415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_456_n 0.00666349f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_28 VNB N_VGND_c_457_n 0.00469169f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_29 VNB N_VGND_c_458_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_459_n 0.0228178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_460_n 0.00336608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_461_n 0.0203085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_462_n 0.00324283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_463_n 0.0196806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_464_n 0.00324283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_465_n 0.0142408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_466_n 0.244283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_467_n 0.018858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_468_n 0.0207275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VPB N_B_N_c_79_n 0.0403857f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_41 VPB N_B_N_c_80_n 0.0325653f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_42 VPB B_N 0.0295284f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_43 VPB N_B_N_c_78_n 0.0101702f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_44 VPB N_A_27_53#_c_109_n 0.0190122f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_45 VPB N_A_27_53#_c_103_n 0.0140754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_53#_c_104_n 0.0072327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_53#_c_108_n 0.0100117f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_48 VPB N_A_27_53#_c_113_n 0.0156704f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.16
cc_49 VPB N_A_c_164_n 0.0257831f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_50 VPB N_A_229_297#_c_201_n 0.0164974f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_51 VPB N_A_229_297#_c_202_n 0.0159111f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_52 VPB N_A_229_297#_c_203_n 0.0158526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_229_297#_c_204_n 0.019194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_229_297#_c_205_n 0.010652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_229_297#_c_198_n 0.00177712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_229_297#_c_207_n 0.00666923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_229_297#_c_208_n 0.00111937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_229_297#_c_209_n 0.00261924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_229_297#_c_200_n 0.0462269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_321_n 0.00995082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_322_n 0.0191035f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_323_n 0.00534879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_324_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.16
cc_64 VPB N_VPWR_c_325_n 0.00518f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.87
cc_65 VPB N_VPWR_c_326_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_327_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_328_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_329_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_330_n 0.0480363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_331_n 0.0140765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_320_n 0.0611893f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_333_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_X_c_386_n 0.0199149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_X_c_387_n 0.0034365f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB X 0.00854832f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 N_B_N_c_78_n N_A_27_53#_c_103_n 0.0117538f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B_N_M1000_g N_A_27_53#_c_105_n 0.00300084f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_78 N_B_N_M1000_g N_A_27_53#_c_106_n 0.0196695f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_79 N_B_N_c_78_n N_A_27_53#_c_106_n 0.00111307f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_80 B_N N_A_27_53#_c_107_n 0.0275042f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_81 N_B_N_c_78_n N_A_27_53#_c_107_n 0.00803194f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B_N_M1000_g N_A_27_53#_c_108_n 0.00895928f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_83 B_N N_A_27_53#_c_108_n 0.0170242f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_84 N_B_N_c_79_n N_A_27_53#_c_113_n 0.0165589f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_85 N_B_N_c_80_n N_A_27_53#_c_113_n 0.00705181f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_86 B_N N_A_27_53#_c_113_n 0.0389673f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_87 N_B_N_c_80_n N_VPWR_c_322_n 0.00654989f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_88 B_N N_VPWR_c_322_n 0.0225917f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_89 N_B_N_c_80_n N_VPWR_c_330_n 0.00743866f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_90 N_B_N_c_80_n N_VPWR_c_320_n 0.0148061f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_91 B_N N_VPWR_c_320_n 0.0041505f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_92 N_B_N_M1000_g N_VGND_c_466_n 0.00754515f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_93 N_B_N_M1000_g N_VGND_c_467_n 0.00413798f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_94 N_B_N_M1000_g N_VGND_c_468_n 0.00501457f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_95 N_A_27_53#_c_102_n N_A_c_163_n 0.011608f $X=1.47 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_96 N_A_27_53#_c_109_n N_A_c_164_n 0.0666158f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_27_53#_c_104_n N_A_c_164_n 0.0278976f $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A_27_53#_c_104_n A 0.00145041f $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_27_53#_c_109_n N_A_229_297#_c_205_n 0.0234665f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_100 N_A_27_53#_c_113_n N_A_229_297#_c_205_n 0.0568606f $X=0.73 $Y=2.2 $X2=0
+ $Y2=0
cc_101 N_A_27_53#_c_102_n N_A_229_297#_c_198_n 0.00284611f $X=1.47 $Y=0.995
+ $X2=0 $Y2=0
cc_102 N_A_27_53#_c_109_n N_A_229_297#_c_198_n 0.00139725f $X=1.505 $Y=1.41
+ $X2=0 $Y2=0
cc_103 N_A_27_53#_c_103_n N_A_229_297#_c_198_n 0.00853799f $X=1.395 $Y=1.16
+ $X2=0 $Y2=0
cc_104 N_A_27_53#_c_104_n N_A_229_297#_c_198_n 0.0124219f $X=1.395 $Y=0.995
+ $X2=0 $Y2=0
cc_105 N_A_27_53#_c_108_n N_A_229_297#_c_198_n 0.0250557f $X=0.73 $Y=1.325 $X2=0
+ $Y2=0
cc_106 N_A_27_53#_c_113_n N_A_229_297#_c_198_n 0.00418496f $X=0.73 $Y=2.2 $X2=0
+ $Y2=0
cc_107 N_A_27_53#_c_102_n N_A_229_297#_c_219_n 0.0127846f $X=1.47 $Y=0.995 $X2=0
+ $Y2=0
cc_108 N_A_27_53#_c_109_n N_A_229_297#_c_207_n 0.00446962f $X=1.505 $Y=1.41
+ $X2=0 $Y2=0
cc_109 N_A_27_53#_c_104_n N_A_229_297#_c_207_n 3.24848e-19 $X=1.395 $Y=0.995
+ $X2=0 $Y2=0
cc_110 N_A_27_53#_c_109_n N_A_229_297#_c_209_n 0.00291914f $X=1.505 $Y=1.41
+ $X2=0 $Y2=0
cc_111 N_A_27_53#_c_103_n N_A_229_297#_c_209_n 0.00858393f $X=1.395 $Y=1.16
+ $X2=0 $Y2=0
cc_112 N_A_27_53#_c_108_n N_A_229_297#_c_209_n 0.0109731f $X=0.73 $Y=1.325 $X2=0
+ $Y2=0
cc_113 N_A_27_53#_c_113_n N_A_229_297#_c_209_n 0.0102315f $X=0.73 $Y=2.2 $X2=0
+ $Y2=0
cc_114 N_A_27_53#_c_102_n N_A_229_297#_c_199_n 0.0069639f $X=1.47 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_A_27_53#_c_104_n N_A_229_297#_c_199_n 0.00157803f $X=1.395 $Y=0.995
+ $X2=0 $Y2=0
cc_116 N_A_27_53#_c_108_n N_A_229_297#_c_199_n 0.00814809f $X=0.73 $Y=1.325
+ $X2=0 $Y2=0
cc_117 N_A_27_53#_c_113_n N_VPWR_c_322_n 0.0167625f $X=0.73 $Y=2.2 $X2=0 $Y2=0
cc_118 N_A_27_53#_c_109_n N_VPWR_c_330_n 0.00483853f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_27_53#_c_113_n N_VPWR_c_330_n 0.0118139f $X=0.73 $Y=2.2 $X2=0 $Y2=0
cc_120 N_A_27_53#_M1001_d N_VPWR_c_320_n 0.00635031f $X=0.585 $Y=2.065 $X2=0
+ $Y2=0
cc_121 N_A_27_53#_c_109_n N_VPWR_c_320_n 0.00854743f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_122 N_A_27_53#_c_113_n N_VPWR_c_320_n 0.00646998f $X=0.73 $Y=2.2 $X2=0 $Y2=0
cc_123 N_A_27_53#_c_102_n N_VGND_c_459_n 0.00402575f $X=1.47 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_A_27_53#_c_102_n N_VGND_c_466_n 0.00693531f $X=1.47 $Y=0.995 $X2=0
+ $Y2=0
cc_125 N_A_27_53#_c_105_n N_VGND_c_466_n 0.0117861f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_27_53#_c_106_n N_VGND_c_466_n 0.00503364f $X=0.645 $Y=0.82 $X2=0
+ $Y2=0
cc_127 N_A_27_53#_c_108_n N_VGND_c_466_n 0.00106095f $X=0.73 $Y=1.325 $X2=0
+ $Y2=0
cc_128 N_A_27_53#_c_105_n N_VGND_c_467_n 0.0192939f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_129 N_A_27_53#_c_106_n N_VGND_c_467_n 0.00299761f $X=0.645 $Y=0.82 $X2=0
+ $Y2=0
cc_130 N_A_27_53#_c_102_n N_VGND_c_468_n 0.00700085f $X=1.47 $Y=0.995 $X2=0
+ $Y2=0
cc_131 N_A_27_53#_c_103_n N_VGND_c_468_n 0.0058713f $X=1.395 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_27_53#_c_108_n N_VGND_c_468_n 0.0327468f $X=0.73 $Y=1.325 $X2=0 $Y2=0
cc_133 N_A_c_163_n N_A_229_297#_c_194_n 0.0155072f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_164_n N_A_229_297#_c_201_n 0.0281441f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_164_n N_A_229_297#_c_205_n 0.00356582f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_c_163_n N_A_229_297#_c_198_n 0.00173941f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_164_n N_A_229_297#_c_198_n 0.00177124f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_138 A N_A_229_297#_c_198_n 0.016247f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_139 N_A_c_163_n N_A_229_297#_c_219_n 0.0060188f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_c_164_n N_A_229_297#_c_207_n 0.0207545f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_141 A N_A_229_297#_c_207_n 0.0536724f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_142 A N_A_229_297#_c_238_n 0.0116153f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A_c_164_n N_A_229_297#_c_208_n 2.0275e-19 $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_144 A N_A_229_297#_c_208_n 0.00176792f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A_c_163_n N_A_229_297#_c_199_n 0.00290011f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_146 A N_A_229_297#_c_199_n 0.00939662f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A_c_164_n N_A_229_297#_c_200_n 0.0254411f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_148 A N_A_229_297#_c_200_n 0.0140488f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A_c_164_n N_VPWR_c_323_n 0.0117805f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_164_n N_VPWR_c_330_n 0.00702461f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_164_n N_VPWR_c_320_n 0.0127233f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_163_n N_VGND_c_456_n 0.0086257f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_153 A N_VGND_c_456_n 0.0147599f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A_c_163_n N_VGND_c_459_n 0.00543342f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_163_n N_VGND_c_466_n 0.0100364f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_229_297#_c_207_n N_VPWR_M1007_d 0.00287935f $X=2.69 $Y=1.53 $X2=0
+ $Y2=0
cc_157 N_A_229_297#_c_201_n N_VPWR_c_323_n 0.00315364f $X=2.455 $Y=1.41 $X2=0
+ $Y2=0
cc_158 N_A_229_297#_c_205_n N_VPWR_c_323_n 0.0213641f $X=1.27 $Y=1.63 $X2=0
+ $Y2=0
cc_159 N_A_229_297#_c_207_n N_VPWR_c_323_n 0.0162556f $X=2.69 $Y=1.53 $X2=0
+ $Y2=0
cc_160 N_A_229_297#_c_202_n N_VPWR_c_324_n 0.00300743f $X=2.925 $Y=1.41 $X2=0
+ $Y2=0
cc_161 N_A_229_297#_c_203_n N_VPWR_c_324_n 0.00300743f $X=3.395 $Y=1.41 $X2=0
+ $Y2=0
cc_162 N_A_229_297#_c_204_n N_VPWR_c_325_n 0.00479105f $X=3.865 $Y=1.41 $X2=0
+ $Y2=0
cc_163 N_A_229_297#_c_201_n N_VPWR_c_326_n 0.00702461f $X=2.455 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_229_297#_c_202_n N_VPWR_c_326_n 0.00702461f $X=2.925 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_A_229_297#_c_203_n N_VPWR_c_328_n 0.00702461f $X=3.395 $Y=1.41 $X2=0
+ $Y2=0
cc_166 N_A_229_297#_c_204_n N_VPWR_c_328_n 0.00702461f $X=3.865 $Y=1.41 $X2=0
+ $Y2=0
cc_167 N_A_229_297#_c_205_n N_VPWR_c_330_n 0.0342422f $X=1.27 $Y=1.63 $X2=0
+ $Y2=0
cc_168 N_A_229_297#_M1005_s N_VPWR_c_320_n 0.00217517f $X=1.145 $Y=1.485 $X2=0
+ $Y2=0
cc_169 N_A_229_297#_c_201_n N_VPWR_c_320_n 0.0125915f $X=2.455 $Y=1.41 $X2=0
+ $Y2=0
cc_170 N_A_229_297#_c_202_n N_VPWR_c_320_n 0.00693457f $X=2.925 $Y=1.41 $X2=0
+ $Y2=0
cc_171 N_A_229_297#_c_203_n N_VPWR_c_320_n 0.00693457f $X=3.395 $Y=1.41 $X2=0
+ $Y2=0
cc_172 N_A_229_297#_c_204_n N_VPWR_c_320_n 0.0134797f $X=3.865 $Y=1.41 $X2=0
+ $Y2=0
cc_173 N_A_229_297#_c_205_n N_VPWR_c_320_n 0.0192181f $X=1.27 $Y=1.63 $X2=0
+ $Y2=0
cc_174 N_A_229_297#_c_207_n A_319_297# 0.00442604f $X=2.69 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A_229_297#_c_207_n N_X_M1002_s 0.00189183f $X=2.69 $Y=1.53 $X2=0 $Y2=0
cc_176 N_A_229_297#_c_194_n N_X_c_390_n 0.00499768f $X=2.43 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_229_297#_c_195_n N_X_c_390_n 0.00672047f $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_229_297#_c_196_n N_X_c_390_n 5.78063e-19 $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_229_297#_c_207_n N_X_c_393_n 0.014924f $X=2.69 $Y=1.53 $X2=0 $Y2=0
cc_180 N_A_229_297#_c_200_n N_X_c_393_n 6.22666e-19 $X=3.865 $Y=1.202 $X2=0
+ $Y2=0
cc_181 N_A_229_297#_c_195_n N_X_c_381_n 0.0087433f $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_229_297#_c_196_n N_X_c_381_n 0.00879805f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_229_297#_c_238_n N_X_c_381_n 3.39565e-19 $X=2.775 $Y=1.245 $X2=0
+ $Y2=0
cc_184 N_A_229_297#_c_273_p N_X_c_381_n 0.0387503f $X=3.635 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_229_297#_c_200_n N_X_c_381_n 0.00345061f $X=3.865 $Y=1.202 $X2=0
+ $Y2=0
cc_186 N_A_229_297#_c_194_n N_X_c_382_n 0.00286107f $X=2.43 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_229_297#_c_195_n N_X_c_382_n 0.00113678f $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_229_297#_c_207_n N_X_c_382_n 0.00759496f $X=2.69 $Y=1.53 $X2=0 $Y2=0
cc_189 N_A_229_297#_c_238_n N_X_c_382_n 0.0142226f $X=2.775 $Y=1.245 $X2=0 $Y2=0
cc_190 N_A_229_297#_c_200_n N_X_c_382_n 0.00414235f $X=3.865 $Y=1.202 $X2=0
+ $Y2=0
cc_191 N_A_229_297#_c_195_n N_X_c_405_n 5.59948e-19 $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_229_297#_c_196_n N_X_c_405_n 0.00641775f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_229_297#_c_204_n N_X_c_386_n 0.0193054f $X=3.865 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_229_297#_c_200_n N_X_c_386_n 6.71711e-19 $X=3.865 $Y=1.202 $X2=0
+ $Y2=0
cc_195 N_A_229_297#_c_197_n N_X_c_383_n 0.0140086f $X=3.89 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_229_297#_c_273_p N_X_c_383_n 3.20053e-19 $X=3.635 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_229_297#_c_202_n N_X_c_411_n 0.013137f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_229_297#_c_207_n N_X_c_411_n 0.00179336f $X=2.69 $Y=1.53 $X2=0 $Y2=0
cc_199 N_A_229_297#_c_273_p N_X_c_411_n 0.00502147f $X=3.635 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_229_297#_c_200_n N_X_c_411_n 9.61223e-19 $X=3.865 $Y=1.202 $X2=0
+ $Y2=0
cc_201 N_A_229_297#_c_202_n N_X_c_387_n 0.00685448f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_229_297#_c_203_n N_X_c_387_n 0.0215096f $X=3.395 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_229_297#_c_207_n N_X_c_387_n 0.0121608f $X=2.69 $Y=1.53 $X2=0 $Y2=0
cc_204 N_A_229_297#_c_273_p N_X_c_387_n 0.0487655f $X=3.635 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_229_297#_c_200_n N_X_c_387_n 0.0134576f $X=3.865 $Y=1.202 $X2=0 $Y2=0
cc_206 N_A_229_297#_c_196_n N_X_c_384_n 0.00116733f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_229_297#_c_273_p N_X_c_384_n 0.0302634f $X=3.635 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_229_297#_c_200_n N_X_c_384_n 0.00485436f $X=3.865 $Y=1.202 $X2=0
+ $Y2=0
cc_209 N_A_229_297#_c_204_n X 0.00133905f $X=3.865 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_229_297#_c_197_n X 0.019437f $X=3.89 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_229_297#_c_273_p X 0.00919972f $X=3.635 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_229_297#_c_194_n N_VGND_c_456_n 0.00303405f $X=2.43 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_229_297#_c_219_n N_VGND_c_456_n 0.0303769f $X=1.68 $Y=0.4 $X2=0 $Y2=0
cc_214 N_A_229_297#_c_195_n N_VGND_c_457_n 0.00431919f $X=2.9 $Y=0.995 $X2=0
+ $Y2=0
cc_215 N_A_229_297#_c_196_n N_VGND_c_457_n 0.00276126f $X=3.37 $Y=0.995 $X2=0
+ $Y2=0
cc_216 N_A_229_297#_c_197_n N_VGND_c_458_n 0.00438629f $X=3.89 $Y=0.995 $X2=0
+ $Y2=0
cc_217 N_A_229_297#_c_219_n N_VGND_c_459_n 0.0168234f $X=1.68 $Y=0.4 $X2=0 $Y2=0
cc_218 N_A_229_297#_c_199_n N_VGND_c_459_n 0.00142085f $X=1.592 $Y=0.905 $X2=0
+ $Y2=0
cc_219 N_A_229_297#_c_194_n N_VGND_c_461_n 0.00542757f $X=2.43 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_229_297#_c_195_n N_VGND_c_461_n 0.00425814f $X=2.9 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_229_297#_c_196_n N_VGND_c_463_n 0.00425814f $X=3.37 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_229_297#_c_197_n N_VGND_c_463_n 0.00439206f $X=3.89 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_229_297#_M1004_d N_VGND_c_466_n 0.00218509f $X=1.545 $Y=0.235 $X2=0
+ $Y2=0
cc_224 N_A_229_297#_c_194_n N_VGND_c_466_n 0.0099246f $X=2.43 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_229_297#_c_195_n N_VGND_c_466_n 0.00611499f $X=2.9 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_229_297#_c_196_n N_VGND_c_466_n 0.00610757f $X=3.37 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_229_297#_c_197_n N_VGND_c_466_n 0.00727186f $X=3.89 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_229_297#_c_219_n N_VGND_c_466_n 0.0135032f $X=1.68 $Y=0.4 $X2=0 $Y2=0
cc_229 N_A_229_297#_c_199_n N_VGND_c_466_n 0.00306781f $X=1.592 $Y=0.905 $X2=0
+ $Y2=0
cc_230 N_A_229_297#_c_219_n N_VGND_c_468_n 0.0215368f $X=1.68 $Y=0.4 $X2=0 $Y2=0
cc_231 N_VPWR_c_320_n A_319_297# 0.00983149f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_232 N_VPWR_c_320_n N_X_M1002_s 0.0031047f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_233 N_VPWR_c_320_n N_X_M1011_s 0.00307556f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_234 N_VPWR_c_326_n N_X_c_428_n 0.0149311f $X=3.035 $Y=2.72 $X2=0 $Y2=0
cc_235 N_VPWR_c_320_n N_X_c_428_n 0.00955092f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_236 N_VPWR_c_328_n N_X_c_430_n 0.014675f $X=3.975 $Y=2.72 $X2=0 $Y2=0
cc_237 N_VPWR_c_320_n N_X_c_430_n 0.00948039f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_238 N_VPWR_M1012_d N_X_c_386_n 0.00487431f $X=3.955 $Y=1.485 $X2=0 $Y2=0
cc_239 N_VPWR_c_325_n N_X_c_386_n 0.0174922f $X=4.1 $Y=1.96 $X2=0 $Y2=0
cc_240 N_VPWR_c_324_n N_X_c_411_n 0.014185f $X=3.16 $Y=2.3 $X2=0 $Y2=0
cc_241 N_VPWR_c_320_n N_X_c_411_n 0.00762318f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_242 N_VPWR_M1006_d N_X_c_387_n 0.00557493f $X=3.015 $Y=1.485 $X2=0 $Y2=0
cc_243 N_VPWR_c_320_n N_X_c_387_n 0.00753105f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_244 N_X_c_381_n N_VGND_M1009_s 0.0025752f $X=3.415 $Y=0.82 $X2=0 $Y2=0
cc_245 N_X_c_383_n N_VGND_M1013_s 0.00525022f $X=4.105 $Y=0.82 $X2=0 $Y2=0
cc_246 N_X_c_382_n N_VGND_c_456_n 0.00788213f $X=2.855 $Y=0.82 $X2=0 $Y2=0
cc_247 N_X_c_390_n N_VGND_c_457_n 0.0159144f $X=2.69 $Y=0.4 $X2=0 $Y2=0
cc_248 N_X_c_381_n N_VGND_c_457_n 0.0118167f $X=3.415 $Y=0.82 $X2=0 $Y2=0
cc_249 N_X_c_383_n N_VGND_c_458_n 0.0123826f $X=4.105 $Y=0.82 $X2=0 $Y2=0
cc_250 N_X_c_390_n N_VGND_c_461_n 0.0182313f $X=2.69 $Y=0.4 $X2=0 $Y2=0
cc_251 N_X_c_381_n N_VGND_c_461_n 0.00260082f $X=3.415 $Y=0.82 $X2=0 $Y2=0
cc_252 N_X_c_381_n N_VGND_c_463_n 0.00193763f $X=3.415 $Y=0.82 $X2=0 $Y2=0
cc_253 N_X_c_405_n N_VGND_c_463_n 0.0188919f $X=3.63 $Y=0.4 $X2=0 $Y2=0
cc_254 N_X_c_383_n N_VGND_c_463_n 0.00248202f $X=4.105 $Y=0.82 $X2=0 $Y2=0
cc_255 N_X_c_383_n N_VGND_c_465_n 0.0049839f $X=4.105 $Y=0.82 $X2=0 $Y2=0
cc_256 N_X_M1008_d N_VGND_c_466_n 0.00257593f $X=2.505 $Y=0.235 $X2=0 $Y2=0
cc_257 N_X_M1010_d N_VGND_c_466_n 0.0030688f $X=3.445 $Y=0.235 $X2=0 $Y2=0
cc_258 N_X_c_390_n N_VGND_c_466_n 0.0138527f $X=2.69 $Y=0.4 $X2=0 $Y2=0
cc_259 N_X_c_381_n N_VGND_c_466_n 0.00963305f $X=3.415 $Y=0.82 $X2=0 $Y2=0
cc_260 N_X_c_405_n N_VGND_c_466_n 0.014059f $X=3.63 $Y=0.4 $X2=0 $Y2=0
cc_261 N_X_c_383_n N_VGND_c_466_n 0.0141878f $X=4.105 $Y=0.82 $X2=0 $Y2=0
