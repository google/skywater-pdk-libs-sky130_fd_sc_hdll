# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nor4b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.340000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.075000 2.650000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.860000 1.075000 3.660000 1.285000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.205000 1.075000 5.885000 1.285000 ;
        RECT 5.615000 1.285000 5.885000 1.955000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.219500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.895000 0.725000 ;
        RECT 0.515000 0.725000 4.270000 0.905000 ;
        RECT 1.455000 0.255000 1.835000 0.725000 ;
        RECT 2.950000 0.255000 3.330000 0.725000 ;
        RECT 3.890000 0.255000 4.270000 0.725000 ;
        RECT 3.980000 1.455000 4.490000 1.625000 ;
        RECT 3.980000 1.625000 4.230000 2.125000 ;
        RECT 4.065000 0.905000 4.270000 1.075000 ;
        RECT 4.065000 1.075000 4.490000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  1.455000 2.305000 1.625000 ;
      RECT 0.085000  1.625000 0.425000 2.465000 ;
      RECT 0.645000  1.795000 0.855000 2.635000 ;
      RECT 1.075000  1.625000 1.325000 2.465000 ;
      RECT 1.115000  0.085000 1.285000 0.555000 ;
      RECT 1.545000  1.795000 1.755000 2.295000 ;
      RECT 1.545000  2.295000 3.290000 2.465000 ;
      RECT 1.925000  1.625000 2.305000 2.125000 ;
      RECT 2.055000  0.085000 2.780000 0.555000 ;
      RECT 2.475000  1.455000 3.760000 1.625000 ;
      RECT 2.475000  1.625000 2.860000 2.125000 ;
      RECT 3.080000  1.795000 3.290000 2.295000 ;
      RECT 3.510000  1.625000 3.760000 2.295000 ;
      RECT 3.510000  2.295000 4.695000 2.465000 ;
      RECT 3.550000  0.085000 3.720000 0.555000 ;
      RECT 4.450000  1.795000 4.695000 2.295000 ;
      RECT 4.490000  0.085000 4.695000 0.895000 ;
      RECT 4.720000  1.075000 5.035000 1.245000 ;
      RECT 4.865000  0.380000 5.220000 0.905000 ;
      RECT 4.865000  0.905000 5.035000 1.075000 ;
      RECT 4.865000  1.245000 5.035000 2.035000 ;
      RECT 4.865000  2.035000 5.220000 2.450000 ;
      RECT 5.440000  0.085000 5.690000 0.825000 ;
      RECT 5.440000  2.135000 5.690000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4b_2
END LIBRARY
