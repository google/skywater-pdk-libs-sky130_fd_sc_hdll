* File: sky130_fd_sc_hdll__inv_6.pxi.spice
* Created: Wed Sep  2 08:33:18 2020
* 
x_PM_SKY130_FD_SC_HDLL__INV_6%A N_A_c_60_n N_A_M1000_g N_A_c_52_n N_A_M1001_g
+ N_A_c_61_n N_A_M1002_g N_A_c_53_n N_A_M1005_g N_A_c_62_n N_A_M1003_g
+ N_A_c_54_n N_A_M1006_g N_A_c_63_n N_A_M1004_g N_A_c_55_n N_A_M1008_g
+ N_A_c_64_n N_A_M1007_g N_A_c_56_n N_A_M1009_g N_A_c_65_n N_A_M1010_g
+ N_A_c_57_n N_A_M1011_g A A A A N_A_c_59_n A A A A
+ PM_SKY130_FD_SC_HDLL__INV_6%A
x_PM_SKY130_FD_SC_HDLL__INV_6%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_M1004_d
+ N_VPWR_M1010_d N_VPWR_c_163_n N_VPWR_c_164_n N_VPWR_c_165_n N_VPWR_c_166_n
+ N_VPWR_c_167_n N_VPWR_c_168_n N_VPWR_c_169_n N_VPWR_c_170_n N_VPWR_c_171_n
+ VPWR N_VPWR_c_172_n N_VPWR_c_162_n N_VPWR_c_174_n N_VPWR_c_175_n
+ PM_SKY130_FD_SC_HDLL__INV_6%VPWR
x_PM_SKY130_FD_SC_HDLL__INV_6%Y N_Y_M1001_s N_Y_M1006_s N_Y_M1009_s N_Y_M1000_s
+ N_Y_M1003_s N_Y_M1007_s N_Y_c_227_n N_Y_c_231_n N_Y_c_234_n N_Y_c_219_n
+ N_Y_c_220_n N_Y_c_242_n N_Y_c_246_n N_Y_c_250_n N_Y_c_221_n N_Y_c_255_n
+ N_Y_c_258_n N_Y_c_259_n N_Y_c_222_n Y Y Y Y N_Y_c_273_n Y
+ PM_SKY130_FD_SC_HDLL__INV_6%Y
x_PM_SKY130_FD_SC_HDLL__INV_6%VGND N_VGND_M1001_d N_VGND_M1005_d N_VGND_M1008_d
+ N_VGND_M1011_d N_VGND_c_327_n N_VGND_c_328_n N_VGND_c_329_n N_VGND_c_330_n
+ N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n VGND N_VGND_c_334_n
+ N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n N_VGND_c_339_n
+ VGND PM_SKY130_FD_SC_HDLL__INV_6%VGND
cc_1 VNB N_A_c_52_n 0.0224567f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_A_c_53_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_A_c_54_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_4 VNB N_A_c_55_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_A_c_56_n 0.0167382f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.995
cc_6 VNB N_A_c_57_n 0.0191128f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.995
cc_7 VNB A 0.00932659f $X=-0.19 $Y=-0.24 $X2=2.395 $Y2=1.105
cc_8 VNB N_A_c_59_n 0.129622f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.202
cc_9 VNB N_VPWR_c_162_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_10 VNB N_Y_c_219_n 0.00380351f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.985
cc_11 VNB N_Y_c_220_n 0.00137522f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.995
cc_12 VNB N_Y_c_221_n 0.00380351f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.105
cc_13 VNB N_Y_c_222_n 0.00113459f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_14 VNB Y 0.0182299f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.202
cc_15 VNB Y 0.0117385f $X=-0.19 $Y=-0.24 $X2=2.01 $Y2=1.2
cc_16 VNB N_VGND_c_327_n 0.011417f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_17 VNB N_VGND_c_328_n 0.0191933f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_18 VNB N_VGND_c_329_n 0.0201447f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_19 VNB N_VGND_c_330_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_20 VNB N_VGND_c_331_n 0.0206128f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_21 VNB N_VGND_c_332_n 0.00417249f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.985
cc_22 VNB N_VGND_c_333_n 0.00230383f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.41
cc_23 VNB N_VGND_c_334_n 0.01593f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.56
cc_24 VNB N_VGND_c_335_n 0.018164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_336_n 0.214466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_337_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.16
cc_27 VNB N_VGND_c_338_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_28 VNB N_VGND_c_339_n 0.00420379f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_29 VPB N_A_c_60_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_30 VPB N_A_c_61_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_31 VPB N_A_c_62_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_32 VPB N_A_c_63_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_33 VPB N_A_c_64_n 0.0162574f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_34 VPB N_A_c_65_n 0.0196202f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_35 VPB A 7.73822e-19 $X=-0.19 $Y=1.305 $X2=2.395 $Y2=1.105
cc_36 VPB N_A_c_59_n 0.0799008f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.202
cc_37 VPB N_VPWR_c_163_n 0.0110239f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_38 VPB N_VPWR_c_164_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_39 VPB N_VPWR_c_165_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_40 VPB N_VPWR_c_166_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_41 VPB N_VPWR_c_167_n 0.0206409f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_42 VPB N_VPWR_c_168_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.4 $Y2=0.56
cc_43 VPB N_VPWR_c_169_n 0.00474148f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.985
cc_44 VPB N_VPWR_c_170_n 0.0206409f $X=-0.19 $Y=1.305 $X2=2.87 $Y2=0.56
cc_45 VPB N_VPWR_c_171_n 0.0032427f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.105
cc_46 VPB N_VPWR_c_172_n 0.0185316f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_47 VPB N_VPWR_c_162_n 0.0601043f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_48 VPB N_VPWR_c_174_n 0.00324069f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.202
cc_49 VPB N_VPWR_c_175_n 0.00324069f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.202
cc_50 VPB Y 0.00833318f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.202
cc_51 VPB Y 0.00985087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 N_A_c_60_n N_VPWR_c_164_n 0.00736507f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_53 A N_VPWR_c_164_n 0.00477961f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A_c_59_n N_VPWR_c_164_n 0.00137444f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_55 N_A_c_60_n N_VPWR_c_165_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_56 N_A_c_61_n N_VPWR_c_165_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_57 N_A_c_61_n N_VPWR_c_166_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_58 N_A_c_62_n N_VPWR_c_166_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A_c_62_n N_VPWR_c_167_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_c_63_n N_VPWR_c_167_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_c_63_n N_VPWR_c_168_n 0.0052072f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_62 N_A_c_64_n N_VPWR_c_168_n 0.004751f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_63 N_A_c_65_n N_VPWR_c_169_n 0.00570803f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A_c_64_n N_VPWR_c_170_n 0.00597712f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_c_65_n N_VPWR_c_170_n 0.00673617f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_c_60_n N_VPWR_c_162_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_c_61_n N_VPWR_c_162_n 0.0118438f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A_c_62_n N_VPWR_c_162_n 0.00999457f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_c_63_n N_VPWR_c_162_n 0.0118438f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_c_64_n N_VPWR_c_162_n 0.00999457f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A_c_65_n N_VPWR_c_162_n 0.0131262f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_c_60_n N_Y_c_227_n 0.00347232f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A_c_61_n N_Y_c_227_n 5.79575e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 A N_Y_c_227_n 0.0253353f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_c_59_n N_Y_c_227_n 0.00651614f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_76 N_A_c_60_n N_Y_c_231_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_c_61_n N_Y_c_231_n 0.0106251f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_c_62_n N_Y_c_231_n 6.24674e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_c_53_n N_Y_c_234_n 0.00504502f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_c_53_n N_Y_c_219_n 0.0126725f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_c_54_n N_Y_c_219_n 0.0131218f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_82 A N_Y_c_219_n 0.0557164f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A_c_59_n N_Y_c_219_n 0.00369961f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_84 N_A_c_52_n N_Y_c_220_n 0.00138578f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_85 A N_Y_c_220_n 0.0140163f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_c_59_n N_Y_c_220_n 0.0033272f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_87 N_A_c_61_n N_Y_c_242_n 0.0137916f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_c_62_n N_Y_c_242_n 0.0101048f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_89 A N_Y_c_242_n 0.0356113f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A_c_59_n N_Y_c_242_n 0.00635951f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_91 N_A_c_61_n N_Y_c_246_n 6.48386e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_c_62_n N_Y_c_246_n 0.0130707f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A_c_63_n N_Y_c_246_n 0.0106081f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_c_64_n N_Y_c_246_n 6.26411e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_c_55_n N_Y_c_250_n 0.00504502f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_c_55_n N_Y_c_221_n 0.0131218f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_c_56_n N_Y_c_221_n 0.0131218f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_98 A N_Y_c_221_n 0.0682828f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_99 N_A_c_59_n N_Y_c_221_n 0.00369961f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_100 N_A_c_63_n N_Y_c_255_n 5.85735e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_64_n N_Y_c_255_n 0.0128705f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_c_65_n N_Y_c_255_n 0.0253519f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_57_n N_Y_c_258_n 0.00449507f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_c_62_n N_Y_c_259_n 0.00210477f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_c_63_n N_Y_c_259_n 5.79575e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_106 A N_Y_c_259_n 0.0253353f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_107 N_A_c_59_n N_Y_c_259_n 0.00651614f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_108 A N_Y_c_222_n 0.0140163f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_109 N_A_c_59_n N_Y_c_222_n 0.0033272f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_110 N_A_c_64_n Y 4.02863e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_56_n Y 4.70607e-19 $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_c_65_n Y 0.00386107f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_c_57_n Y 0.00414834f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_114 A Y 0.0200758f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A_c_59_n Y 0.0209959f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_116 N_A_c_57_n Y 0.0135152f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A_c_59_n Y 0.00350525f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_118 N_A_c_63_n N_Y_c_273_n 0.0137916f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_64_n N_Y_c_273_n 0.0101048f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_120 A N_Y_c_273_n 0.0551661f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A_c_59_n N_Y_c_273_n 0.00635951f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_122 N_A_c_64_n Y 0.00267709f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_c_65_n Y 0.0174335f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_59_n Y 0.00638266f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_125 N_A_c_52_n N_VGND_c_328_n 0.00451231f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_126 A N_VGND_c_328_n 0.00350557f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_127 N_A_c_59_n N_VGND_c_328_n 0.00214651f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_128 N_A_c_52_n N_VGND_c_329_n 0.00585385f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_c_53_n N_VGND_c_329_n 0.00437852f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_53_n N_VGND_c_330_n 0.00276126f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_54_n N_VGND_c_330_n 0.00405406f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_54_n N_VGND_c_331_n 0.00437852f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_55_n N_VGND_c_331_n 0.00437852f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_55_n N_VGND_c_332_n 0.00276126f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_56_n N_VGND_c_332_n 0.00267891f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_c_56_n N_VGND_c_333_n 6.15983e-19 $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_57_n N_VGND_c_333_n 0.0119564f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_c_56_n N_VGND_c_334_n 0.00437852f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_c_57_n N_VGND_c_334_n 0.00203537f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_c_52_n N_VGND_c_336_n 0.0116629f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_c_53_n N_VGND_c_336_n 0.00614065f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_c_54_n N_VGND_c_336_n 0.00626341f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_c_55_n N_VGND_c_336_n 0.00614065f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_c_56_n N_VGND_c_336_n 0.00626341f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_57_n N_VGND_c_336_n 0.0028209f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_146 N_VPWR_c_162_n N_Y_M1000_s 0.00231261f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_147 N_VPWR_c_162_n N_Y_M1003_s 0.00231261f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_148 N_VPWR_c_162_n N_Y_M1007_s 0.00231261f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_149 N_VPWR_c_164_n N_Y_c_227_n 0.0133617f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_150 N_VPWR_c_164_n N_Y_c_231_n 0.0596857f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_151 N_VPWR_c_165_n N_Y_c_231_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_152 N_VPWR_c_166_n N_Y_c_231_n 0.0385613f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_153 N_VPWR_c_162_n N_Y_c_231_n 0.0140101f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_M1002_d N_Y_c_242_n 0.00325884f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_155 N_VPWR_c_166_n N_Y_c_242_n 0.0136682f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_156 N_VPWR_c_166_n N_Y_c_246_n 0.0470327f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_157 N_VPWR_c_167_n N_Y_c_246_n 0.0223557f $X=2.055 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_c_168_n N_Y_c_246_n 0.0385613f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_159 N_VPWR_c_162_n N_Y_c_246_n 0.0140101f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_160 N_VPWR_c_168_n N_Y_c_255_n 0.0470327f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_161 N_VPWR_c_169_n N_Y_c_255_n 0.0177504f $X=3.08 $Y=2.34 $X2=0 $Y2=0
cc_162 N_VPWR_c_170_n N_Y_c_255_n 0.0223557f $X=2.995 $Y=2.72 $X2=0 $Y2=0
cc_163 N_VPWR_c_162_n N_Y_c_255_n 0.0140101f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_164 N_VPWR_M1010_d Y 6.97377e-19 $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_165 N_VPWR_M1004_d N_Y_c_273_n 0.00325884f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_166 N_VPWR_c_168_n N_Y_c_273_n 0.0136682f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_167 N_VPWR_M1010_d Y 0.00663034f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_168 N_VPWR_c_169_n Y 0.00623505f $X=3.08 $Y=2.34 $X2=0 $Y2=0
cc_169 N_Y_c_219_n N_VGND_M1005_d 0.00255004f $X=1.585 $Y=0.815 $X2=0 $Y2=0
cc_170 N_Y_c_221_n N_VGND_M1008_d 0.00255004f $X=2.525 $Y=0.815 $X2=0 $Y2=0
cc_171 Y N_VGND_M1011_d 0.00345704f $X=3.085 $Y=0.85 $X2=0 $Y2=0
cc_172 N_Y_c_234_n N_VGND_c_329_n 0.0115672f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_173 N_Y_c_219_n N_VGND_c_329_n 0.00345617f $X=1.585 $Y=0.815 $X2=0 $Y2=0
cc_174 N_Y_c_219_n N_VGND_c_330_n 0.0121134f $X=1.585 $Y=0.815 $X2=0 $Y2=0
cc_175 N_Y_c_219_n N_VGND_c_331_n 0.00346295f $X=1.585 $Y=0.815 $X2=0 $Y2=0
cc_176 N_Y_c_250_n N_VGND_c_331_n 0.0115672f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_177 N_Y_c_221_n N_VGND_c_331_n 0.00345617f $X=2.525 $Y=0.815 $X2=0 $Y2=0
cc_178 N_Y_c_221_n N_VGND_c_332_n 0.0121134f $X=2.525 $Y=0.815 $X2=0 $Y2=0
cc_179 N_Y_c_258_n N_VGND_c_333_n 0.0216214f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_180 Y N_VGND_c_333_n 0.0180302f $X=3.085 $Y=0.85 $X2=0 $Y2=0
cc_181 N_Y_c_221_n N_VGND_c_334_n 0.00548535f $X=2.525 $Y=0.815 $X2=0 $Y2=0
cc_182 N_Y_c_258_n N_VGND_c_334_n 0.011304f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_183 Y N_VGND_c_335_n 0.00148445f $X=3.085 $Y=0.85 $X2=0 $Y2=0
cc_184 N_Y_M1001_s N_VGND_c_336_n 0.00477343f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_185 N_Y_M1006_s N_VGND_c_336_n 0.00327321f $X=1.535 $Y=0.235 $X2=0 $Y2=0
cc_186 N_Y_M1009_s N_VGND_c_336_n 0.00331787f $X=2.475 $Y=0.235 $X2=0 $Y2=0
cc_187 N_Y_c_234_n N_VGND_c_336_n 0.0064623f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_188 N_Y_c_219_n N_VGND_c_336_n 0.0149247f $X=1.585 $Y=0.815 $X2=0 $Y2=0
cc_189 N_Y_c_250_n N_VGND_c_336_n 0.0064623f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_190 N_Y_c_221_n N_VGND_c_336_n 0.0191258f $X=2.525 $Y=0.815 $X2=0 $Y2=0
cc_191 N_Y_c_258_n N_VGND_c_336_n 0.00640911f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_192 Y N_VGND_c_336_n 0.0038121f $X=3.085 $Y=0.85 $X2=0 $Y2=0
