* File: sky130_fd_sc_hdll__or4b_2.pex.spice
* Created: Thu Aug 27 19:25:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR4B_2%D_N 1 3 6 8 13
c28 6 0 3.04036e-19 $X=0.52 $Y=0.445
c29 1 0 2.19607e-19 $X=0.495 $Y=1.41
r30 13 14 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r31 11 13 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r33 4 14 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r35 1 13 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r36 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_2%A_186_21# 1 2 3 10 12 13 15 16 18 19 21 22
+ 28 30 34 38 39 41 43 44
c118 44 0 3.00167e-19 $X=3.525 $Y=1.612
c119 39 0 1.66962e-19 $X=1.49 $Y=1.16
c120 19 0 1.40478e-19 $X=1.5 $Y=1.41
r121 47 48 57.0452 $w=3.76e-07 $l=4.45e-07 $layer=POLY_cond $X=1.03 $Y=1.202
+ $X2=1.475 $Y2=1.202
r122 46 47 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=1.005 $Y=1.202
+ $X2=1.03 $Y2=1.202
r123 43 44 10.1862 $w=3.33e-07 $l=2.15e-07 $layer=LI1_cond $X=3.74 $Y=1.612
+ $X2=3.525 $Y2=1.612
r124 39 50 1.28191 $w=3.76e-07 $l=1e-08 $layer=POLY_cond $X=1.49 $Y=1.202
+ $X2=1.5 $Y2=1.202
r125 39 48 1.92287 $w=3.76e-07 $l=1.5e-08 $layer=POLY_cond $X=1.49 $Y=1.202
+ $X2=1.475 $Y2=1.202
r126 38 40 18.2016 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=1.16
+ $X2=1.57 $Y2=1.53
r127 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.16 $X2=1.49 $Y2=1.16
r128 36 38 18.4476 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=1.57 $Y=0.785
+ $X2=1.57 $Y2=1.16
r129 32 34 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.22 $Y=0.7
+ $X2=3.22 $Y2=0.47
r130 31 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=0.785
+ $X2=2.27 $Y2=0.785
r131 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.135 $Y=0.785
+ $X2=3.22 $Y2=0.7
r132 30 31 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.135 $Y=0.785
+ $X2=2.355 $Y2=0.785
r133 26 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.27 $Y=0.7 $X2=2.27
+ $Y2=0.785
r134 26 28 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.27 $Y=0.7
+ $X2=2.27 $Y2=0.47
r135 25 40 2.94836 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=1.53
+ $X2=1.57 $Y2=1.53
r136 25 44 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=1.735 $Y=1.53
+ $X2=3.525 $Y2=1.53
r137 23 36 2.94836 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=0.785
+ $X2=1.57 $Y2=0.785
r138 22 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=0.785
+ $X2=2.27 $Y2=0.785
r139 22 23 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.185 $Y=0.785
+ $X2=1.735 $Y2=0.785
r140 19 50 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.5 $Y2=1.202
r141 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.5 $Y2=1.985
r142 16 48 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=1.202
r143 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=0.56
r144 13 47 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.202
r145 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.985
r146 10 46 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=1.202
r147 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.56
r148 3 43 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=3.595
+ $Y=1.485 $X2=3.74 $Y2=1.655
r149 2 34 182 $w=1.7e-07 $l=3.14166e-07 $layer=licon1_NDIFF $count=1 $X=3.035
+ $Y=0.235 $X2=3.22 $Y2=0.47
r150 1 28 182 $w=1.7e-07 $l=3.14166e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.235 $X2=2.27 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_2%A 3 5 7 8 15
c35 8 0 1.93068e-19 $X=2.185 $Y=1.105
r36 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=1.16 $X2=2.07 $Y2=1.16
r37 8 15 11.0909 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=2.27 $Y=1.175 $X2=2.07
+ $Y2=1.175
r38 5 11 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.035 $Y=1.41
+ $X2=2.095 $Y2=1.16
r39 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.035 $Y=1.41
+ $X2=2.035 $Y2=1.695
r40 1 11 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.01 $Y=0.995
+ $X2=2.095 $Y2=1.16
r41 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.01 $Y=0.995 $X2=2.01
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_2%B 3 6 8 10 11 20
c42 10 0 1.50083e-19 $X=2.56 $Y=1.41
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=2.3 $X2=2.48 $Y2=2.3
r44 11 20 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=2.78 $Y=2.27
+ $X2=2.785 $Y2=2.27
r45 11 15 11.9218 $w=2.88e-07 $l=3e-07 $layer=LI1_cond $X=2.78 $Y=2.27 $X2=2.48
+ $Y2=2.27
r46 9 10 35.1901 $w=1.8e-07 $l=8.5e-08 $layer=POLY_cond $X=2.56 $Y=1.325
+ $X2=2.56 $Y2=1.41
r47 8 10 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.565 $Y=1.695
+ $X2=2.565 $Y2=1.41
r48 6 14 50.163 $w=3.01e-07 $l=3.00167e-07 $layer=POLY_cond $X=2.565 $Y=2.035
+ $X2=2.49 $Y2=2.3
r49 6 8 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=2.565 $Y=2.035
+ $X2=2.565 $Y2=1.695
r50 3 9 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.54 $Y=0.445 $X2=2.54
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_2%C 3 5 7 8 9 20
c32 5 0 1.93068e-19 $X=2.985 $Y=1.41
r33 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.02
+ $Y=1.16 $X2=3.02 $Y2=1.16
r34 9 20 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=3.8 $Y=1.175
+ $X2=3.785 $Y2=1.175
r35 8 20 27.45 $w=1.98e-07 $l=4.95e-07 $layer=LI1_cond $X=3.29 $Y=1.175
+ $X2=3.785 $Y2=1.175
r36 8 14 14.9727 $w=1.98e-07 $l=2.7e-07 $layer=LI1_cond $X=3.29 $Y=1.175
+ $X2=3.02 $Y2=1.175
r37 5 13 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=3.02 $Y2=1.16
r38 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=2.985 $Y2=1.695
r39 1 13 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.96 $Y=0.995
+ $X2=3.02 $Y2=1.16
r40 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.96 $Y=0.995 $X2=2.96
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_2%A_27_47# 1 2 9 12 14 16 19 21 25 26 29 31
+ 34 35 37 41 44
c112 44 0 1.66962e-19 $X=1.702 $Y=1.87
c113 31 0 1.40478e-19 $X=3.16 $Y=1.87
c114 29 0 3.79655e-20 $X=1.54 $Y=2.08
c115 16 0 1.50083e-19 $X=3.5 $Y=1.41
r116 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=2.3 $X2=3.44 $Y2=2.3
r117 35 37 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.33 $Y=2.3
+ $X2=3.44 $Y2=2.3
r118 34 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=2.215
+ $X2=3.33 $Y2=2.3
r119 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.245 $Y=1.955
+ $X2=3.245 $Y2=2.215
r120 32 44 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=1.865 $Y=1.87
+ $X2=1.702 $Y2=1.87
r121 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.16 $Y=1.87
+ $X2=3.245 $Y2=1.955
r122 31 32 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=3.16 $Y=1.87
+ $X2=1.865 $Y2=1.87
r123 30 42 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.815 $Y=2.08
+ $X2=0.662 $Y2=2.08
r124 29 44 7.44655 $w=3.23e-07 $l=2.1e-07 $layer=LI1_cond $X=1.702 $Y=2.08
+ $X2=1.702 $Y2=1.87
r125 29 30 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.54 $Y=2.08
+ $X2=0.815 $Y2=2.08
r126 27 41 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.73 $Y=0.905
+ $X2=0.73 $Y2=1.605
r127 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.73 $Y2=0.905
r128 25 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.35 $Y2=0.82
r129 21 42 12.5824 $w=3.03e-07 $l=3.33e-07 $layer=LI1_cond $X=0.662 $Y=1.747
+ $X2=0.662 $Y2=2.08
r130 21 41 7.60552 $w=3.03e-07 $l=1.42e-07 $layer=LI1_cond $X=0.662 $Y=1.747
+ $X2=0.662 $Y2=1.605
r131 21 23 10.1091 $w=2.83e-07 $l=2.5e-07 $layer=LI1_cond $X=0.51 $Y=1.747
+ $X2=0.26 $Y2=1.747
r132 17 26 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.217 $Y=0.735
+ $X2=0.35 $Y2=0.82
r133 17 19 10.2198 $w=2.63e-07 $l=2.35e-07 $layer=LI1_cond $X=0.217 $Y=0.735
+ $X2=0.217 $Y2=0.5
r134 15 16 35.1901 $w=1.8e-07 $l=8.5e-08 $layer=POLY_cond $X=3.5 $Y=1.325
+ $X2=3.5 $Y2=1.41
r135 14 16 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.505 $Y=1.695
+ $X2=3.505 $Y2=1.41
r136 12 38 50.8629 $w=2.91e-07 $l=2.97061e-07 $layer=POLY_cond $X=3.505 $Y=2.035
+ $X2=3.437 $Y2=2.3
r137 12 14 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=3.505 $Y=2.035
+ $X2=3.505 $Y2=1.695
r138 9 15 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.48 $Y=0.445
+ $X2=3.48 $Y2=1.325
r139 2 23 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.72
r140 1 19 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_2%VPWR 1 2 8 11 14 16 29 30 33
r51 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 33 36 9.09823 $w=3.78e-07 $l=3e-07 $layer=LI1_cond $X=0.705 $Y=2.42
+ $X2=0.705 $Y2=2.72
r53 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r54 27 30 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.91 $Y2=2.72
r55 26 29 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.91 $Y2=2.72
r56 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 24 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 24 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 21 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r61 21 23 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 16 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r63 16 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 14 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 14 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r66 12 26 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.965 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 11 23 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.63 $Y=2.72 $X2=1.61
+ $Y2=2.72
r68 11 12 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.797 $Y=2.72
+ $X2=1.965 $Y2=2.72
r69 8 11 10.3204 $w=3.33e-07 $l=3e-07 $layer=LI1_cond $X=1.797 $Y=2.42 $X2=1.797
+ $Y2=2.72
r70 2 8 600 $w=1.7e-07 $l=1.03469e-06 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.485 $X2=1.8 $Y2=2.42
r71 1 33 600 $w=1.7e-07 $l=3.17884e-07 $layer=licon1_PDIFF $count=1 $X=0.535
+ $Y=2.185 $X2=0.73 $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_2%X 1 2 8 10 14 16
c27 14 0 1.81642e-19 $X=1.265 $Y=1.66
c28 10 0 1.38594e-19 $X=1.185 $Y=0.79
c29 8 0 1.65442e-19 $X=1.127 $Y=1.495
r30 11 14 4.81931 $w=3.28e-07 $l=1.38e-07 $layer=LI1_cond $X=1.127 $Y=1.66
+ $X2=1.265 $Y2=1.66
r31 9 16 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.185 $Y=0.625
+ $X2=1.185 $Y2=0.51
r32 9 10 7.16023 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=0.625
+ $X2=1.185 $Y2=0.79
r33 8 11 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=1.127 $Y=1.495
+ $X2=1.127 $Y2=1.66
r34 8 10 37.7894 $w=2.13e-07 $l=7.05e-07 $layer=LI1_cond $X=1.127 $Y=1.495
+ $X2=1.127 $Y2=0.79
r35 2 14 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.66
r36 1 16 182 $w=1.7e-07 $l=3.60832e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_2%VGND 1 2 3 4 17 19 23 25 27 30 31 32 38 43
+ 47 54 56
r72 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r73 47 50 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=1.75 $Y=0 $X2=1.75
+ $Y2=0.4
r74 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r75 44 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r76 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r77 41 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r78 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r79 38 53 4.94378 $w=1.7e-07 $l=3.07e-07 $layer=LI1_cond $X=3.525 $Y=0 $X2=3.832
+ $Y2=0
r80 38 40 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.525 $Y=0 $X2=3.45
+ $Y2=0
r81 37 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r82 37 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r83 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r84 34 47 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=1.75
+ $Y2=0
r85 34 36 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=2.53
+ $Y2=0
r86 32 44 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r87 32 56 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r88 30 36 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.53
+ $Y2=0
r89 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.75
+ $Y2=0
r90 29 40 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.45
+ $Y2=0
r91 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.75
+ $Y2=0
r92 25 53 3.25291 $w=3.8e-07 $l=1.53734e-07 $layer=LI1_cond $X=3.715 $Y=0.085
+ $X2=3.832 $Y2=0
r93 25 27 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=3.715 $Y=0.085
+ $X2=3.715 $Y2=0.5
r94 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=0.085
+ $X2=2.75 $Y2=0
r95 21 23 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.75 $Y=0.085
+ $X2=2.75 $Y2=0.4
r96 20 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=0 $X2=0.765
+ $Y2=0
r97 19 47 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.75
+ $Y2=0
r98 19 20 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=0.85
+ $Y2=0
r99 15 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0
r100 15 17 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0.4
r101 4 27 182 $w=1.7e-07 $l=3.45326e-07 $layer=licon1_NDIFF $count=1 $X=3.555
+ $Y=0.235 $X2=3.74 $Y2=0.5
r102 3 23 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.235 $X2=2.75 $Y2=0.4
r103 2 50 182 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.235 $X2=1.75 $Y2=0.4
r104 1 17 182 $w=1.7e-07 $l=2.38642e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.765 $Y2=0.4
.ends

