* File: sky130_fd_sc_hdll__o21ai_2.pxi.spice
* Created: Wed Sep  2 08:43:31 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21AI_2%A1 N_A1_c_57_n N_A1_M1002_g N_A1_c_58_n
+ N_A1_M1000_g N_A1_c_59_n N_A1_M1005_g N_A1_c_60_n N_A1_M1008_g N_A1_c_64_n
+ N_A1_c_61_n A1 A1 PM_SKY130_FD_SC_HDLL__O21AI_2%A1
x_PM_SKY130_FD_SC_HDLL__O21AI_2%A2 N_A2_c_131_n N_A2_M1003_g N_A2_c_127_n
+ N_A2_M1009_g N_A2_c_132_n N_A2_M1007_g N_A2_c_128_n N_A2_M1010_g A2
+ N_A2_c_129_n N_A2_c_130_n A2 PM_SKY130_FD_SC_HDLL__O21AI_2%A2
x_PM_SKY130_FD_SC_HDLL__O21AI_2%B1 N_B1_c_178_n N_B1_M1004_g N_B1_c_179_n
+ N_B1_c_186_n N_B1_M1001_g N_B1_c_180_n N_B1_c_181_n N_B1_M1006_g N_B1_c_187_n
+ N_B1_M1011_g N_B1_c_182_n N_B1_c_183_n B1 B1 N_B1_c_185_n B1 B1
+ PM_SKY130_FD_SC_HDLL__O21AI_2%B1
x_PM_SKY130_FD_SC_HDLL__O21AI_2%VPWR N_VPWR_M1002_s N_VPWR_M1005_s
+ N_VPWR_M1011_s N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n
+ N_VPWR_c_238_n VPWR N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n
+ N_VPWR_c_233_n PM_SKY130_FD_SC_HDLL__O21AI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O21AI_2%A_120_297# N_A_120_297#_M1002_d
+ N_A_120_297#_M1007_d N_A_120_297#_c_290_n N_A_120_297#_c_291_n
+ N_A_120_297#_c_298_n N_A_120_297#_c_293_n
+ PM_SKY130_FD_SC_HDLL__O21AI_2%A_120_297#
x_PM_SKY130_FD_SC_HDLL__O21AI_2%Y N_Y_M1004_d N_Y_M1003_s N_Y_M1001_d
+ N_Y_c_319_n Y Y Y Y N_Y_c_311_n Y Y N_Y_c_308_n Y N_Y_c_315_n
+ PM_SKY130_FD_SC_HDLL__O21AI_2%Y
x_PM_SKY130_FD_SC_HDLL__O21AI_2%A_29_47# N_A_29_47#_M1000_d N_A_29_47#_M1009_d
+ N_A_29_47#_M1008_d N_A_29_47#_M1006_s N_A_29_47#_c_353_n N_A_29_47#_c_358_n
+ N_A_29_47#_c_354_n N_A_29_47#_c_362_n N_A_29_47#_c_355_n N_A_29_47#_c_367_n
+ N_A_29_47#_c_368_n N_A_29_47#_c_384_n N_A_29_47#_c_356_n N_A_29_47#_c_357_n
+ PM_SKY130_FD_SC_HDLL__O21AI_2%A_29_47#
x_PM_SKY130_FD_SC_HDLL__O21AI_2%VGND N_VGND_M1000_s N_VGND_M1010_s
+ N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n N_VGND_c_425_n VGND
+ N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n
+ PM_SKY130_FD_SC_HDLL__O21AI_2%VGND
cc_1 VNB N_A1_c_57_n 0.0502326f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.41
cc_2 VNB N_A1_c_58_n 0.0197439f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.96
cc_3 VNB N_A1_c_59_n 0.0263665f $X=-0.19 $Y=-0.24 $X2=2.02 $Y2=1.41
cc_4 VNB N_A1_c_60_n 0.017934f $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=0.995
cc_5 VNB N_A1_c_61_n 0.00505416f $X=-0.19 $Y=-0.24 $X2=2.015 $Y2=1.16
cc_6 VNB N_A2_c_127_n 0.0173119f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.96
cc_7 VNB N_A2_c_128_n 0.0181744f $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=0.995
cc_8 VNB N_A2_c_129_n 0.005399f $X=-0.19 $Y=-0.24 $X2=2.022 $Y2=1.53
cc_9 VNB N_A2_c_130_n 0.0398859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B1_c_178_n 0.0149577f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.41
cc_11 VNB N_B1_c_179_n 0.00760459f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.56
cc_12 VNB N_B1_c_180_n 0.0132857f $X=-0.19 $Y=-0.24 $X2=2.02 $Y2=1.985
cc_13 VNB N_B1_c_181_n 0.017933f $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=0.56
cc_14 VNB N_B1_c_182_n 0.00794252f $X=-0.19 $Y=-0.24 $X2=2.015 $Y2=1.16
cc_15 VNB N_B1_c_183_n 0.0114381f $X=-0.19 $Y=-0.24 $X2=2.022 $Y2=1.53
cc_16 VNB B1 0.0217359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B1_c_185_n 0.0332966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_233_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_308_n 0.00290144f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.445
cc_20 VNB N_A_29_47#_c_353_n 0.018052f $X=-0.19 $Y=-0.24 $X2=2.022 $Y2=1.16
cc_21 VNB N_A_29_47#_c_354_n 0.00939546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_29_47#_c_355_n 0.00429425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_29_47#_c_356_n 0.00157304f $X=-0.19 $Y=-0.24 $X2=2.04 $Y2=1.16
cc_24 VNB N_A_29_47#_c_357_n 0.0133315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_422_n 0.00472864f $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=0.56
cc_26 VNB N_VGND_c_423_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=2.022 $Y2=1.16
cc_27 VNB N_VGND_c_424_n 0.0212061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_425_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=2.022 $Y2=1.53
cc_29 VNB N_VGND_c_426_n 0.0459305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_427_n 0.201981f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_31 VNB N_VGND_c_428_n 0.0225816f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.445
cc_32 VPB N_A1_c_57_n 0.0347837f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_33 VPB N_A1_c_59_n 0.0277137f $X=-0.19 $Y=1.305 $X2=2.02 $Y2=1.41
cc_34 VPB N_A1_c_64_n 0.00751513f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.53
cc_35 VPB N_A1_c_61_n 0.00313036f $X=-0.19 $Y=1.305 $X2=2.015 $Y2=1.16
cc_36 VPB A1 0.00518033f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_37 VPB A1 0.00726806f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.445
cc_38 VPB N_A2_c_131_n 0.0161434f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_39 VPB N_A2_c_132_n 0.0166599f $X=-0.19 $Y=1.305 $X2=2.02 $Y2=1.41
cc_40 VPB N_A2_c_130_n 0.0218533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_B1_c_186_n 0.023275f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=0.56
cc_42 VPB N_B1_c_187_n 0.0207798f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.53
cc_43 VPB N_B1_c_183_n 0.00662917f $X=-0.19 $Y=1.305 $X2=2.022 $Y2=1.53
cc_44 VPB B1 0.00787477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_B1_c_185_n 0.0161094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_234_n 0.0107179f $X=-0.19 $Y=1.305 $X2=2.085 $Y2=0.995
cc_47 VPB N_VPWR_c_235_n 0.0306206f $X=-0.19 $Y=1.305 $X2=2.085 $Y2=0.56
cc_48 VPB N_VPWR_c_236_n 0.00297154f $X=-0.19 $Y=1.305 $X2=2.015 $Y2=1.16
cc_49 VPB N_VPWR_c_237_n 0.0117652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_238_n 0.039619f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_239_n 0.0372076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_240_n 0.0216916f $X=-0.19 $Y=1.305 $X2=2.04 $Y2=1.16
cc_53 VPB N_VPWR_c_241_n 0.00591924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_233_n 0.0457802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_Y_c_308_n 0.00165722f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.445
cc_56 N_A1_c_57_n N_A2_c_131_n 0.0214937f $X=0.51 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_57 N_A1_c_64_n N_A2_c_131_n 0.0174357f $X=1.75 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_58 N_A1_c_58_n N_A2_c_127_n 0.0212261f $X=0.535 $Y=0.96 $X2=0 $Y2=0
cc_59 N_A1_c_59_n N_A2_c_132_n 0.0340265f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A1_c_64_n N_A2_c_132_n 0.011627f $X=1.75 $Y=1.53 $X2=0 $Y2=0
cc_61 N_A1_c_61_n N_A2_c_132_n 0.00114406f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A1_c_60_n N_A2_c_128_n 0.0182248f $X=2.085 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A1_c_57_n N_A2_c_129_n 0.00179314f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A1_c_59_n N_A2_c_129_n 2.10609e-19 $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A1_c_64_n N_A2_c_129_n 0.0643732f $X=1.75 $Y=1.53 $X2=0 $Y2=0
cc_66 N_A1_c_61_n N_A2_c_129_n 0.016536f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_67 A1 N_A2_c_129_n 0.0137629f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A1_c_57_n N_A2_c_130_n 0.0269456f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A1_c_59_n N_A2_c_130_n 0.0189272f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A1_c_64_n N_A2_c_130_n 0.0100673f $X=1.75 $Y=1.53 $X2=0 $Y2=0
cc_71 N_A1_c_61_n N_A2_c_130_n 0.0044123f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_72 A1 N_A2_c_130_n 9.42695e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_73 N_A1_c_60_n N_B1_c_178_n 0.0118108f $X=2.085 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_74 N_A1_c_59_n N_B1_c_186_n 0.0343275f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A1_c_61_n N_B1_c_186_n 0.00216394f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A1_c_59_n N_B1_c_182_n 0.0215846f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A1_c_61_n N_B1_c_182_n 0.00332146f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_78 A1 N_VPWR_M1002_s 0.00302366f $X=0.14 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_79 N_A1_c_61_n N_VPWR_M1005_s 0.00300391f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A1_c_57_n N_VPWR_c_235_n 0.0149911f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_81 A1 N_VPWR_c_235_n 0.0228119f $X=0.14 $Y=1.445 $X2=0 $Y2=0
cc_82 N_A1_c_59_n N_VPWR_c_236_n 0.0106655f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A1_c_57_n N_VPWR_c_239_n 0.00642146f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A1_c_59_n N_VPWR_c_239_n 0.00382138f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A1_c_57_n N_VPWR_c_233_n 0.0107572f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A1_c_59_n N_VPWR_c_233_n 0.00474159f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A1_c_64_n N_A_120_297#_M1002_d 0.00197722f $X=1.75 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_88 N_A1_c_64_n N_A_120_297#_M1007_d 0.00172995f $X=1.75 $Y=1.53 $X2=0 $Y2=0
cc_89 N_A1_c_61_n N_A_120_297#_M1007_d 0.0016577f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A1_c_64_n N_A_120_297#_c_290_n 0.0151327f $X=1.75 $Y=1.53 $X2=0 $Y2=0
cc_91 N_A1_c_64_n N_Y_M1003_s 0.00198204f $X=1.75 $Y=1.53 $X2=0 $Y2=0
cc_92 N_A1_c_59_n N_Y_c_311_n 0.015186f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A1_c_61_n N_Y_c_311_n 0.0334652f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A1_c_59_n N_Y_c_308_n 4.13784e-19 $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A1_c_61_n N_Y_c_308_n 0.0253557f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A1_c_59_n N_Y_c_315_n 6.68213e-19 $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A1_c_64_n N_Y_c_315_n 0.0361847f $X=1.75 $Y=1.53 $X2=0 $Y2=0
cc_98 N_A1_c_58_n N_A_29_47#_c_358_n 0.0122325f $X=0.535 $Y=0.96 $X2=0 $Y2=0
cc_99 N_A1_c_64_n N_A_29_47#_c_358_n 0.00498497f $X=1.75 $Y=1.53 $X2=0 $Y2=0
cc_100 N_A1_c_57_n N_A_29_47#_c_354_n 0.00825477f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_101 A1 N_A_29_47#_c_354_n 0.0255131f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_102 N_A1_c_58_n N_A_29_47#_c_362_n 5.79399e-19 $X=0.535 $Y=0.96 $X2=0 $Y2=0
cc_103 N_A1_c_59_n N_A_29_47#_c_355_n 0.00564397f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A1_c_60_n N_A_29_47#_c_355_n 0.0103516f $X=2.085 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A1_c_64_n N_A_29_47#_c_355_n 0.00480305f $X=1.75 $Y=1.53 $X2=0 $Y2=0
cc_106 N_A1_c_61_n N_A_29_47#_c_355_n 0.0356606f $X=2.015 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A1_c_60_n N_A_29_47#_c_367_n 0.00245764f $X=2.085 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A1_c_60_n N_A_29_47#_c_368_n 0.0050626f $X=2.085 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A1_c_58_n N_VGND_c_422_n 0.00274874f $X=0.535 $Y=0.96 $X2=0 $Y2=0
cc_110 N_A1_c_60_n N_VGND_c_423_n 0.00522011f $X=2.085 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A1_c_60_n N_VGND_c_426_n 0.0042335f $X=2.085 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A1_c_58_n N_VGND_c_427_n 0.0070535f $X=0.535 $Y=0.96 $X2=0 $Y2=0
cc_113 N_A1_c_60_n N_VGND_c_427_n 0.00635527f $X=2.085 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A1_c_58_n N_VGND_c_428_n 0.00436487f $X=0.535 $Y=0.96 $X2=0 $Y2=0
cc_115 N_A2_c_131_n N_VPWR_c_235_n 9.73093e-19 $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A2_c_132_n N_VPWR_c_236_n 0.00100104f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A2_c_131_n N_VPWR_c_239_n 0.00429453f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A2_c_132_n N_VPWR_c_239_n 0.00429453f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A2_c_131_n N_VPWR_c_233_n 0.00614026f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A2_c_132_n N_VPWR_c_233_n 0.0063433f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A2_c_131_n N_A_120_297#_c_291_n 0.0143719f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A2_c_132_n N_A_120_297#_c_291_n 0.0113879f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A2_c_132_n N_A_120_297#_c_293_n 0.00411326f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A2_c_132_n N_Y_c_311_n 0.0107806f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A2_c_132_n N_Y_c_315_n 0.00370818f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A2_c_127_n N_A_29_47#_c_358_n 0.00633817f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A2_c_129_n N_A_29_47#_c_358_n 0.0209679f $X=1.35 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A2_c_130_n N_A_29_47#_c_358_n 0.00294319f $X=1.47 $Y=1.202 $X2=0 $Y2=0
cc_129 N_A2_c_127_n N_A_29_47#_c_362_n 0.0083113f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A2_c_128_n N_A_29_47#_c_355_n 0.0109911f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A2_c_129_n N_A_29_47#_c_355_n 0.0101817f $X=1.35 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A2_c_128_n N_A_29_47#_c_368_n 7.28393e-19 $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A2_c_127_n N_A_29_47#_c_356_n 0.00230239f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A2_c_129_n N_A_29_47#_c_356_n 0.0237681f $X=1.35 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A2_c_130_n N_A_29_47#_c_356_n 0.00379646f $X=1.47 $Y=1.202 $X2=0 $Y2=0
cc_136 N_A2_c_127_n N_VGND_c_422_n 0.00358434f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A2_c_128_n N_VGND_c_423_n 0.00408861f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A2_c_127_n N_VGND_c_424_n 0.00398595f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A2_c_128_n N_VGND_c_424_n 0.00436487f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A2_c_127_n N_VGND_c_427_n 0.00589518f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A2_c_128_n N_VGND_c_427_n 0.00652478f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B1_c_186_n N_VPWR_c_236_n 0.00328209f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B1_c_187_n N_VPWR_c_238_n 0.0199662f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_144 B1 N_VPWR_c_238_n 0.0227481f $X=3.3 $Y=0.765 $X2=0 $Y2=0
cc_145 N_B1_c_185_n N_VPWR_c_238_n 0.00149204f $X=3.365 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B1_c_186_n N_VPWR_c_240_n 0.0053025f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B1_c_187_n N_VPWR_c_240_n 0.00430719f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B1_c_186_n N_VPWR_c_233_n 0.00709264f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B1_c_187_n N_VPWR_c_233_n 0.00719535f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B1_c_186_n N_Y_c_319_n 0.0072067f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B1_c_187_n N_Y_c_319_n 0.0140411f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B1_c_187_n Y 0.00392665f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_153 N_B1_c_186_n N_Y_c_311_n 0.0189657f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_154 N_B1_c_178_n N_Y_c_308_n 0.00320852f $X=2.515 $Y=0.96 $X2=0 $Y2=0
cc_155 N_B1_c_179_n N_Y_c_308_n 0.0028639f $X=2.54 $Y=1.31 $X2=0 $Y2=0
cc_156 N_B1_c_186_n N_Y_c_308_n 0.0058249f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_157 N_B1_c_180_n N_Y_c_308_n 0.0130904f $X=2.92 $Y=1.062 $X2=0 $Y2=0
cc_158 N_B1_c_181_n N_Y_c_308_n 0.0133525f $X=2.995 $Y=0.96 $X2=0 $Y2=0
cc_159 N_B1_c_187_n N_Y_c_308_n 0.0144271f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_160 N_B1_c_183_n N_Y_c_308_n 0.0171896f $X=2.92 $Y=0.96 $X2=0 $Y2=0
cc_161 B1 N_Y_c_308_n 0.0448478f $X=3.3 $Y=0.765 $X2=0 $Y2=0
cc_162 B1 N_A_29_47#_M1006_s 0.00387643f $X=3.3 $Y=0.765 $X2=0 $Y2=0
cc_163 N_B1_c_178_n N_A_29_47#_c_355_n 0.00318705f $X=2.515 $Y=0.96 $X2=0 $Y2=0
cc_164 N_B1_c_178_n N_A_29_47#_c_367_n 5.89792e-19 $X=2.515 $Y=0.96 $X2=0 $Y2=0
cc_165 N_B1_c_178_n N_A_29_47#_c_368_n 0.00459058f $X=2.515 $Y=0.96 $X2=0 $Y2=0
cc_166 N_B1_c_181_n N_A_29_47#_c_368_n 7.39444e-19 $X=2.995 $Y=0.96 $X2=0 $Y2=0
cc_167 N_B1_c_178_n N_A_29_47#_c_384_n 0.0107519f $X=2.515 $Y=0.96 $X2=0 $Y2=0
cc_168 N_B1_c_180_n N_A_29_47#_c_384_n 8.91958e-19 $X=2.92 $Y=1.062 $X2=0 $Y2=0
cc_169 N_B1_c_181_n N_A_29_47#_c_384_n 0.0111274f $X=2.995 $Y=0.96 $X2=0 $Y2=0
cc_170 N_B1_c_183_n N_A_29_47#_c_384_n 0.00402622f $X=2.92 $Y=0.96 $X2=0 $Y2=0
cc_171 N_B1_c_181_n N_A_29_47#_c_357_n 0.00660852f $X=2.995 $Y=0.96 $X2=0 $Y2=0
cc_172 B1 N_A_29_47#_c_357_n 0.0205835f $X=3.3 $Y=0.765 $X2=0 $Y2=0
cc_173 N_B1_c_185_n N_A_29_47#_c_357_n 0.0010079f $X=3.365 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B1_c_178_n N_VGND_c_426_n 0.00357842f $X=2.515 $Y=0.96 $X2=0 $Y2=0
cc_175 N_B1_c_181_n N_VGND_c_426_n 0.00357877f $X=2.995 $Y=0.96 $X2=0 $Y2=0
cc_176 N_B1_c_178_n N_VGND_c_427_n 0.00543359f $X=2.515 $Y=0.96 $X2=0 $Y2=0
cc_177 N_B1_c_181_n N_VGND_c_427_n 0.00656954f $X=2.995 $Y=0.96 $X2=0 $Y2=0
cc_178 B1 N_VGND_c_427_n 0.00216432f $X=3.3 $Y=0.765 $X2=0 $Y2=0
cc_179 N_VPWR_c_233_n N_A_120_297#_M1002_d 0.00426758f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_180 N_VPWR_c_233_n N_A_120_297#_M1007_d 0.00330737f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_239_n N_A_120_297#_c_291_n 0.0444999f $X=2.06 $Y=2.72 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_233_n N_A_120_297#_c_291_n 0.0280854f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_239_n N_A_120_297#_c_298_n 0.014286f $X=2.06 $Y=2.72 $X2=0 $Y2=0
cc_184 N_VPWR_c_233_n N_A_120_297#_c_298_n 0.00846213f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_236_n N_A_120_297#_c_293_n 0.0196339f $X=2.275 $Y=2.34 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_239_n N_A_120_297#_c_293_n 0.012523f $X=2.06 $Y=2.72 $X2=0 $Y2=0
cc_187 N_VPWR_c_233_n N_A_120_297#_c_293_n 0.00710678f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_233_n N_Y_M1003_s 0.00240926f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_189 N_VPWR_c_233_n N_Y_M1001_d 0.0027532f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_190 N_VPWR_c_238_n N_Y_c_319_n 0.0386292f $X=3.365 $Y=1.735 $X2=0 $Y2=0
cc_191 N_VPWR_c_240_n N_Y_c_319_n 0.0266734f $X=3.28 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_233_n N_Y_c_319_n 0.0150868f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_238_n Y 0.0145383f $X=3.365 $Y=1.735 $X2=0 $Y2=0
cc_194 N_VPWR_M1005_s N_Y_c_311_n 0.00764918f $X=2.11 $Y=1.485 $X2=0 $Y2=0
cc_195 N_VPWR_c_236_n N_Y_c_311_n 0.0178393f $X=2.275 $Y=2.34 $X2=0 $Y2=0
cc_196 N_VPWR_c_239_n N_Y_c_311_n 0.00217898f $X=2.06 $Y=2.72 $X2=0 $Y2=0
cc_197 N_VPWR_c_240_n N_Y_c_311_n 0.00284211f $X=3.28 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_233_n N_Y_c_311_n 0.0126147f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_238_n N_Y_c_308_n 0.0165884f $X=3.365 $Y=1.735 $X2=0 $Y2=0
cc_200 N_A_120_297#_c_291_n N_Y_M1003_s 0.00372897f $X=1.675 $Y=2.38 $X2=0.51
+ $Y2=1.985
cc_201 N_A_120_297#_M1007_d N_Y_c_311_n 0.00573175f $X=1.56 $Y=1.485 $X2=0 $Y2=0
cc_202 N_A_120_297#_c_291_n N_Y_c_311_n 0.00804752f $X=1.675 $Y=2.38 $X2=0 $Y2=0
cc_203 N_A_120_297#_c_293_n N_Y_c_311_n 0.0139655f $X=1.76 $Y=2.3 $X2=0 $Y2=0
cc_204 N_A_120_297#_c_291_n N_Y_c_315_n 0.0143524f $X=1.675 $Y=2.38 $X2=0 $Y2=0
cc_205 N_Y_c_308_n N_A_29_47#_c_355_n 0.0112777f $X=2.78 $Y=0.76 $X2=0 $Y2=0
cc_206 N_Y_c_308_n N_A_29_47#_c_368_n 0.00748984f $X=2.78 $Y=0.76 $X2=0 $Y2=0
cc_207 N_Y_M1004_d N_A_29_47#_c_384_n 0.00517242f $X=2.59 $Y=0.235 $X2=0 $Y2=0
cc_208 N_Y_c_308_n N_A_29_47#_c_384_n 0.0233868f $X=2.78 $Y=0.76 $X2=0 $Y2=0
cc_209 N_Y_M1004_d N_VGND_c_427_n 0.00265018f $X=2.59 $Y=0.235 $X2=0 $Y2=0
cc_210 N_A_29_47#_c_358_n N_VGND_M1000_s 0.00485811f $X=1.015 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_211 N_A_29_47#_c_355_n N_VGND_M1010_s 0.00979481f $X=2.135 $Y=0.8 $X2=0 $Y2=0
cc_212 N_A_29_47#_c_358_n N_VGND_c_422_n 0.0130378f $X=1.015 $Y=0.8 $X2=0 $Y2=0
cc_213 N_A_29_47#_c_362_n N_VGND_c_422_n 0.0207137f $X=1.23 $Y=0.4 $X2=0 $Y2=0
cc_214 N_A_29_47#_c_355_n N_VGND_c_423_n 0.0131159f $X=2.135 $Y=0.8 $X2=0 $Y2=0
cc_215 N_A_29_47#_c_367_n N_VGND_c_423_n 0.00884087f $X=2.3 $Y=0.425 $X2=0 $Y2=0
cc_216 N_A_29_47#_c_368_n N_VGND_c_423_n 0.00585481f $X=2.3 $Y=0.715 $X2=0 $Y2=0
cc_217 N_A_29_47#_c_358_n N_VGND_c_424_n 0.00217503f $X=1.015 $Y=0.8 $X2=0 $Y2=0
cc_218 N_A_29_47#_c_362_n N_VGND_c_424_n 0.0232119f $X=1.23 $Y=0.4 $X2=0 $Y2=0
cc_219 N_A_29_47#_c_355_n N_VGND_c_424_n 0.00339992f $X=2.135 $Y=0.8 $X2=0 $Y2=0
cc_220 N_A_29_47#_c_355_n N_VGND_c_426_n 0.0037456f $X=2.135 $Y=0.8 $X2=0 $Y2=0
cc_221 N_A_29_47#_c_367_n N_VGND_c_426_n 0.0189784f $X=2.3 $Y=0.425 $X2=0 $Y2=0
cc_222 N_A_29_47#_c_384_n N_VGND_c_426_n 0.0463135f $X=3.28 $Y=0.34 $X2=0 $Y2=0
cc_223 N_A_29_47#_c_357_n N_VGND_c_426_n 0.016642f $X=3.405 $Y=0.34 $X2=0 $Y2=0
cc_224 N_A_29_47#_M1000_d N_VGND_c_427_n 0.00265179f $X=0.145 $Y=0.235 $X2=0
+ $Y2=0
cc_225 N_A_29_47#_M1009_d N_VGND_c_427_n 0.00274151f $X=1.09 $Y=0.235 $X2=0
+ $Y2=0
cc_226 N_A_29_47#_M1008_d N_VGND_c_427_n 0.00223231f $X=2.16 $Y=0.235 $X2=0
+ $Y2=0
cc_227 N_A_29_47#_M1006_s N_VGND_c_427_n 0.00340507f $X=3.07 $Y=0.235 $X2=0
+ $Y2=0
cc_228 N_A_29_47#_c_353_n N_VGND_c_427_n 0.0126066f $X=0.27 $Y=0.4 $X2=0 $Y2=0
cc_229 N_A_29_47#_c_358_n N_VGND_c_427_n 0.0103459f $X=1.015 $Y=0.8 $X2=0 $Y2=0
cc_230 N_A_29_47#_c_362_n N_VGND_c_427_n 0.0141177f $X=1.23 $Y=0.4 $X2=0 $Y2=0
cc_231 N_A_29_47#_c_355_n N_VGND_c_427_n 0.0144381f $X=2.135 $Y=0.8 $X2=0 $Y2=0
cc_232 N_A_29_47#_c_367_n N_VGND_c_427_n 0.0123102f $X=2.3 $Y=0.425 $X2=0 $Y2=0
cc_233 N_A_29_47#_c_384_n N_VGND_c_427_n 0.0291011f $X=3.28 $Y=0.34 $X2=0 $Y2=0
cc_234 N_A_29_47#_c_357_n N_VGND_c_427_n 0.00938745f $X=3.405 $Y=0.34 $X2=0
+ $Y2=0
cc_235 N_A_29_47#_c_353_n N_VGND_c_428_n 0.0219214f $X=0.27 $Y=0.4 $X2=0 $Y2=0
cc_236 N_A_29_47#_c_358_n N_VGND_c_428_n 0.00267476f $X=1.015 $Y=0.8 $X2=0 $Y2=0
