* File: sky130_fd_sc_hdll__o2bb2ai_1.pxi.spice
* Created: Wed Sep  2 08:46:21 2020
* 
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A1_N N_A1_N_c_61_n N_A1_N_M1000_g
+ N_A1_N_c_58_n N_A1_N_M1006_g A1_N N_A1_N_c_60_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A1_N
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A2_N N_A2_N_c_81_n N_A2_N_M1004_g
+ N_A2_N_c_82_n N_A2_N_M1008_g A2_N N_A2_N_c_83_n N_A2_N_c_84_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A2_N
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A_120_297# N_A_120_297#_M1004_d
+ N_A_120_297#_M1000_d N_A_120_297#_c_123_n N_A_120_297#_M1002_g
+ N_A_120_297#_c_117_n N_A_120_297#_M1005_g N_A_120_297#_c_118_n
+ N_A_120_297#_c_119_n N_A_120_297#_c_151_p N_A_120_297#_c_133_n
+ N_A_120_297#_c_135_n N_A_120_297#_c_126_n N_A_120_297#_c_120_n
+ N_A_120_297#_c_121_n N_A_120_297#_c_122_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A_120_297#
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_1%B2 N_B2_c_181_n N_B2_M1007_g N_B2_c_182_n
+ N_B2_M1009_g N_B2_c_183_n B2 PM_SKY130_FD_SC_HDLL__O2BB2AI_1%B2
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_1%B1 N_B1_c_223_n N_B1_M1001_g N_B1_c_226_n
+ N_B1_M1003_g B1 N_B1_c_224_n N_B1_c_225_n PM_SKY130_FD_SC_HDLL__O2BB2AI_1%B1
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_1%VPWR N_VPWR_M1000_s N_VPWR_M1008_d
+ N_VPWR_M1003_d N_VPWR_c_250_n N_VPWR_c_251_n N_VPWR_c_252_n N_VPWR_c_253_n
+ N_VPWR_c_254_n VPWR N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_249_n
+ N_VPWR_c_258_n N_VPWR_c_259_n PM_SKY130_FD_SC_HDLL__O2BB2AI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_1%Y N_Y_M1005_s N_Y_M1002_d N_Y_c_293_n
+ N_Y_c_303_n N_Y_c_295_n Y PM_SKY130_FD_SC_HDLL__O2BB2AI_1%Y
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_1%VGND N_VGND_M1006_s N_VGND_M1009_d
+ N_VGND_c_329_n N_VGND_c_330_n N_VGND_c_331_n VGND N_VGND_c_332_n
+ N_VGND_c_333_n N_VGND_c_334_n N_VGND_c_335_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_1%VGND
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A_396_47# N_A_396_47#_M1005_d
+ N_A_396_47#_M1001_d N_A_396_47#_c_376_n N_A_396_47#_c_373_n
+ N_A_396_47#_c_374_n N_A_396_47#_c_375_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_1%A_396_47#
cc_1 VNB N_A1_N_c_58_n 0.0213679f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.995
cc_2 VNB A1_N 0.0156928f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A1_N_c_60_n 0.0406751f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.202
cc_4 VNB N_A2_N_c_81_n 0.0195988f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.41
cc_5 VNB N_A2_N_c_82_n 0.0209616f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.995
cc_6 VNB N_A2_N_c_83_n 0.00269804f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.202
cc_7 VNB N_A2_N_c_84_n 0.00150095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_120_297#_c_117_n 0.0207951f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_9 VNB N_A_120_297#_c_118_n 0.0289798f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.202
cc_10 VNB N_A_120_297#_c_119_n 0.0133695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_120_297#_c_120_n 0.00879707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_120_297#_c_121_n 0.00701951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_120_297#_c_122_n 0.00236927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B2_c_181_n 0.020245f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.41
cc_15 VNB N_B2_c_182_n 0.0168395f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.995
cc_16 VNB N_B2_c_183_n 0.00493557f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_17 VNB B2 2.49476e-19 $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.202
cc_18 VNB N_B1_c_223_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.41
cc_19 VNB N_B1_c_224_n 0.0424395f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_20 VNB N_B1_c_225_n 0.00789198f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.202
cc_21 VNB N_VPWR_c_249_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_293_n 0.00129211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_329_n 0.0115155f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_24 VNB N_VGND_c_330_n 0.0284516f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.202
cc_25 VNB N_VGND_c_331_n 0.00467422f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.202
cc_26 VNB N_VGND_c_332_n 0.0562662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_333_n 0.0295869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_334_n 0.220202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_335_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_396_47#_c_373_n 0.0153705f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_31 VNB N_A_396_47#_c_374_n 0.00206507f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.202
cc_32 VNB N_A_396_47#_c_375_n 0.0179666f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_A1_N_c_61_n 0.020476f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_34 VPB N_A1_N_c_60_n 0.0197692f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.202
cc_35 VPB N_A2_N_c_82_n 0.0281648f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=0.995
cc_36 VPB N_A2_N_c_83_n 0.00278414f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.202
cc_37 VPB N_A_120_297#_c_123_n 0.0182751f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_38 VPB N_A_120_297#_c_118_n 0.0134344f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.202
cc_39 VPB N_A_120_297#_c_119_n 0.0068042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_120_297#_c_126_n 0.0028476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_120_297#_c_121_n 0.00217316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_B2_c_181_n 0.0243401f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_43 VPB B2 0.00162687f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.202
cc_44 VPB N_B1_c_226_n 0.0204535f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=0.995
cc_45 VPB N_B1_c_224_n 0.019884f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_46 VPB N_VPWR_c_250_n 0.0117686f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_47 VPB N_VPWR_c_251_n 0.00822434f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.202
cc_48 VPB N_VPWR_c_252_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_253_n 0.00757742f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_254_n 0.00816174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_255_n 0.0325453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_256_n 0.0174178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_249_n 0.0606104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_258_n 0.0132428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_259_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_Y_c_293_n 0.00124792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_Y_c_295_n 0.00679585f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 N_A1_N_c_58_n N_A2_N_c_81_n 0.0295378f $X=0.535 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_59 N_A1_N_c_61_n N_A2_N_c_82_n 0.0200829f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A1_N_c_60_n N_A2_N_c_82_n 0.0295378f $X=0.51 $Y=1.202 $X2=0 $Y2=0
cc_61 A1_N N_A2_N_c_83_n 0.0226327f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_62 N_A1_N_c_60_n N_A2_N_c_83_n 0.00992465f $X=0.51 $Y=1.202 $X2=0 $Y2=0
cc_63 N_A1_N_c_58_n N_A2_N_c_84_n 0.0181955f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_64 A1_N N_A2_N_c_84_n 6.63121e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_65 N_A1_N_c_58_n N_A_120_297#_c_120_n 4.13142e-19 $X=0.535 $Y=0.995 $X2=0
+ $Y2=0
cc_66 N_A1_N_c_61_n N_VPWR_c_251_n 0.00606123f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_67 A1_N N_VPWR_c_251_n 0.020778f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A1_N_c_60_n N_VPWR_c_251_n 0.00606334f $X=0.51 $Y=1.202 $X2=0 $Y2=0
cc_69 N_A1_N_c_61_n N_VPWR_c_252_n 0.00702461f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A1_N_c_61_n N_VPWR_c_249_n 0.0133595f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A1_N_c_58_n N_VGND_c_330_n 0.0160492f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_72 A1_N N_VGND_c_330_n 0.0278031f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_73 N_A1_N_c_60_n N_VGND_c_330_n 0.00239594f $X=0.51 $Y=1.202 $X2=0 $Y2=0
cc_74 N_A1_N_c_58_n N_VGND_c_332_n 0.0057945f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_75 N_A1_N_c_58_n N_VGND_c_334_n 0.0115449f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A2_N_c_82_n N_A_120_297#_c_123_n 0.00631184f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A2_N_c_82_n N_A_120_297#_c_118_n 0.0202683f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A2_N_c_83_n N_A_120_297#_c_118_n 3.12322e-19 $X=1.015 $Y=1.16 $X2=0
+ $Y2=0
cc_79 N_A2_N_c_82_n N_A_120_297#_c_119_n 7.92819e-19 $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A2_N_c_82_n N_A_120_297#_c_133_n 0.0195897f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A2_N_c_83_n N_A_120_297#_c_133_n 0.0147715f $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A2_N_c_83_n N_A_120_297#_c_135_n 0.0183514f $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A2_N_c_82_n N_A_120_297#_c_126_n 0.00406803f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A2_N_c_81_n N_A_120_297#_c_120_n 0.00641981f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_85 N_A2_N_c_82_n N_A_120_297#_c_120_n 0.00310147f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A2_N_c_83_n N_A_120_297#_c_120_n 0.00543737f $X=1.015 $Y=1.16 $X2=0
+ $Y2=0
cc_87 N_A2_N_c_82_n N_A_120_297#_c_121_n 0.00202421f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A2_N_c_83_n N_A_120_297#_c_121_n 0.0267416f $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A2_N_c_81_n N_A_120_297#_c_122_n 0.00246602f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_90 N_A2_N_c_84_n N_A_120_297#_c_122_n 0.005333f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A2_N_c_82_n N_VPWR_c_252_n 0.00702461f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A2_N_c_82_n N_VPWR_c_253_n 0.00391982f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A2_N_c_82_n N_VPWR_c_249_n 0.0131729f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A2_N_c_81_n N_VGND_c_332_n 0.00542362f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A2_N_c_84_n N_VGND_c_332_n 0.0115142f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A2_N_c_81_n N_VGND_c_334_n 0.0110558f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A2_N_c_84_n N_VGND_c_334_n 0.00828176f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A2_N_c_84_n A_122_47# 0.00253371f $X=0.715 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_99 N_A_120_297#_c_123_n N_B2_c_181_n 0.00853155f $X=1.88 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_100 N_A_120_297#_c_119_n N_B2_c_181_n 0.024337f $X=1.88 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_101 N_A_120_297#_c_117_n N_B2_c_182_n 0.0237042f $X=1.905 $Y=0.995 $X2=0
+ $Y2=0
cc_102 N_A_120_297#_c_119_n N_B2_c_183_n 0.00142853f $X=1.88 $Y=1.202 $X2=0
+ $Y2=0
cc_103 N_A_120_297#_c_119_n B2 3.7952e-19 $X=1.88 $Y=1.202 $X2=0 $Y2=0
cc_104 N_A_120_297#_c_133_n N_VPWR_M1008_d 0.00980592f $X=1.27 $Y=1.58 $X2=0
+ $Y2=0
cc_105 N_A_120_297#_c_126_n N_VPWR_M1008_d 2.11684e-19 $X=1.355 $Y=1.495 $X2=0
+ $Y2=0
cc_106 N_A_120_297#_c_151_p N_VPWR_c_252_n 0.0149311f $X=0.745 $Y=1.96 $X2=0
+ $Y2=0
cc_107 N_A_120_297#_c_123_n N_VPWR_c_253_n 0.00399885f $X=1.88 $Y=1.41 $X2=0
+ $Y2=0
cc_108 N_A_120_297#_c_118_n N_VPWR_c_253_n 0.00642345f $X=1.78 $Y=1.16 $X2=0
+ $Y2=0
cc_109 N_A_120_297#_c_133_n N_VPWR_c_253_n 0.0268351f $X=1.27 $Y=1.58 $X2=0
+ $Y2=0
cc_110 N_A_120_297#_c_121_n N_VPWR_c_253_n 0.00489511f $X=1.495 $Y=1.16 $X2=0
+ $Y2=0
cc_111 N_A_120_297#_c_123_n N_VPWR_c_255_n 0.00673617f $X=1.88 $Y=1.41 $X2=0
+ $Y2=0
cc_112 N_A_120_297#_M1000_d N_VPWR_c_249_n 0.00370124f $X=0.6 $Y=1.485 $X2=0
+ $Y2=0
cc_113 N_A_120_297#_c_123_n N_VPWR_c_249_n 0.012529f $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_120_297#_c_151_p N_VPWR_c_249_n 0.00955092f $X=0.745 $Y=1.96 $X2=0
+ $Y2=0
cc_115 N_A_120_297#_c_123_n N_Y_c_293_n 0.00168464f $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_120_297#_c_117_n N_Y_c_293_n 0.00717388f $X=1.905 $Y=0.995 $X2=0
+ $Y2=0
cc_117 N_A_120_297#_c_118_n N_Y_c_293_n 0.00566751f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_120_297#_c_119_n N_Y_c_293_n 0.011905f $X=1.88 $Y=1.202 $X2=0 $Y2=0
cc_119 N_A_120_297#_c_126_n N_Y_c_293_n 0.00580501f $X=1.355 $Y=1.495 $X2=0
+ $Y2=0
cc_120 N_A_120_297#_c_120_n N_Y_c_293_n 0.00990191f $X=1.165 $Y=0.39 $X2=0 $Y2=0
cc_121 N_A_120_297#_c_121_n N_Y_c_293_n 0.0223977f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_120_297#_c_117_n N_Y_c_303_n 0.00733714f $X=1.905 $Y=0.995 $X2=0
+ $Y2=0
cc_123 N_A_120_297#_c_118_n N_Y_c_303_n 0.00621802f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_120_297#_c_120_n N_Y_c_303_n 0.0300001f $X=1.165 $Y=0.39 $X2=0 $Y2=0
cc_125 N_A_120_297#_c_123_n N_Y_c_295_n 0.0161195f $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_120_297#_c_119_n N_Y_c_295_n 6.01036e-19 $X=1.88 $Y=1.202 $X2=0 $Y2=0
cc_127 N_A_120_297#_c_126_n N_Y_c_295_n 0.00224979f $X=1.355 $Y=1.495 $X2=0
+ $Y2=0
cc_128 N_A_120_297#_c_123_n Y 0.0145162f $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_120_297#_c_117_n N_VGND_c_332_n 0.00456303f $X=1.905 $Y=0.995 $X2=0
+ $Y2=0
cc_130 N_A_120_297#_c_120_n N_VGND_c_332_n 0.0247545f $X=1.165 $Y=0.39 $X2=0
+ $Y2=0
cc_131 N_A_120_297#_M1004_d N_VGND_c_334_n 0.00210425f $X=1.03 $Y=0.235 $X2=0
+ $Y2=0
cc_132 N_A_120_297#_c_117_n N_VGND_c_334_n 0.00879357f $X=1.905 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_120_297#_c_120_n N_VGND_c_334_n 0.0163948f $X=1.165 $Y=0.39 $X2=0
+ $Y2=0
cc_134 N_A_120_297#_c_117_n N_A_396_47#_c_376_n 0.00213513f $X=1.905 $Y=0.995
+ $X2=0 $Y2=0
cc_135 N_A_120_297#_c_117_n N_A_396_47#_c_374_n 0.00140151f $X=1.905 $Y=0.995
+ $X2=0 $Y2=0
cc_136 N_B2_c_182_n N_B1_c_223_n 0.0229524f $X=2.395 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_137 N_B2_c_181_n N_B1_c_226_n 0.0484622f $X=2.37 $Y=1.41 $X2=0 $Y2=0
cc_138 B2 N_B1_c_226_n 0.00890526f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_139 N_B2_c_181_n N_B1_c_224_n 0.0229524f $X=2.37 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B2_c_183_n N_B1_c_224_n 0.0018113f $X=2.445 $Y=1.175 $X2=0 $Y2=0
cc_141 B2 N_B1_c_224_n 0.00287505f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_142 N_B2_c_183_n N_B1_c_225_n 0.0123516f $X=2.445 $Y=1.175 $X2=0 $Y2=0
cc_143 B2 N_B1_c_225_n 4.85142e-19 $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_144 B2 N_VPWR_c_254_n 0.0221446f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_145 N_B2_c_181_n N_VPWR_c_255_n 0.00681977f $X=2.37 $Y=1.41 $X2=0 $Y2=0
cc_146 B2 N_VPWR_c_255_n 0.00781729f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_147 N_B2_c_181_n N_VPWR_c_249_n 0.012267f $X=2.37 $Y=1.41 $X2=0 $Y2=0
cc_148 B2 N_VPWR_c_249_n 0.0062765f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_149 N_B2_c_181_n N_Y_c_293_n 0.00133866f $X=2.37 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B2_c_182_n N_Y_c_293_n 5.81918e-19 $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B2_c_183_n N_Y_c_293_n 0.0127513f $X=2.445 $Y=1.175 $X2=0 $Y2=0
cc_152 B2 N_Y_c_293_n 0.00461559f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_153 N_B2_c_181_n N_Y_c_295_n 0.00217332f $X=2.37 $Y=1.41 $X2=0 $Y2=0
cc_154 N_B2_c_183_n N_Y_c_295_n 0.00942836f $X=2.445 $Y=1.175 $X2=0 $Y2=0
cc_155 B2 N_Y_c_295_n 0.00912214f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_156 B2 A_492_297# 0.0113049f $X=2.445 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_157 N_B2_c_182_n N_VGND_c_331_n 0.00268723f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_158 N_B2_c_182_n N_VGND_c_332_n 0.00429718f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_159 N_B2_c_182_n N_VGND_c_334_n 0.00601131f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B2_c_182_n N_A_396_47#_c_376_n 0.00473705f $X=2.395 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_B2_c_182_n N_A_396_47#_c_373_n 0.00865583f $X=2.395 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_B2_c_183_n N_A_396_47#_c_373_n 0.0206867f $X=2.445 $Y=1.175 $X2=0 $Y2=0
cc_163 N_B2_c_181_n N_A_396_47#_c_374_n 0.00322706f $X=2.37 $Y=1.41 $X2=0 $Y2=0
cc_164 N_B2_c_182_n N_A_396_47#_c_374_n 0.0019969f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_165 N_B2_c_183_n N_A_396_47#_c_374_n 0.0158983f $X=2.445 $Y=1.175 $X2=0 $Y2=0
cc_166 N_B2_c_182_n N_A_396_47#_c_375_n 5.15568e-19 $X=2.395 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_B1_c_226_n N_VPWR_c_254_n 0.00558657f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_168 N_B1_c_224_n N_VPWR_c_254_n 0.00606334f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_169 N_B1_c_225_n N_VPWR_c_254_n 0.0202873f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B1_c_226_n N_VPWR_c_255_n 0.00702461f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_171 N_B1_c_226_n N_VPWR_c_249_n 0.0137956f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B1_c_223_n N_VGND_c_331_n 0.00268723f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B1_c_223_n N_VGND_c_333_n 0.00424138f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B1_c_223_n N_VGND_c_334_n 0.00707055f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B1_c_223_n N_A_396_47#_c_376_n 4.7333e-19 $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B1_c_223_n N_A_396_47#_c_373_n 0.0135486f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B1_c_224_n N_A_396_47#_c_373_n 0.00913298f $X=2.84 $Y=1.202 $X2=0 $Y2=0
cc_178 N_B1_c_225_n N_A_396_47#_c_373_n 0.0303643f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B1_c_223_n N_A_396_47#_c_375_n 0.00612654f $X=2.815 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_249_n N_Y_M1002_d 0.00264678f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_181 N_VPWR_c_255_n Y 0.0188775f $X=2.95 $Y=2.72 $X2=0 $Y2=0
cc_182 N_VPWR_c_249_n Y 0.01228f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_183 N_VPWR_c_249_n A_492_297# 0.00706335f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_184 N_Y_c_303_n N_VGND_c_332_n 0.0090392f $X=1.845 $Y=0.61 $X2=0 $Y2=0
cc_185 N_Y_M1005_s N_VGND_c_334_n 0.00414732f $X=1.56 $Y=0.235 $X2=0 $Y2=0
cc_186 N_Y_c_303_n N_VGND_c_334_n 0.0103575f $X=1.845 $Y=0.61 $X2=0 $Y2=0
cc_187 N_Y_c_303_n N_A_396_47#_c_376_n 0.0223649f $X=1.845 $Y=0.61 $X2=0 $Y2=0
cc_188 N_Y_c_293_n N_A_396_47#_c_374_n 0.00911194f $X=1.845 $Y=1.445 $X2=0 $Y2=0
cc_189 N_Y_c_303_n N_A_396_47#_c_374_n 0.00530028f $X=1.845 $Y=0.61 $X2=0 $Y2=0
cc_190 N_Y_c_295_n N_A_396_47#_c_374_n 0.00187199f $X=2.112 $Y=1.665 $X2=0 $Y2=0
cc_191 N_VGND_c_334_n A_122_47# 0.00412129f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_192 N_VGND_c_334_n N_A_396_47#_M1005_d 0.00714495f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_193 N_VGND_c_334_n N_A_396_47#_M1001_d 0.0025127f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_c_332_n N_A_396_47#_c_376_n 0.00714743f $X=2.52 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_c_334_n N_A_396_47#_c_376_n 0.00838703f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_M1009_d N_A_396_47#_c_373_n 0.00162089f $X=2.47 $Y=0.235 $X2=0
+ $Y2=0
cc_197 N_VGND_c_331_n N_A_396_47#_c_373_n 0.0122559f $X=2.605 $Y=0.39 $X2=0
+ $Y2=0
cc_198 N_VGND_c_332_n N_A_396_47#_c_373_n 0.00198695f $X=2.52 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_333_n N_A_396_47#_c_373_n 0.00198695f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_200 N_VGND_c_334_n N_A_396_47#_c_373_n 0.00835832f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_201 N_VGND_c_333_n N_A_396_47#_c_375_n 0.0216641f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_334_n N_A_396_47#_c_375_n 0.0141809f $X=3.45 $Y=0 $X2=0 $Y2=0
