# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o221a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o221a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 1.075000 3.325000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235000 1.075000 2.615000 1.705000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 1.075000 1.330000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 1.075000 1.905000 1.705000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.345000 1.325000 ;
    END
  END C1
  PIN VGND
    ANTENNADIFFAREA  0.546000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.970000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545000 0.265000 3.925000 0.735000 ;
        RECT 3.545000 0.735000 4.490000 0.905000 ;
        RECT 3.545000 1.875000 4.490000 2.045000 ;
        RECT 3.545000 2.045000 3.845000 2.465000 ;
        RECT 4.180000 0.905000 4.490000 1.875000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.170000  0.255000 0.500000 0.635000 ;
      RECT 0.170000  0.635000 0.765000 0.805000 ;
      RECT 0.250000  1.495000 1.350000 1.670000 ;
      RECT 0.250000  1.670000 0.580000 2.465000 ;
      RECT 0.545000  0.805000 0.765000 1.445000 ;
      RECT 0.545000  1.445000 1.350000 1.495000 ;
      RECT 0.670000  0.295000 2.005000 0.465000 ;
      RECT 0.800000  1.850000 1.010000 2.635000 ;
      RECT 1.135000  0.645000 1.570000 0.735000 ;
      RECT 1.135000  0.735000 2.985000 0.905000 ;
      RECT 1.180000  1.670000 1.350000 1.875000 ;
      RECT 1.180000  1.875000 2.965000 2.045000 ;
      RECT 1.700000  2.045000 2.455000 2.465000 ;
      RECT 2.265000  0.085000 2.435000 0.555000 ;
      RECT 2.605000  0.270000 2.985000 0.735000 ;
      RECT 2.795000  1.455000 3.715000 1.625000 ;
      RECT 2.795000  1.625000 2.965000 1.875000 ;
      RECT 3.145000  1.795000 3.375000 2.635000 ;
      RECT 3.205000  0.085000 3.375000 0.905000 ;
      RECT 3.495000  1.075000 3.875000 1.285000 ;
      RECT 3.495000  1.285000 3.715000 1.455000 ;
      RECT 4.015000  2.215000 4.405000 2.635000 ;
      RECT 4.145000  0.085000 4.315000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221a_2
END LIBRARY
