* NGSPICE file created from sky130_fd_sc_hdll__mux2i_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
M1000 Y A1 a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=1.215e+12p ps=1.043e+07u
M1001 VGND a_1311_21# a_109_47# VNB nshort w=650000u l=150000u
+  ad=1.03025e+12p pd=9.67e+06u as=9.3275e+11p ps=8.07e+06u
M1002 Y A0 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=1.16e+12p ps=1.032e+07u
M1003 VPWR a_1311_21# a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.475e+12p pd=1.295e+07u as=0p ps=0u
M1004 a_109_47# a_1311_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_117_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND S a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=8.645e+11p ps=7.86e+06u
M1007 a_493_297# A1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_485_47# S VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR S a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_109_47# A0 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=9.295e+11p ps=9.36e+06u
M1011 Y A1 a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A0 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A1 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_493_297# a_1311_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_117_297# A0 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND S a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_493_297# A1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_1311_21# a_493_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_485_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_117_297# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_109_47# a_1311_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A0 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_493_297# a_1311_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_485_47# S VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A0 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A1 a_485_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_485_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_1311_21# a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1311_21# S VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1030 a_117_297# A0 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR S a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_109_47# A0 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1311_21# S VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
.ends

