* File: sky130_fd_sc_hdll__a211o_1.pxi.spice
* Created: Thu Aug 27 18:51:24 2020
* 
x_PM_SKY130_FD_SC_HDLL__A211O_1%A_80_21# N_A_80_21#_M1006_d N_A_80_21#_M1009_d
+ N_A_80_21#_M1000_d N_A_80_21#_c_52_n N_A_80_21#_M1003_g N_A_80_21#_c_56_n
+ N_A_80_21#_M1002_g N_A_80_21#_c_53_n N_A_80_21#_c_64_p N_A_80_21#_c_124_p
+ N_A_80_21#_c_58_n N_A_80_21#_c_103_p N_A_80_21#_c_65_p N_A_80_21#_c_54_n
+ N_A_80_21#_c_59_n N_A_80_21#_c_89_p N_A_80_21#_c_78_p N_A_80_21#_c_55_n
+ PM_SKY130_FD_SC_HDLL__A211O_1%A_80_21#
x_PM_SKY130_FD_SC_HDLL__A211O_1%A2 N_A2_c_151_n N_A2_M1005_g N_A2_c_148_n
+ N_A2_M1007_g A2 A2 N_A2_c_150_n A2 PM_SKY130_FD_SC_HDLL__A211O_1%A2
x_PM_SKY130_FD_SC_HDLL__A211O_1%A1 N_A1_c_181_n N_A1_M1008_g N_A1_c_182_n
+ N_A1_M1006_g A1 A1 PM_SKY130_FD_SC_HDLL__A211O_1%A1
x_PM_SKY130_FD_SC_HDLL__A211O_1%B1 N_B1_c_211_n N_B1_M1001_g N_B1_c_212_n
+ N_B1_M1004_g B1 B1 PM_SKY130_FD_SC_HDLL__A211O_1%B1
x_PM_SKY130_FD_SC_HDLL__A211O_1%C1 N_C1_c_241_n N_C1_M1009_g N_C1_c_244_n
+ N_C1_M1000_g C1 N_C1_c_242_n C1 PM_SKY130_FD_SC_HDLL__A211O_1%C1
x_PM_SKY130_FD_SC_HDLL__A211O_1%X N_X_M1003_s N_X_M1002_s X X X X X X
+ N_X_c_268_n X PM_SKY130_FD_SC_HDLL__A211O_1%X
x_PM_SKY130_FD_SC_HDLL__A211O_1%VPWR N_VPWR_M1002_d N_VPWR_M1005_d
+ N_VPWR_c_285_n VPWR N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_284_n
+ N_VPWR_c_289_n N_VPWR_c_290_n N_VPWR_c_291_n VPWR
+ PM_SKY130_FD_SC_HDLL__A211O_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A211O_1%A_227_297# N_A_227_297#_M1005_s
+ N_A_227_297#_M1008_d N_A_227_297#_c_334_n N_A_227_297#_c_335_n
+ N_A_227_297#_c_339_n N_A_227_297#_c_340_n N_A_227_297#_c_342_n
+ PM_SKY130_FD_SC_HDLL__A211O_1%A_227_297#
x_PM_SKY130_FD_SC_HDLL__A211O_1%VGND N_VGND_M1003_d N_VGND_M1001_d VGND
+ N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n
+ N_VGND_c_369_n VGND PM_SKY130_FD_SC_HDLL__A211O_1%VGND
cc_1 VNB N_A_80_21#_c_52_n 0.0231018f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A_80_21#_c_53_n 0.00225869f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=1.16
cc_3 VNB N_A_80_21#_c_54_n 0.00773822f $X=-0.19 $Y=-0.24 $X2=3.31 $Y2=0.72
cc_4 VNB N_A_80_21#_c_55_n 0.0405625f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.202
cc_5 VNB N_A2_c_148_n 0.0222779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB A2 0.00583268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A2_c_150_n 0.0320015f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.985
cc_8 VNB N_A1_c_181_n 0.0236901f $X=-0.19 $Y=-0.24 $X2=2.26 $Y2=0.235
cc_9 VNB N_A1_c_182_n 0.0184721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB A1 0.00588498f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.985
cc_11 VNB N_B1_c_211_n 0.0175445f $X=-0.19 $Y=-0.24 $X2=2.26 $Y2=0.235
cc_12 VNB N_B1_c_212_n 0.023855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB B1 0.00198956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_C1_c_241_n 0.0230181f $X=-0.19 $Y=-0.24 $X2=2.26 $Y2=0.235
cc_15 VNB N_C1_c_242_n 0.0354259f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_16 VNB C1 0.0129734f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=1.505
cc_17 VNB N_X_c_268_n 0.0421698f $X=-0.19 $Y=-0.24 $X2=0.845 $Y2=0.72
cc_18 VNB N_VPWR_c_284_n 0.155873f $X=-0.19 $Y=-0.24 $X2=2.357 $Y2=0.53
cc_19 VNB N_VGND_c_364_n 0.033917f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_20 VNB N_VGND_c_365_n 0.0171009f $X=-0.19 $Y=-0.24 $X2=2.195 $Y2=0.72
cc_21 VNB N_VGND_c_366_n 0.201946f $X=-0.19 $Y=-0.24 $X2=0.845 $Y2=0.72
cc_22 VNB N_VGND_c_367_n 0.019692f $X=-0.19 $Y=-0.24 $X2=2.357 $Y2=0.625
cc_23 VNB N_VGND_c_368_n 0.0222886f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.85
cc_24 VNB N_VGND_c_369_n 0.00939383f $X=-0.19 $Y=-0.24 $X2=3.422 $Y2=0.53
cc_25 VPB N_A_80_21#_c_56_n 0.0214006f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_26 VPB N_A_80_21#_c_53_n 0.00319497f $X=-0.19 $Y=1.305 $X2=0.735 $Y2=1.16
cc_27 VPB N_A_80_21#_c_58_n 0.0228096f $X=-0.19 $Y=1.305 $X2=3.205 $Y2=1.595
cc_28 VPB N_A_80_21#_c_59_n 0.0290872f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.85
cc_29 VPB N_A_80_21#_c_55_n 0.0162194f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.202
cc_30 VPB N_A2_c_151_n 0.0207525f $X=-0.19 $Y=1.305 $X2=2.26 $Y2=0.235
cc_31 VPB A2 0.00222587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A2_c_150_n 0.0151258f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_33 VPB N_A1_c_181_n 0.0280466f $X=-0.19 $Y=1.305 $X2=2.26 $Y2=0.235
cc_34 VPB A1 0.00218477f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_35 VPB N_B1_c_212_n 0.0270517f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB B1 0.00198956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_C1_c_244_n 0.0217197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_C1_c_242_n 0.0165117f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_39 VPB C1 0.00223262f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.505
cc_40 VPB X 0.0294769f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_41 VPB N_X_c_268_n 0.00882641f $X=-0.19 $Y=1.305 $X2=0.845 $Y2=0.72
cc_42 VPB X 0.0065071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_285_n 0.00790262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_286_n 0.0153767f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_45 VPB N_VPWR_c_287_n 0.0453429f $X=-0.19 $Y=1.305 $X2=2.357 $Y2=0.625
cc_46 VPB N_VPWR_c_284_n 0.0537992f $X=-0.19 $Y=1.305 $X2=2.357 $Y2=0.53
cc_47 VPB N_VPWR_c_289_n 0.00583344f $X=-0.19 $Y=1.305 $X2=3.31 $Y2=0.72
cc_48 VPB N_VPWR_c_290_n 0.0154544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_291_n 0.00923591f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.202
cc_50 VPB N_A_227_297#_c_334_n 0.00283489f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_227_297#_c_335_n 0.0034964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 N_A_80_21#_c_53_n N_A2_c_151_n 0.00226662f $X=0.735 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_53 N_A_80_21#_c_58_n N_A2_c_151_n 0.0154778f $X=3.205 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_54 N_A_80_21#_c_53_n N_A2_c_148_n 0.00406595f $X=0.735 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_80_21#_c_64_p N_A2_c_148_n 0.0160373f $X=2.195 $Y=0.72 $X2=0 $Y2=0
cc_56 N_A_80_21#_c_65_p N_A2_c_148_n 0.00166353f $X=2.405 $Y=0.53 $X2=0 $Y2=0
cc_57 N_A_80_21#_c_53_n A2 0.0270712f $X=0.735 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_80_21#_c_64_p A2 0.0449055f $X=2.195 $Y=0.72 $X2=0 $Y2=0
cc_59 N_A_80_21#_c_58_n A2 0.0448371f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_60 N_A_80_21#_c_55_n A2 0.00243729f $X=0.5 $Y=1.202 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_53_n N_A2_c_150_n 0.00241891f $X=0.735 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_64_p N_A2_c_150_n 0.00718142f $X=2.195 $Y=0.72 $X2=0 $Y2=0
cc_63 N_A_80_21#_c_58_n N_A2_c_150_n 0.00591483f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_55_n N_A2_c_150_n 0.0160667f $X=0.5 $Y=1.202 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_64_p N_A1_c_181_n 0.0038311f $X=2.195 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_66 N_A_80_21#_c_58_n N_A1_c_181_n 0.0159428f $X=3.205 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_67 N_A_80_21#_c_64_p N_A1_c_182_n 0.00791421f $X=2.195 $Y=0.72 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_65_p N_A1_c_182_n 0.0100957f $X=2.405 $Y=0.53 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_78_p N_A1_c_182_n 0.00315047f $X=2.357 $Y=0.72 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_64_p A1 0.0215584f $X=2.195 $Y=0.72 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_58_n A1 0.0336551f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_78_p A1 0.0131342f $X=2.357 $Y=0.72 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_54_n N_B1_c_211_n 0.0134653f $X=3.31 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_74 N_A_80_21#_c_58_n N_B1_c_212_n 0.0215941f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_54_n N_B1_c_212_n 0.0038311f $X=3.31 $Y=0.72 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_59_n N_B1_c_212_n 0.00275944f $X=3.41 $Y=1.85 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_58_n B1 0.0311114f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_54_n B1 0.0311261f $X=3.31 $Y=0.72 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_54_n N_C1_c_241_n 0.0168396f $X=3.31 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_80_21#_c_89_p N_C1_c_241_n 0.00538893f $X=3.41 $Y=0.53 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_80_21#_c_58_n N_C1_c_244_n 0.022253f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_59_n N_C1_c_244_n 0.0184497f $X=3.41 $Y=1.85 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_58_n N_C1_c_242_n 0.00611079f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_54_n N_C1_c_242_n 0.00764341f $X=3.31 $Y=0.72 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_58_n C1 0.0184833f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_54_n C1 0.0177994f $X=3.31 $Y=0.72 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_52_n N_X_c_268_n 0.0161551f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_56_n N_X_c_268_n 0.00265688f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_53_n N_X_c_268_n 0.0461845f $X=0.735 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_55_n N_X_c_268_n 0.0151531f $X=0.5 $Y=1.202 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_56_n X 0.00249812f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_53_n N_VPWR_M1002_d 3.22661e-19 $X=0.735 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_80_21#_c_58_n N_VPWR_M1002_d 6.41771e-19 $X=3.205 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_80_21#_c_103_p N_VPWR_M1002_d 0.00446661f $X=0.845 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_80_21#_c_58_n N_VPWR_M1005_d 0.0136877f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_56_n N_VPWR_c_285_n 0.0192899f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_58_n N_VPWR_c_285_n 0.00395007f $X=3.205 $Y=1.595 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_103_p N_VPWR_c_285_n 0.0142107f $X=0.845 $Y=1.595 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_55_n N_VPWR_c_285_n 9.00282e-19 $X=0.5 $Y=1.202 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_56_n N_VPWR_c_286_n 0.00447018f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_59_n N_VPWR_c_287_n 0.0203764f $X=3.41 $Y=1.85 $X2=0 $Y2=0
cc_102 N_A_80_21#_M1000_d N_VPWR_c_284_n 0.00222762f $X=3.26 $Y=1.485 $X2=0
+ $Y2=0
cc_103 N_A_80_21#_c_56_n N_VPWR_c_284_n 0.00855297f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_59_n N_VPWR_c_284_n 0.0127069f $X=3.41 $Y=1.85 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_58_n N_A_227_297#_M1005_s 0.00518781f $X=3.205 $Y=1.595
+ $X2=-0.19 $Y2=-0.24
cc_106 N_A_80_21#_c_58_n N_A_227_297#_M1008_d 0.00689361f $X=3.205 $Y=1.595
+ $X2=0 $Y2=0
cc_107 N_A_80_21#_c_58_n N_A_227_297#_c_334_n 0.0200841f $X=3.205 $Y=1.595 $X2=0
+ $Y2=0
cc_108 N_A_80_21#_c_58_n N_A_227_297#_c_339_n 0.050075f $X=3.205 $Y=1.595 $X2=0
+ $Y2=0
cc_109 N_A_80_21#_c_58_n N_A_227_297#_c_340_n 0.0154327f $X=3.205 $Y=1.595 $X2=0
+ $Y2=0
cc_110 N_A_80_21#_c_59_n N_A_227_297#_c_340_n 0.00608274f $X=3.41 $Y=1.85 $X2=0
+ $Y2=0
cc_111 N_A_80_21#_c_59_n N_A_227_297#_c_342_n 0.00880832f $X=3.41 $Y=1.85 $X2=0
+ $Y2=0
cc_112 N_A_80_21#_c_58_n A_546_297# 0.0114769f $X=3.205 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_113 N_A_80_21#_c_53_n N_VGND_M1003_d 0.001211f $X=0.735 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A_80_21#_c_64_p N_VGND_M1003_d 0.0194434f $X=2.195 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_115 N_A_80_21#_c_124_p N_VGND_M1003_d 0.00539361f $X=0.845 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_116 N_A_80_21#_c_54_n N_VGND_M1001_d 0.0055812f $X=3.31 $Y=0.72 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_64_p N_VGND_c_364_n 0.0127336f $X=2.195 $Y=0.72 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_65_p N_VGND_c_364_n 0.0179497f $X=2.405 $Y=0.53 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_54_n N_VGND_c_364_n 0.0028245f $X=3.31 $Y=0.72 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_54_n N_VGND_c_365_n 0.00351404f $X=3.31 $Y=0.72 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_89_p N_VGND_c_365_n 0.0145106f $X=3.41 $Y=0.53 $X2=0 $Y2=0
cc_122 N_A_80_21#_M1006_d N_VGND_c_366_n 0.00231366f $X=2.26 $Y=0.235 $X2=0
+ $Y2=0
cc_123 N_A_80_21#_M1009_d N_VGND_c_366_n 0.00285424f $X=3.22 $Y=0.235 $X2=0
+ $Y2=0
cc_124 N_A_80_21#_c_52_n N_VGND_c_366_n 0.0122215f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_64_p N_VGND_c_366_n 0.0241299f $X=2.195 $Y=0.72 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_124_p N_VGND_c_366_n 0.00247904f $X=0.845 $Y=0.72 $X2=0
+ $Y2=0
cc_127 N_A_80_21#_c_65_p N_VGND_c_366_n 0.0120156f $X=2.405 $Y=0.53 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_54_n N_VGND_c_366_n 0.0120267f $X=3.31 $Y=0.72 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_89_p N_VGND_c_366_n 0.00849891f $X=3.41 $Y=0.53 $X2=0 $Y2=0
cc_130 N_A_80_21#_c_52_n N_VGND_c_367_n 0.00549284f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_131 N_A_80_21#_c_124_p N_VGND_c_367_n 9.58021e-19 $X=0.845 $Y=0.72 $X2=0
+ $Y2=0
cc_132 N_A_80_21#_c_52_n N_VGND_c_368_n 0.00991501f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_80_21#_c_64_p N_VGND_c_368_n 0.0417213f $X=2.195 $Y=0.72 $X2=0 $Y2=0
cc_134 N_A_80_21#_c_124_p N_VGND_c_368_n 0.0158738f $X=0.845 $Y=0.72 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_55_n N_VGND_c_368_n 7.26772e-19 $X=0.5 $Y=1.202 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_54_n N_VGND_c_369_n 0.0209815f $X=3.31 $Y=0.72 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_89_p N_VGND_c_369_n 0.0114768f $X=3.41 $Y=0.53 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_64_p A_320_47# 0.0171987f $X=2.195 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_139 N_A2_c_151_n N_A1_c_181_n 0.0260897f $X=1.5 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_140 A2 N_A1_c_181_n 0.00112958f $X=1.465 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_141 N_A2_c_150_n N_A1_c_181_n 0.0145321f $X=1.5 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_142 N_A2_c_148_n N_A1_c_182_n 0.0216402f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_143 A2 A1 0.0301398f $X=1.465 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A2_c_150_n A1 0.00103003f $X=1.5 $Y=1.202 $X2=0 $Y2=0
cc_145 N_A2_c_151_n N_VPWR_c_285_n 0.00202168f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_151_n N_VPWR_c_284_n 0.0051021f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A2_c_151_n N_VPWR_c_290_n 0.00324069f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A2_c_151_n N_VPWR_c_291_n 0.0100641f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A2_c_151_n N_A_227_297#_c_339_n 0.0137899f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A2_c_148_n N_VGND_c_364_n 0.0042361f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A2_c_148_n N_VGND_c_366_n 0.00763232f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A2_c_148_n N_VGND_c_368_n 0.00904025f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A1_c_182_n N_B1_c_211_n 0.0212715f $X=2.185 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A1_c_181_n N_B1_c_212_n 0.0428624f $X=2.16 $Y=1.41 $X2=0 $Y2=0
cc_155 A1 N_B1_c_212_n 0.00247635f $X=2.105 $Y=1.19 $X2=0 $Y2=0
cc_156 N_A1_c_181_n B1 3.12382e-19 $X=2.16 $Y=1.41 $X2=0 $Y2=0
cc_157 A1 B1 0.0247209f $X=2.105 $Y=1.19 $X2=0 $Y2=0
cc_158 N_A1_c_181_n N_VPWR_c_287_n 0.00465273f $X=2.16 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A1_c_181_n N_VPWR_c_284_n 0.00528712f $X=2.16 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A1_c_181_n N_VPWR_c_291_n 0.0120416f $X=2.16 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A1_c_181_n N_A_227_297#_c_339_n 0.0142343f $X=2.16 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A1_c_182_n N_VGND_c_364_n 0.00397444f $X=2.185 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_c_182_n N_VGND_c_366_n 0.00617099f $X=2.185 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B1_c_211_n N_C1_c_241_n 0.0228548f $X=2.615 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_165 N_B1_c_212_n N_C1_c_244_n 0.042218f $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B1_c_212_n N_C1_c_242_n 0.0253584f $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_167 B1 N_C1_c_242_n 0.00874817f $X=2.855 $Y=1.105 $X2=0 $Y2=0
cc_168 N_B1_c_212_n C1 2.11477e-19 $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_169 B1 C1 0.0198324f $X=2.855 $Y=1.105 $X2=0 $Y2=0
cc_170 N_B1_c_212_n N_VPWR_c_287_n 0.00681403f $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_171 N_B1_c_212_n N_VPWR_c_284_n 0.0124207f $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B1_c_212_n N_VPWR_c_291_n 0.00103643f $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_173 N_B1_c_212_n N_A_227_297#_c_340_n 0.00471889f $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B1_c_212_n N_A_227_297#_c_342_n 0.00716211f $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B1_c_211_n N_VGND_c_364_n 0.0042361f $X=2.615 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B1_c_211_n N_VGND_c_366_n 0.00596762f $X=2.615 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B1_c_211_n N_VGND_c_369_n 0.00464734f $X=2.615 $Y=0.995 $X2=0 $Y2=0
cc_178 N_C1_c_244_n N_VPWR_c_287_n 0.00621235f $X=3.17 $Y=1.41 $X2=0 $Y2=0
cc_179 N_C1_c_244_n N_VPWR_c_284_n 0.0118946f $X=3.17 $Y=1.41 $X2=0 $Y2=0
cc_180 N_C1_c_244_n N_A_227_297#_c_340_n 6.83796e-19 $X=3.17 $Y=1.41 $X2=0 $Y2=0
cc_181 N_C1_c_244_n N_A_227_297#_c_342_n 0.00107437f $X=3.17 $Y=1.41 $X2=0 $Y2=0
cc_182 N_C1_c_241_n N_VGND_c_365_n 0.0039537f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_183 N_C1_c_241_n N_VGND_c_366_n 0.00558493f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_184 N_C1_c_241_n N_VGND_c_369_n 0.00785612f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_185 X N_VPWR_c_286_n 0.017406f $X=0.135 $Y=1.785 $X2=0 $Y2=0
cc_186 N_X_M1002_s N_VPWR_c_284_n 0.00412825f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_187 X N_VPWR_c_284_n 0.0100753f $X=0.135 $Y=1.785 $X2=0 $Y2=0
cc_188 N_X_M1003_s N_VGND_c_366_n 0.00213747f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_189 N_X_c_268_n N_VGND_c_366_n 0.0125813f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_190 N_X_c_268_n N_VGND_c_367_n 0.0201263f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_191 N_X_c_268_n N_VGND_c_368_n 0.0123783f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_192 N_VPWR_c_284_n N_A_227_297#_M1005_s 0.0024001f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_193 N_VPWR_c_284_n N_A_227_297#_M1008_d 0.00257715f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_285_n N_A_227_297#_c_334_n 0.0148677f $X=0.74 $Y=2 $X2=0 $Y2=0
cc_195 N_VPWR_c_285_n N_A_227_297#_c_335_n 0.0274913f $X=0.74 $Y=2 $X2=0 $Y2=0
cc_196 N_VPWR_c_284_n N_A_227_297#_c_335_n 0.00984593f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_290_n N_A_227_297#_c_335_n 0.0168929f $X=1.525 $Y=2.535 $X2=0
+ $Y2=0
cc_198 N_VPWR_M1005_d N_A_227_297#_c_339_n 0.00924429f $X=1.59 $Y=1.485 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_287_n N_A_227_297#_c_339_n 0.00335192f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_284_n N_A_227_297#_c_339_n 0.0123194f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_290_n N_A_227_297#_c_339_n 0.00249844f $X=1.525 $Y=2.535 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_291_n N_A_227_297#_c_339_n 0.0339748f $X=2.085 $Y=2.535 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_287_n N_A_227_297#_c_342_n 0.0149642f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_284_n N_A_227_297#_c_342_n 0.00970974f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_284_n A_546_297# 0.014961f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_206 N_VGND_c_366_n A_320_47# 0.00590778f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
