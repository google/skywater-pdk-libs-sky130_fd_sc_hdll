* File: sky130_fd_sc_hdll__muxb8to1_4.spice
* Created: Wed Sep  2 08:36:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__muxb8to1_4.pex.spice"
.subckt sky130_fd_sc_hdll__muxb8to1_4  VNB VPB S[0] S[1] D[0] D[1] D[2] D[3]
+ S[2] S[3] S[4] S[5] D[4] D[5] D[6] D[7] S[6] S[7] VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* S[7]	S[7]
* S[6]	S[6]
* D[7]	D[7]
* D[6]	D[6]
* D[5]	D[5]
* D[4]	D[4]
* S[5]	S[5]
* S[4]	S[4]
* S[3]	S[3]
* S[2]	S[2]
* D[3]	D[3]
* D[2]	D[2]
* D[1]	D[1]
* D[0]	D[0]
* S[1]	S[1]
* S[0]	S[0]
* VPB	VPB
* VNB	VNB
MM1043 N_VGND_M1043_d N_S[0]_M1043_g N_A_142_325#_M1043_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1084 N_A_142_599#_M1084_d N_S[1]_M1084_g N_VGND_M1084_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1067 N_VGND_M1067_d N_S[0]_M1067_g N_A_142_325#_M1043_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1138 N_A_142_599#_M1084_d N_S[1]_M1138_g N_VGND_M1138_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_405_66#_M1003_d N_S[0]_M1003_g N_Z_M1003_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1029 N_A_405_918#_M1029_d N_S[1]_M1029_g N_Z_M1029_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1100 N_A_405_66#_M1100_d N_S[0]_M1100_g N_Z_M1003_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1058 N_A_405_918#_M1058_d N_S[1]_M1058_g N_Z_M1029_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1109 N_A_405_66#_M1100_d N_S[0]_M1109_g N_Z_M1109_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1083 N_A_405_918#_M1058_d N_S[1]_M1083_g N_Z_M1083_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1133 N_A_405_66#_M1133_d N_S[0]_M1133_g N_Z_M1109_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1102 N_A_405_918#_M1102_d N_S[1]_M1102_g N_Z_M1083_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1065 N_A_405_66#_M1065_d N_D[0]_M1065_g N_VGND_M1065_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1030 N_A_405_918#_M1030_d N_D[1]_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1097 N_A_405_66#_M1065_d N_D[0]_M1097_g N_VGND_M1097_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.6 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1059 N_A_405_918#_M1030_d N_D[1]_M1059_g N_VGND_M1059_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.6 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1151 N_A_405_66#_M1151_d N_D[0]_M1151_g N_VGND_M1097_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.1 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1068 N_A_405_918#_M1068_d N_D[1]_M1068_g N_VGND_M1059_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.1 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1156 N_A_405_66#_M1151_d N_D[0]_M1156_g N_VGND_M1156_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.13975 PD=0.92 PS=1.08 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75001.5 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1157 N_A_405_918#_M1068_d N_D[1]_M1157_g N_VGND_M1157_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.13975 PD=0.92 PS=1.08 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75001.5 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1156_s N_D[2]_M1013_g N_A_1315_47#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.13975 AS=0.08775 PD=1.08 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75002.1 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1015 N_A_1315_911#_M1015_d N_D[3]_M1015_g N_VGND_M1157_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.13975 PD=0.92 PS=1.08 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75002.1 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1037 N_VGND_M1037_d N_D[2]_M1037_g N_A_1315_47#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.5 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1047 N_A_1315_911#_M1015_d N_D[3]_M1047_g N_VGND_M1047_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.5 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1069 N_VGND_M1037_d N_D[2]_M1069_g N_A_1315_47#_M1069_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1104 N_A_1315_911#_M1104_d N_D[3]_M1104_g N_VGND_M1047_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1150 N_VGND_M1150_d N_D[2]_M1150_g N_A_1315_47#_M1069_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1136 N_A_1315_911#_M1104_d N_D[3]_M1136_g N_VGND_M1136_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1024 N_Z_M1024_d N_S[2]_M1024_g N_A_1315_47#_M1024_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1016 N_Z_M1016_d N_S[3]_M1016_g N_A_1315_911#_M1016_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1028 N_Z_M1024_d N_S[2]_M1028_g N_A_1315_47#_M1028_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1020 N_Z_M1016_d N_S[3]_M1020_g N_A_1315_911#_M1020_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1044 N_Z_M1044_d N_S[2]_M1044_g N_A_1315_47#_M1028_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1048 N_Z_M1048_d N_S[3]_M1048_g N_A_1315_911#_M1020_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1057 N_Z_M1044_d N_S[2]_M1057_g N_A_1315_47#_M1057_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1135 N_Z_M1048_d N_S[3]_M1135_g N_A_1315_911#_M1135_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1094 N_VGND_M1094_d N_S[2]_M1094_g N_A_1755_265#_M1094_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1060 N_VGND_M1060_d N_S[3]_M1060_g N_A_1755_793#_M1060_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1103 N_VGND_M1103_d N_S[2]_M1103_g N_A_1755_265#_M1094_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1140 N_VGND_M1140_d N_S[3]_M1140_g N_A_1755_793#_M1060_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1121 N_VGND_M1121_d N_S[4]_M1121_g N_A_2626_325#_M1121_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1074 N_VGND_M1074_d N_S[5]_M1074_g N_A_2626_599#_M1074_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1129 N_VGND_M1129_d N_S[4]_M1129_g N_A_2626_325#_M1121_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1154 N_VGND_M1154_d N_S[5]_M1154_g N_A_2626_599#_M1074_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_2889_66#_M1006_d N_S[4]_M1006_g N_Z_M1006_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1009 N_Z_M1009_d N_S[5]_M1009_g N_A_2889_918#_M1009_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1022 N_A_2889_66#_M1022_d N_S[4]_M1022_g N_Z_M1006_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1038 N_Z_M1009_d N_S[5]_M1038_g N_A_2889_918#_M1038_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1035 N_A_2889_66#_M1022_d N_S[4]_M1035_g N_Z_M1035_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1112 N_Z_M1112_d N_S[5]_M1112_g N_A_2889_918#_M1038_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1066 N_A_2889_66#_M1066_d N_S[4]_M1066_g N_Z_M1035_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1142 N_Z_M1112_d N_S[5]_M1142_g N_A_2889_918#_M1142_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1027 N_VGND_M1027_d N_D[4]_M1027_g N_A_2889_66#_M1027_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1033 N_VGND_M1033_d N_D[5]_M1033_g N_A_2889_918#_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1034 N_VGND_M1034_d N_D[4]_M1034_g N_A_2889_66#_M1027_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1077 N_VGND_M1077_d N_D[5]_M1077_g N_A_2889_918#_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1045 N_VGND_M1034_d N_D[4]_M1045_g N_A_2889_66#_M1045_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1106 N_VGND_M1077_d N_D[5]_M1106_g N_A_2889_918#_M1106_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1079 N_VGND_M1079_d N_D[4]_M1079_g N_A_2889_66#_M1045_s VNB NSHORT L=0.15
+ W=0.65 AD=0.13975 AS=0.08775 PD=1.08 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1107 N_VGND_M1107_d N_D[5]_M1107_g N_A_2889_918#_M1106_s VNB NSHORT L=0.15
+ W=0.65 AD=0.13975 AS=0.08775 PD=1.08 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1005 N_A_3799_47#_M1005_d N_D[6]_M1005_g N_VGND_M1079_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.13975 PD=0.92 PS=1.08 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75002.1 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1107_d N_D[7]_M1014_g N_A_3799_911#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.13975 AS=0.08775 PD=1.08 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75002.1 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1081 N_A_3799_47#_M1005_d N_D[6]_M1081_g N_VGND_M1081_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.5 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1025_d N_D[7]_M1025_g N_A_3799_911#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.5 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1111 N_A_3799_47#_M1111_d N_D[6]_M1111_g N_VGND_M1081_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1026 N_VGND_M1025_d N_D[7]_M1026_g N_A_3799_911#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1159 N_A_3799_47#_M1111_d N_D[6]_M1159_g N_VGND_M1159_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1098 N_VGND_M1098_d N_D[7]_M1098_g N_A_3799_911#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1089 N_A_3799_47#_M1089_d N_S[6]_M1089_g N_Z_M1089_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1008 N_Z_M1008_d N_S[7]_M1008_g N_A_3799_911#_M1008_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1101 N_A_3799_47#_M1101_d N_S[6]_M1101_g N_Z_M1089_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1063 N_Z_M1008_d N_S[7]_M1063_g N_A_3799_911#_M1063_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1122 N_A_3799_47#_M1101_d N_S[6]_M1122_g N_Z_M1122_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1091 N_Z_M1091_d N_S[7]_M1091_g N_A_3799_911#_M1063_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1132 N_A_3799_47#_M1132_d N_S[6]_M1132_g N_Z_M1122_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1144 N_Z_M1091_d N_S[7]_M1144_g N_A_3799_911#_M1144_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1032 N_A_4239_265#_M1032_d N_S[6]_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1114 N_A_4239_793#_M1114_d N_S[7]_M1114_g N_VGND_M1114_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1061 N_A_4239_265#_M1032_d N_S[6]_M1061_g N_VGND_M1061_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1149 N_A_4239_793#_M1114_d N_S[7]_M1149_g N_VGND_M1149_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_S[0]_M1001_g N_A_142_325#_M1001_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1052 N_VPWR_M1052_d N_S[1]_M1052_g N_A_142_599#_M1052_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1040 N_VPWR_M1040_d N_S[0]_M1040_g N_A_142_325#_M1001_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1088 N_VPWR_M1088_d N_S[1]_M1088_g N_A_142_599#_M1052_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1010 N_A_355_311#_M1010_d N_A_142_325#_M1010_g N_Z_M1010_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1054 N_A_355_613#_M1054_d N_A_142_599#_M1054_g N_Z_M1054_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1019 N_A_355_311#_M1019_d N_A_142_325#_M1019_g N_Z_M1010_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1080 N_A_355_613#_M1080_d N_A_142_599#_M1080_g N_Z_M1054_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1051 N_A_355_311#_M1019_d N_A_142_325#_M1051_g N_Z_M1051_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1092 N_A_355_613#_M1080_d N_A_142_599#_M1092_g N_Z_M1092_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1147 N_A_355_311#_M1147_d N_A_142_325#_M1147_g N_Z_M1051_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1123 N_A_355_613#_M1123_d N_A_142_599#_M1123_g N_Z_M1092_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1012 N_A_355_311#_M1012_d N_D[0]_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1017 N_A_355_613#_M1017_d N_D[1]_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1049 N_A_355_311#_M1012_d N_D[0]_M1049_g N_VPWR_M1049_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1055 N_A_355_613#_M1017_d N_D[1]_M1055_g N_VPWR_M1055_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1086 N_A_355_311#_M1086_d N_D[0]_M1086_g N_VPWR_M1049_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1093 N_A_355_613#_M1093_d N_D[1]_M1093_g N_VPWR_M1055_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1137 N_A_355_311#_M1086_d N_D[0]_M1137_g N_VPWR_M1137_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.175 PD=1.29 PS=1.35 NRD=0.9653 NRS=6.8753 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1141 N_A_355_613#_M1093_d N_D[1]_M1141_g N_VPWR_M1141_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.175 PD=1.29 PS=1.35 NRD=0.9653 NRS=6.8753 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1071 N_VPWR_M1137_s N_D[2]_M1071_g N_A_1313_297#_M1071_s VPB PHIGHVT L=0.18
+ W=1 AD=0.175 AS=0.145 PD=1.35 PS=1.29 NRD=6.8753 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1000 N_A_1313_591#_M1000_d N_D[3]_M1000_g N_VPWR_M1141_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.175 PD=1.29 PS=1.35 NRD=0.9653 NRS=6.8753 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1090 N_VPWR_M1090_d N_D[2]_M1090_g N_A_1313_297#_M1071_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1076 N_A_1313_591#_M1000_d N_D[3]_M1076_g N_VPWR_M1076_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1118 N_VPWR_M1090_d N_D[2]_M1118_g N_A_1313_297#_M1118_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1095 N_A_1313_591#_M1095_d N_D[3]_M1095_g N_VPWR_M1076_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1158 N_VPWR_M1158_d N_D[2]_M1158_g N_A_1313_297#_M1118_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1120 N_A_1313_591#_M1095_d N_D[3]_M1120_g N_VPWR_M1120_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1050 N_Z_M1050_d N_A_1755_265#_M1050_g N_A_1313_297#_M1050_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1031 N_Z_M1031_d N_A_1755_793#_M1031_g N_A_1313_591#_M1031_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1073 N_Z_M1050_d N_A_1755_265#_M1073_g N_A_1313_297#_M1073_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1036 N_Z_M1031_d N_A_1755_793#_M1036_g N_A_1313_591#_M1036_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1116 N_Z_M1116_d N_A_1755_265#_M1116_g N_A_1313_297#_M1073_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1124 N_Z_M1124_d N_A_1755_793#_M1124_g N_A_1313_591#_M1036_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1126 N_Z_M1116_d N_A_1755_265#_M1126_g N_A_1313_297#_M1126_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1152 N_Z_M1124_d N_A_1755_793#_M1152_g N_A_1313_591#_M1152_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1072 N_VPWR_M1072_d N_S[2]_M1072_g N_A_1755_265#_M1072_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1007 N_A_1755_793#_M1007_d N_S[3]_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1115 N_VPWR_M1115_d N_S[2]_M1115_g N_A_1755_265#_M1072_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1125 N_A_1755_793#_M1007_d N_S[3]_M1125_g N_VPWR_M1125_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1128 N_VPWR_M1128_d N_S[4]_M1128_g N_A_2626_325#_M1128_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1018 N_VPWR_M1018_d N_S[5]_M1018_g N_A_2626_599#_M1018_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1155 N_VPWR_M1155_d N_S[4]_M1155_g N_A_2626_325#_M1128_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1039 N_VPWR_M1039_d N_S[5]_M1039_g N_A_2626_599#_M1018_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1004 N_Z_M1004_d N_A_2626_325#_M1004_g N_A_2839_311#_M1004_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1021 N_A_2839_613#_M1021_d N_A_2626_599#_M1021_g N_Z_M1021_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1110 N_Z_M1004_d N_A_2626_325#_M1110_g N_A_2839_311#_M1110_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1041 N_A_2839_613#_M1041_d N_A_2626_599#_M1041_g N_Z_M1021_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1131 N_Z_M1131_d N_A_2626_325#_M1131_g N_A_2839_311#_M1110_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1056 N_A_2839_613#_M1041_d N_A_2626_599#_M1056_g N_Z_M1056_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1146 N_Z_M1131_d N_A_2626_325#_M1146_g N_A_2839_311#_M1146_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1078 N_A_2839_613#_M1078_d N_A_2626_599#_M1078_g N_Z_M1056_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1042 N_VPWR_M1042_d N_D[4]_M1042_g N_A_2839_311#_M1042_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1046 N_VPWR_M1046_d N_D[5]_M1046_g N_A_2839_613#_M1046_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1062 N_VPWR_M1062_d N_D[4]_M1062_g N_A_2839_311#_M1042_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1070 N_VPWR_M1070_d N_D[5]_M1070_g N_A_2839_613#_M1046_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1105 N_VPWR_M1062_d N_D[4]_M1105_g N_A_2839_311#_M1105_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1113 N_VPWR_M1070_d N_D[5]_M1113_g N_A_2839_613#_M1113_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1127 N_VPWR_M1127_d N_D[4]_M1127_g N_A_2839_311#_M1105_s VPB PHIGHVT L=0.18
+ W=1 AD=0.175 AS=0.145 PD=1.35 PS=1.29 NRD=6.8753 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1134 N_VPWR_M1134_d N_D[5]_M1134_g N_A_2839_613#_M1113_s VPB PHIGHVT L=0.18
+ W=1 AD=0.175 AS=0.145 PD=1.35 PS=1.29 NRD=6.8753 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1082 N_A_3797_297#_M1082_d N_D[6]_M1082_g N_VPWR_M1127_d VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.175 PD=1.29 PS=1.35 NRD=0.9653 NRS=6.8753 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1087 N_A_3797_591#_M1087_d N_D[7]_M1087_g N_VPWR_M1134_d VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.175 PD=1.29 PS=1.35 NRD=0.9653 NRS=6.8753 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1108 N_A_3797_297#_M1082_d N_D[6]_M1108_g N_VPWR_M1108_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1117 N_A_3797_591#_M1087_d N_D[7]_M1117_g N_VPWR_M1117_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1130 N_A_3797_297#_M1130_d N_D[6]_M1130_g N_VPWR_M1108_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1139 N_A_3797_591#_M1139_d N_D[7]_M1139_g N_VPWR_M1117_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1145 N_A_3797_297#_M1130_d N_D[6]_M1145_g N_VPWR_M1145_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1153 N_A_3797_591#_M1139_d N_D[7]_M1153_g N_VPWR_M1153_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1002 N_A_3797_297#_M1002_d N_A_4239_265#_M1002_g N_Z_M1002_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1011 N_A_3797_591#_M1011_d N_A_4239_793#_M1011_g N_Z_M1011_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1023 N_A_3797_297#_M1023_d N_A_4239_265#_M1023_g N_Z_M1002_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1053 N_A_3797_591#_M1053_d N_A_4239_793#_M1053_g N_Z_M1011_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1099 N_A_3797_297#_M1023_d N_A_4239_265#_M1099_g N_Z_M1099_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1075 N_A_3797_591#_M1053_d N_A_4239_793#_M1075_g N_Z_M1075_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1143 N_A_3797_297#_M1143_d N_A_4239_265#_M1143_g N_Z_M1099_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1096 N_A_3797_591#_M1096_d N_A_4239_793#_M1096_g N_Z_M1075_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1064 N_VPWR_M1064_d N_S[6]_M1064_g N_A_4239_265#_M1064_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1119 N_VPWR_M1119_d N_S[7]_M1119_g N_A_4239_793#_M1119_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1085 N_VPWR_M1085_d N_S[6]_M1085_g N_A_4239_265#_M1064_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1148 N_VPWR_M1148_d N_S[7]_M1148_g N_A_4239_793#_M1119_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
DX160_noxref VNB VPB NWDIODE A=71.3726 P=56.1
c_903 VPB 0 9.66518e-19 $X=18.545 $Y=2.635
*
.include "sky130_fd_sc_hdll__muxb8to1_4.pxi.spice"
*
.ends
*
*
