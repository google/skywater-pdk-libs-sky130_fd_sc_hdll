* File: sky130_fd_sc_hdll__dfstp_4.pxi.spice
* Created: Wed Sep  2 08:28:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%CLK N_CLK_c_239_n N_CLK_c_240_n N_CLK_M1007_g
+ N_CLK_c_234_n N_CLK_M1025_g N_CLK_c_235_n CLK CLK N_CLK_c_237_n N_CLK_c_238_n
+ PM_SKY130_FD_SC_HDLL__DFSTP_4%CLK
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%A_27_47# N_A_27_47#_M1025_s N_A_27_47#_M1007_s
+ N_A_27_47#_c_289_n N_A_27_47#_c_290_n N_A_27_47#_M1032_g N_A_27_47#_M1002_g
+ N_A_27_47#_c_276_n N_A_27_47#_M1003_g N_A_27_47#_c_291_n N_A_27_47#_M1024_g
+ N_A_27_47#_c_292_n N_A_27_47#_M1035_g N_A_27_47#_c_277_n N_A_27_47#_M1005_g
+ N_A_27_47#_c_517_p N_A_27_47#_c_278_n N_A_27_47#_c_279_n N_A_27_47#_c_293_n
+ N_A_27_47#_c_402_p N_A_27_47#_c_280_n N_A_27_47#_c_281_n N_A_27_47#_c_282_n
+ N_A_27_47#_c_283_n N_A_27_47#_c_284_n N_A_27_47#_c_285_n N_A_27_47#_c_297_n
+ N_A_27_47#_c_286_n N_A_27_47#_c_298_n N_A_27_47#_c_299_n N_A_27_47#_c_445_p
+ N_A_27_47#_c_300_n N_A_27_47#_c_301_n N_A_27_47#_c_302_n N_A_27_47#_c_287_n
+ N_A_27_47#_c_304_n N_A_27_47#_c_288_n PM_SKY130_FD_SC_HDLL__DFSTP_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%D N_D_c_537_n N_D_M1019_g N_D_M1017_g D D
+ N_D_c_539_n PM_SKY130_FD_SC_HDLL__DFSTP_4%D
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%A_211_363# N_A_211_363#_M1002_d
+ N_A_211_363#_M1032_d N_A_211_363#_c_593_n N_A_211_363#_c_594_n
+ N_A_211_363#_M1033_g N_A_211_363#_c_575_n N_A_211_363#_c_576_n
+ N_A_211_363#_M1021_g N_A_211_363#_c_578_n N_A_211_363#_c_597_n
+ N_A_211_363#_M1012_g N_A_211_363#_c_598_n N_A_211_363#_M1029_g
+ N_A_211_363#_c_580_n N_A_211_363#_c_581_n N_A_211_363#_c_582_n
+ N_A_211_363#_c_583_n N_A_211_363#_c_584_n N_A_211_363#_c_585_n
+ N_A_211_363#_c_586_n N_A_211_363#_c_587_n N_A_211_363#_c_588_n
+ N_A_211_363#_c_589_n N_A_211_363#_c_590_n N_A_211_363#_c_591_n
+ N_A_211_363#_c_592_n PM_SKY130_FD_SC_HDLL__DFSTP_4%A_211_363#
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%A_702_21# N_A_702_21#_M1030_d
+ N_A_702_21#_M1031_d N_A_702_21#_M1027_g N_A_702_21#_c_779_n
+ N_A_702_21#_M1010_g N_A_702_21#_c_780_n N_A_702_21#_c_858_p
+ N_A_702_21#_c_781_n N_A_702_21#_c_775_n N_A_702_21#_c_776_n
+ N_A_702_21#_c_783_n N_A_702_21#_c_784_n N_A_702_21#_c_777_n
+ PM_SKY130_FD_SC_HDLL__DFSTP_4%A_702_21#
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%SET_B N_SET_B_c_882_n N_SET_B_c_894_n
+ N_SET_B_M1031_g N_SET_B_M1026_g N_SET_B_M1037_g N_SET_B_c_895_n
+ N_SET_B_c_896_n N_SET_B_M1000_g N_SET_B_c_885_n N_SET_B_c_898_n
+ N_SET_B_c_886_n N_SET_B_c_887_n N_SET_B_c_888_n SET_B N_SET_B_c_889_n
+ N_SET_B_c_890_n N_SET_B_c_891_n N_SET_B_c_892_n
+ PM_SKY130_FD_SC_HDLL__DFSTP_4%SET_B
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%A_506_47# N_A_506_47#_M1003_d
+ N_A_506_47#_M1033_d N_A_506_47#_c_1012_n N_A_506_47#_M1030_g
+ N_A_506_47#_c_1013_n N_A_506_47#_c_1022_n N_A_506_47#_c_1023_n
+ N_A_506_47#_M1022_g N_A_506_47#_c_1014_n N_A_506_47#_c_1024_n
+ N_A_506_47#_c_1025_n N_A_506_47#_M1013_g N_A_506_47#_c_1015_n
+ N_A_506_47#_M1020_g N_A_506_47#_c_1016_n N_A_506_47#_c_1042_n
+ N_A_506_47#_c_1046_n N_A_506_47#_c_1026_n N_A_506_47#_c_1017_n
+ N_A_506_47#_c_1018_n N_A_506_47#_c_1019_n N_A_506_47#_c_1020_n
+ N_A_506_47#_c_1021_n PM_SKY130_FD_SC_HDLL__DFSTP_4%A_506_47#
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%A_1288_261# N_A_1288_261#_M1028_d
+ N_A_1288_261#_M1023_d N_A_1288_261#_c_1172_n N_A_1288_261#_M1011_g
+ N_A_1288_261#_M1034_g N_A_1288_261#_c_1205_p N_A_1288_261#_c_1174_n
+ N_A_1288_261#_c_1175_n N_A_1288_261#_c_1178_n N_A_1288_261#_c_1179_n
+ PM_SKY130_FD_SC_HDLL__DFSTP_4%A_1288_261#
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%A_1126_413# N_A_1126_413#_M1012_d
+ N_A_1126_413#_M1035_d N_A_1126_413#_M1000_s N_A_1126_413#_c_1254_n
+ N_A_1126_413#_M1023_g N_A_1126_413#_M1028_g N_A_1126_413#_c_1245_n
+ N_A_1126_413#_c_1246_n N_A_1126_413#_c_1257_n N_A_1126_413#_c_1258_n
+ N_A_1126_413#_M1009_g N_A_1126_413#_M1006_g N_A_1126_413#_c_1248_n
+ N_A_1126_413#_c_1267_n N_A_1126_413#_c_1260_n N_A_1126_413#_c_1275_n
+ N_A_1126_413#_c_1249_n N_A_1126_413#_c_1250_n N_A_1126_413#_c_1262_n
+ N_A_1126_413#_c_1251_n N_A_1126_413#_c_1263_n N_A_1126_413#_c_1264_n
+ N_A_1126_413#_c_1345_n N_A_1126_413#_c_1252_n N_A_1126_413#_c_1253_n
+ PM_SKY130_FD_SC_HDLL__DFSTP_4%A_1126_413#
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%A_1738_47# N_A_1738_47#_M1006_s
+ N_A_1738_47#_M1009_s N_A_1738_47#_M1001_g N_A_1738_47#_c_1416_n
+ N_A_1738_47#_M1004_g N_A_1738_47#_M1015_g N_A_1738_47#_c_1417_n
+ N_A_1738_47#_M1008_g N_A_1738_47#_M1016_g N_A_1738_47#_c_1418_n
+ N_A_1738_47#_M1014_g N_A_1738_47#_M1018_g N_A_1738_47#_c_1419_n
+ N_A_1738_47#_M1036_g N_A_1738_47#_c_1420_n N_A_1738_47#_M1038_g
+ N_A_1738_47#_M1039_g N_A_1738_47#_c_1412_n N_A_1738_47#_c_1413_n
+ N_A_1738_47#_c_1421_n N_A_1738_47#_c_1422_n N_A_1738_47#_c_1414_n
+ N_A_1738_47#_c_1415_n PM_SKY130_FD_SC_HDLL__DFSTP_4%A_1738_47#
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%VPWR N_VPWR_M1007_d N_VPWR_M1019_s
+ N_VPWR_M1010_d N_VPWR_M1022_d N_VPWR_M1011_d N_VPWR_M1000_d N_VPWR_M1009_d
+ N_VPWR_M1008_s N_VPWR_M1036_s N_VPWR_c_1533_n N_VPWR_c_1534_n N_VPWR_c_1535_n
+ N_VPWR_c_1536_n N_VPWR_c_1537_n N_VPWR_c_1538_n N_VPWR_c_1539_n
+ N_VPWR_c_1540_n N_VPWR_c_1541_n N_VPWR_c_1542_n N_VPWR_c_1543_n VPWR VPWR
+ N_VPWR_c_1544_n N_VPWR_c_1545_n N_VPWR_c_1546_n N_VPWR_c_1547_n
+ N_VPWR_c_1548_n N_VPWR_c_1549_n N_VPWR_c_1550_n N_VPWR_c_1532_n
+ N_VPWR_c_1552_n N_VPWR_c_1553_n N_VPWR_c_1554_n N_VPWR_c_1555_n
+ N_VPWR_c_1556_n N_VPWR_c_1557_n N_VPWR_c_1558_n
+ PM_SKY130_FD_SC_HDLL__DFSTP_4%VPWR
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%A_409_329# N_A_409_329#_M1017_d
+ N_A_409_329#_M1019_d N_A_409_329#_c_1728_n N_A_409_329#_c_1733_n
+ N_A_409_329#_c_1729_n N_A_409_329#_c_1735_n N_A_409_329#_c_1731_n
+ N_A_409_329#_c_1737_n N_A_409_329#_c_1738_n
+ PM_SKY130_FD_SC_HDLL__DFSTP_4%A_409_329#
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%Q N_Q_M1001_d N_Q_M1016_d N_Q_M1039_d
+ N_Q_M1004_d N_Q_M1014_d N_Q_M1038_d N_Q_c_1798_n N_Q_c_1799_n N_Q_c_1813_n
+ N_Q_c_1794_n N_Q_c_1821_n N_Q_c_1822_n N_Q_c_1824_n N_Q_c_1800_n N_Q_c_1795_n
+ N_Q_c_1801_n Q Q Q Q Q Q Q Q Q PM_SKY130_FD_SC_HDLL__DFSTP_4%Q
x_PM_SKY130_FD_SC_HDLL__DFSTP_4%VGND N_VGND_M1025_d N_VGND_M1017_s
+ N_VGND_M1027_d N_VGND_M1020_s N_VGND_M1037_d N_VGND_M1006_d N_VGND_M1015_s
+ N_VGND_M1018_s N_VGND_c_1884_n N_VGND_c_1885_n N_VGND_c_1886_n N_VGND_c_1887_n
+ N_VGND_c_1888_n N_VGND_c_1889_n N_VGND_c_1890_n N_VGND_c_1891_n VGND VGND
+ N_VGND_c_1892_n N_VGND_c_1893_n N_VGND_c_1894_n N_VGND_c_1895_n
+ N_VGND_c_1896_n N_VGND_c_1897_n N_VGND_c_1898_n N_VGND_c_1899_n
+ N_VGND_c_1900_n N_VGND_c_1901_n N_VGND_c_1902_n N_VGND_c_1903_n
+ N_VGND_c_1904_n N_VGND_c_1905_n N_VGND_c_1906_n
+ PM_SKY130_FD_SC_HDLL__DFSTP_4%VGND
cc_1 VNB N_CLK_c_234_n 0.0173562f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_2 VNB N_CLK_c_235_n 0.0271087f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_3 VNB CLK 0.0190034f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_CLK_c_237_n 0.0200763f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_CLK_c_238_n 0.0129466f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_6 VNB N_A_27_47#_M1002_g 0.0398926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_276_n 0.0187477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_277_n 0.0163574f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_9 VNB N_A_27_47#_c_278_n 0.00321162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_279_n 0.00649157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_280_n 0.0070415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_281_n 0.00517505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_282_n 0.0371442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_283_n 0.00720088f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_284_n 0.0105433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_285_n 0.0015872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_286_n 0.005579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_287_n 0.0263102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_288_n 0.0294618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_D_c_537_n 0.0289757f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_21 VNB N_D_M1017_g 0.0215162f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_22 VNB N_D_c_539_n 0.00504367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_211_363#_c_575_n 0.0147397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_211_363#_c_576_n 0.00518722f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_25 VNB N_A_211_363#_M1021_g 0.0207711f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_211_363#_c_578_n 0.00815197f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_27 VNB N_A_211_363#_M1012_g 0.0360314f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_28 VNB N_A_211_363#_c_580_n 0.0183966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_211_363#_c_581_n 0.0150246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_211_363#_c_582_n 0.0198942f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_31 VNB N_A_211_363#_c_583_n 0.00136753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_211_363#_c_584_n 0.001138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_211_363#_c_585_n 0.00547903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_211_363#_c_586_n 0.00188917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_211_363#_c_587_n 0.00588109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_211_363#_c_588_n 0.00137055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_211_363#_c_589_n 0.00223774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_211_363#_c_590_n 0.0167125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_211_363#_c_591_n 0.0253335f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_211_363#_c_592_n 0.0167983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_702_21#_M1027_g 0.0439852f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_42 VNB N_A_702_21#_c_775_n 0.00165887f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_43 VNB N_A_702_21#_c_776_n 0.00301395f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_44 VNB N_A_702_21#_c_777_n 0.00546105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_SET_B_c_882_n 0.00818253f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.07
cc_46 VNB N_SET_B_M1026_g 0.0187279f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_47 VNB N_SET_B_M1037_g 0.0193309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_SET_B_c_885_n 0.00846072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_SET_B_c_886_n 0.0136644f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_50 VNB N_SET_B_c_887_n 0.00264744f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_51 VNB N_SET_B_c_888_n 0.00136151f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_52 VNB N_SET_B_c_889_n 0.0347746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_SET_B_c_890_n 0.0288993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_SET_B_c_891_n 0.00798617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_SET_B_c_892_n 0.00955824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_506_47#_c_1012_n 0.0172275f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_57 VNB N_A_506_47#_c_1013_n 0.0151982f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_58 VNB N_A_506_47#_c_1014_n 0.0631852f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_59 VNB N_A_506_47#_c_1015_n 0.0183541f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_60 VNB N_A_506_47#_c_1016_n 0.00602262f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_61 VNB N_A_506_47#_c_1017_n 0.00495474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_506_47#_c_1018_n 0.00363504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_506_47#_c_1019_n 0.00317166f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_506_47#_c_1020_n 9.79949e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_506_47#_c_1021_n 0.0161521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1288_261#_c_1172_n 0.00882161f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=2.135
cc_67 VNB N_A_1288_261#_M1034_g 0.038132f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1288_261#_c_1174_n 0.00771946f $X=-0.19 $Y=-0.24 $X2=0.245
+ $Y2=1.235
cc_69 VNB N_A_1288_261#_c_1175_n 0.00532019f $X=-0.19 $Y=-0.24 $X2=0.265
+ $Y2=1.19
cc_70 VNB N_A_1126_413#_M1028_g 0.0340132f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_71 VNB N_A_1126_413#_c_1245_n 0.0405105f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=1.665
cc_72 VNB N_A_1126_413#_c_1246_n 0.016325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1126_413#_M1006_g 0.0390294f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_74 VNB N_A_1126_413#_c_1248_n 0.00782612f $X=-0.19 $Y=-0.24 $X2=0.265
+ $Y2=1.19
cc_75 VNB N_A_1126_413#_c_1249_n 0.00527277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1126_413#_c_1250_n 0.0010444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1126_413#_c_1251_n 0.0117159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1126_413#_c_1252_n 0.00111309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1126_413#_c_1253_n 0.0046917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1738_47#_M1001_g 0.0188836f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_81 VNB N_A_1738_47#_M1015_g 0.018541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1738_47#_M1016_g 0.0180317f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_83 VNB N_A_1738_47#_M1018_g 0.0190329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1738_47#_M1039_g 0.0215422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1738_47#_c_1412_n 0.0089403f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1738_47#_c_1413_n 0.0121201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1738_47#_c_1414_n 3.08128e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1738_47#_c_1415_n 0.11628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VPWR_c_1532_n 0.497461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_409_329#_c_1728_n 0.00900128f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_91 VNB N_A_409_329#_c_1729_n 0.00223047f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_92 VNB N_Q_c_1794_n 0.00109029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_Q_c_1795_n 0.00109029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB Q 0.0172698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB Q 0.0283742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1884_n 0.0191046f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_97 VNB N_VGND_c_1885_n 0.00784644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1886_n 0.0113467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1887_n 0.0053627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1888_n 0.00224717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1889_n 0.00241972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1890_n 0.0311849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1891_n 0.00545379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1892_n 0.0154125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1893_n 0.051238f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1894_n 0.0211095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1895_n 0.019446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1896_n 0.0136646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1897_n 0.014816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1898_n 0.556476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1899_n 0.00803343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1900_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1901_n 0.0109993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1902_n 0.00747262f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1903_n 0.0455124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1904_n 0.0123511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1905_n 0.00420355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1906_n 0.0060376f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VPB N_CLK_c_239_n 0.0103354f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_120 VPB N_CLK_c_240_n 0.0466088f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_121 VPB CLK 0.018034f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_122 VPB N_CLK_c_237_n 0.0102775f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_123 VPB N_A_27_47#_c_289_n 0.0173254f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_124 VPB N_A_27_47#_c_290_n 0.0249082f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_125 VPB N_A_27_47#_c_291_n 0.0537304f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_126 VPB N_A_27_47#_c_292_n 0.0544621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_27_47#_c_293_n 0.00146669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_47#_c_280_n 0.00397428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_27_47#_c_281_n 0.00304504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_283_n 0.00591262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_297_n 0.00356833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_298_n 0.00289349f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_299_n 0.0143045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_27_47#_c_300_n 0.00218288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_27_47#_c_301_n 0.00768004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_27_47#_c_302_n 0.0108096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_27_47#_c_287_n 0.012089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_27_47#_c_304_n 0.00751374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_D_c_537_n 0.0386914f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.88
cc_140 VPB N_D_c_539_n 0.00467649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_211_363#_c_593_n 0.0293669f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_142 VPB N_A_211_363#_c_594_n 0.0232248f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_143 VPB N_A_211_363#_c_575_n 0.0196158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_211_363#_c_576_n 0.00376696f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_145 VPB N_A_211_363#_c_597_n 0.0226062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_211_363#_c_598_n 0.0224575f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.07
cc_147 VPB N_A_211_363#_c_580_n 0.0126834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_211_363#_c_581_n 0.011213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_211_363#_c_589_n 0.00221192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_211_363#_c_592_n 0.0186828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_702_21#_M1027_g 0.0154962f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_152 VPB N_A_702_21#_c_779_n 0.0579237f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_153 VPB N_A_702_21#_c_780_n 0.00189103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_702_21#_c_781_n 0.00247793f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_155 VPB N_A_702_21#_c_776_n 0.00270641f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_156 VPB N_A_702_21#_c_783_n 0.00506096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_702_21#_c_784_n 0.00112185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_SET_B_c_882_n 0.0322461f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.07
cc_159 VPB N_SET_B_c_894_n 0.021903f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_160 VPB N_SET_B_c_895_n 0.0151303f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.665
cc_161 VPB N_SET_B_c_896_n 0.0275562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_SET_B_c_885_n 0.0135234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_SET_B_c_898_n 0.0107845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_506_47#_c_1022_n 0.0175131f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_165 VPB N_A_506_47#_c_1023_n 0.0204754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_506_47#_c_1024_n 0.0159914f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_167 VPB N_A_506_47#_c_1025_n 0.0208644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_506_47#_c_1026_n 0.0124261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_506_47#_c_1018_n 0.00559159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_506_47#_c_1019_n 0.00300162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_506_47#_c_1020_n 0.00266661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_506_47#_c_1021_n 0.0333235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_1288_261#_c_1172_n 0.0946401f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=2.135
cc_174 VPB N_A_1288_261#_c_1174_n 0.00312406f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_175 VPB N_A_1288_261#_c_1178_n 0.0183631f $X=-0.19 $Y=1.305 $X2=0.265
+ $Y2=1.53
cc_176 VPB N_A_1288_261#_c_1179_n 0.00841164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_1126_413#_c_1254_n 0.0191565f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.445
cc_178 VPB N_A_1126_413#_c_1245_n 0.0342965f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.665
cc_179 VPB N_A_1126_413#_c_1246_n 0.0191057f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_1126_413#_c_1257_n 0.0172705f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_181 VPB N_A_1126_413#_c_1258_n 0.0281414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_1126_413#_c_1248_n 0.00517032f $X=-0.19 $Y=1.305 $X2=0.265
+ $Y2=1.19
cc_183 VPB N_A_1126_413#_c_1260_n 0.00432852f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_1126_413#_c_1249_n 0.00190145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_1126_413#_c_1262_n 0.0151248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1126_413#_c_1263_n 0.00375313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1126_413#_c_1264_n 2.87011e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1126_413#_c_1252_n 2.77041e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1126_413#_c_1253_n 0.00450937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1738_47#_c_1416_n 0.0163846f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=0.805
cc_191 VPB N_A_1738_47#_c_1417_n 0.0160958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1738_47#_c_1418_n 0.0161f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_193 VPB N_A_1738_47#_c_1419_n 0.0159088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1738_47#_c_1420_n 0.01865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_1738_47#_c_1421_n 0.00608957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_1738_47#_c_1422_n 0.00369119f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_1738_47#_c_1415_n 0.0328308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1533_n 0.00108335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1534_n 0.0178983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1535_n 0.00592438f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1536_n 0.00259792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1537_n 0.00330976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1538_n 0.00400449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1539_n 4.16505e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1540_n 0.0216922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1541_n 0.00484211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1542_n 0.0159685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1543_n 0.00487564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1544_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1545_n 0.0467446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1546_n 0.0128873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1547_n 0.0346997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1548_n 0.0313059f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1549_n 0.0174648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1550_n 0.0154229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1532_n 0.068199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1552_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1553_n 0.00513751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1554_n 0.00930315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1555_n 0.00547467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1556_n 0.0131304f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1557_n 0.00538216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1558_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_409_329#_c_1728_n 0.00802517f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_225 VPB N_A_409_329#_c_1731_n 0.00186949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_Q_c_1798_n 0.00218429f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_227 VPB N_Q_c_1799_n 0.00166377f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_228 VPB N_Q_c_1800_n 0.00294772f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_Q_c_1801_n 0.00109154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB Q 0.00828363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB Q 0.0073261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB Q 0.0314153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 N_CLK_c_240_n N_A_27_47#_c_289_n 0.00668506f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_234 CLK N_A_27_47#_c_289_n 8.03089e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_235 N_CLK_c_237_n N_A_27_47#_c_289_n 0.00262072f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_236 N_CLK_c_240_n N_A_27_47#_c_290_n 0.0192779f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_237 N_CLK_c_234_n N_A_27_47#_M1002_g 0.0154184f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_238 N_CLK_c_238_n N_A_27_47#_M1002_g 0.00191451f $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_239 N_CLK_c_234_n N_A_27_47#_c_278_n 0.00643492f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_240 N_CLK_c_235_n N_A_27_47#_c_278_n 0.0108877f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_241 CLK N_A_27_47#_c_278_n 0.00736322f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_242 N_CLK_c_235_n N_A_27_47#_c_279_n 0.0059979f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_243 CLK N_A_27_47#_c_279_n 0.014414f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_244 N_CLK_c_237_n N_A_27_47#_c_279_n 3.2891e-19 $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_245 N_CLK_c_240_n N_A_27_47#_c_293_n 0.0171149f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_246 CLK N_A_27_47#_c_293_n 0.00731943f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_247 N_CLK_c_240_n N_A_27_47#_c_280_n 0.0042845f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_248 N_CLK_c_235_n N_A_27_47#_c_280_n 0.00196813f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_249 CLK N_A_27_47#_c_280_n 0.0429447f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_250 N_CLK_c_237_n N_A_27_47#_c_280_n 7.535e-19 $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_251 N_CLK_c_238_n N_A_27_47#_c_280_n 5.494e-19 $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_252 N_CLK_c_240_n N_A_27_47#_c_297_n 0.007998f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_253 CLK N_A_27_47#_c_297_n 0.0153363f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_254 N_CLK_c_237_n N_A_27_47#_c_297_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_255 N_CLK_c_240_n N_A_27_47#_c_298_n 0.00149934f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_256 CLK N_A_27_47#_c_287_n 0.00184424f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_257 N_CLK_c_237_n N_A_27_47#_c_287_n 0.0131201f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_258 N_CLK_c_240_n N_VPWR_c_1533_n 0.0125197f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_259 N_CLK_c_240_n N_VPWR_c_1544_n 0.00304525f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_260 N_CLK_c_240_n N_VPWR_c_1532_n 0.00454898f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_261 N_CLK_c_234_n N_VGND_c_1892_n 0.00198377f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_262 N_CLK_c_235_n N_VGND_c_1892_n 6.41851e-19 $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_263 N_CLK_c_234_n N_VGND_c_1898_n 0.00367064f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_264 N_CLK_c_234_n N_VGND_c_1899_n 0.0142867f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_281_n N_D_c_537_n 0.00124982f $X=2.585 $Y=0.87 $X2=-0.19
+ $Y2=-0.24
cc_266 N_A_27_47#_c_282_n N_D_c_537_n 0.00157653f $X=2.585 $Y=0.87 $X2=-0.19
+ $Y2=-0.24
cc_267 N_A_27_47#_c_304_n N_D_c_537_n 8.00147e-19 $X=2.965 $Y=1.74 $X2=-0.19
+ $Y2=-0.24
cc_268 N_A_27_47#_c_276_n N_D_M1017_g 0.0212193f $X=2.455 $Y=0.705 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_281_n N_D_M1017_g 0.0012111f $X=2.585 $Y=0.87 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_281_n N_D_c_539_n 0.0464864f $X=2.585 $Y=0.87 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_282_n N_D_c_539_n 2.44236e-19 $X=2.585 $Y=0.87 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_299_n N_D_c_539_n 0.00616551f $X=2.585 $Y=1.825 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_304_n N_D_c_539_n 0.00417777f $X=2.965 $Y=1.74 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_299_n N_A_211_363#_M1032_d 8.51638e-19 $X=2.585 $Y=1.825
+ $X2=0 $Y2=0
cc_275 N_A_27_47#_c_291_n N_A_211_363#_c_593_n 0.0229366f $X=2.96 $Y=1.99 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_281_n N_A_211_363#_c_593_n 0.00637191f $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_277 N_A_27_47#_c_299_n N_A_211_363#_c_593_n 0.00483233f $X=2.585 $Y=1.825
+ $X2=0 $Y2=0
cc_278 N_A_27_47#_c_304_n N_A_211_363#_c_593_n 0.0100464f $X=2.965 $Y=1.74 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_291_n N_A_211_363#_c_594_n 0.0128504f $X=2.96 $Y=1.99 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_299_n N_A_211_363#_c_594_n 0.00214786f $X=2.585 $Y=1.825
+ $X2=0 $Y2=0
cc_281 N_A_27_47#_c_304_n N_A_211_363#_c_594_n 0.00330305f $X=2.965 $Y=1.74
+ $X2=0 $Y2=0
cc_282 N_A_27_47#_c_291_n N_A_211_363#_c_575_n 0.0241913f $X=2.96 $Y=1.99 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_281_n N_A_211_363#_c_575_n 0.0105464f $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_302_n N_A_211_363#_c_575_n 3.63007e-19 $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_285 N_A_27_47#_c_304_n N_A_211_363#_c_575_n 0.00705057f $X=2.965 $Y=1.74
+ $X2=0 $Y2=0
cc_286 N_A_27_47#_c_281_n N_A_211_363#_c_576_n 0.00320692f $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_287 N_A_27_47#_c_282_n N_A_211_363#_c_576_n 0.0265243f $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_276_n N_A_211_363#_M1021_g 0.0140343f $X=2.455 $Y=0.705
+ $X2=0 $Y2=0
cc_289 N_A_27_47#_c_281_n N_A_211_363#_M1021_g 4.17219e-19 $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_290 N_A_27_47#_c_282_n N_A_211_363#_M1021_g 0.0166012f $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_292_n N_A_211_363#_c_597_n 0.0195155f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_283_n N_A_211_363#_c_597_n 0.0021791f $X=5.415 $Y=1.655
+ $X2=0 $Y2=0
cc_293 N_A_27_47#_c_300_n N_A_211_363#_c_597_n 0.00432834f $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_294 N_A_27_47#_c_301_n N_A_211_363#_c_597_n 0.0018637f $X=5.79 $Y=1.825 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_277_n N_A_211_363#_M1012_g 0.0172136f $X=6.645 $Y=0.765
+ $X2=0 $Y2=0
cc_296 N_A_27_47#_c_283_n N_A_211_363#_M1012_g 0.00363369f $X=5.415 $Y=1.655
+ $X2=0 $Y2=0
cc_297 N_A_27_47#_c_284_n N_A_211_363#_M1012_g 0.0116209f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_286_n N_A_211_363#_M1012_g 0.00278087f $X=6.56 $Y=0.81 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_288_n N_A_211_363#_M1012_g 0.0211955f $X=6.645 $Y=0.93 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_292_n N_A_211_363#_c_598_n 0.0138956f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_292_n N_A_211_363#_c_580_n 0.0106611f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_283_n N_A_211_363#_c_580_n 0.00351558f $X=5.415 $Y=1.655
+ $X2=0 $Y2=0
cc_303 N_A_27_47#_c_284_n N_A_211_363#_c_580_n 0.00554481f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_300_n N_A_211_363#_c_580_n 5.18898e-19 $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_305 N_A_27_47#_c_301_n N_A_211_363#_c_580_n 0.00101144f $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_306 N_A_27_47#_c_281_n N_A_211_363#_c_582_n 0.0204078f $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_282_n N_A_211_363#_c_582_n 0.00612283f $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_308 N_A_27_47#_c_281_n N_A_211_363#_c_583_n 0.00929355f $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_c_302_n N_A_211_363#_c_584_n 0.10518f $X=5.645 $Y=1.825 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_M1002_g N_A_211_363#_c_585_n 0.00656242f $X=0.99 $Y=0.445
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_c_278_n N_A_211_363#_c_585_n 0.00346684f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_280_n N_A_211_363#_c_585_n 0.00375448f $X=0.805 $Y=1.235
+ $X2=0 $Y2=0
cc_313 N_A_27_47#_c_281_n N_A_211_363#_c_586_n 3.82096e-19 $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_314 N_A_27_47#_c_276_n N_A_211_363#_c_587_n 5.45585e-19 $X=2.455 $Y=0.705
+ $X2=0 $Y2=0
cc_315 N_A_27_47#_c_291_n N_A_211_363#_c_587_n 3.45225e-19 $X=2.96 $Y=1.99 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_281_n N_A_211_363#_c_587_n 0.0212274f $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_282_n N_A_211_363#_c_587_n 0.0017744f $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_304_n N_A_211_363#_c_587_n 0.00520831f $X=2.965 $Y=1.74
+ $X2=0 $Y2=0
cc_319 N_A_27_47#_c_283_n N_A_211_363#_c_588_n 0.0024665f $X=5.415 $Y=1.655
+ $X2=0 $Y2=0
cc_320 N_A_27_47#_c_284_n N_A_211_363#_c_588_n 0.0014827f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_300_n N_A_211_363#_c_588_n 0.0144661f $X=5.79 $Y=1.825 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_301_n N_A_211_363#_c_588_n 0.00176238f $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_323 N_A_27_47#_c_292_n N_A_211_363#_c_589_n 6.19272e-19 $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_283_n N_A_211_363#_c_589_n 0.0226533f $X=5.415 $Y=1.655
+ $X2=0 $Y2=0
cc_325 N_A_27_47#_c_284_n N_A_211_363#_c_589_n 0.0123304f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_300_n N_A_211_363#_c_589_n 7.50589e-19 $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_301_n N_A_211_363#_c_589_n 0.0118448f $X=5.79 $Y=1.825 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_292_n N_A_211_363#_c_590_n 0.00131967f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_283_n N_A_211_363#_c_590_n 0.0125348f $X=5.415 $Y=1.655
+ $X2=0 $Y2=0
cc_330 N_A_27_47#_c_284_n N_A_211_363#_c_590_n 0.0022936f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_300_n N_A_211_363#_c_590_n 9.71873e-19 $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_c_301_n N_A_211_363#_c_590_n 0.00382035f $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_281_n N_A_211_363#_c_591_n 0.00696604f $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_c_290_n N_A_211_363#_c_592_n 0.00714312f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_M1002_g N_A_211_363#_c_592_n 0.0267456f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_278_n N_A_211_363#_c_592_n 0.00880333f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_402_p N_A_211_363#_c_592_n 0.00890502f $X=0.775 $Y=1.795
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_c_280_n N_A_211_363#_c_592_n 0.0584143f $X=0.805 $Y=1.235
+ $X2=0 $Y2=0
cc_339 N_A_27_47#_c_298_n N_A_211_363#_c_592_n 0.00215885f $X=0.895 $Y=1.825
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_c_299_n N_A_211_363#_c_592_n 0.0250011f $X=2.585 $Y=1.825
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_c_291_n N_A_702_21#_c_779_n 0.0250995f $X=2.96 $Y=1.99 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_302_n N_A_702_21#_c_779_n 0.00386067f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_c_302_n N_A_702_21#_c_780_n 0.0167093f $X=5.645 $Y=1.825 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_292_n N_A_702_21#_c_781_n 7.98086e-19 $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_301_n N_A_702_21#_c_781_n 0.00736761f $X=5.79 $Y=1.825 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_302_n N_A_702_21#_c_781_n 0.0238077f $X=5.645 $Y=1.825 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_292_n N_A_702_21#_c_776_n 2.1576e-19 $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_300_n N_A_702_21#_c_776_n 3.23422e-19 $X=5.79 $Y=1.825 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_301_n N_A_702_21#_c_776_n 0.0109818f $X=5.79 $Y=1.825 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_302_n N_A_702_21#_c_776_n 0.00695052f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_302_n N_A_702_21#_c_783_n 0.0185377f $X=5.645 $Y=1.825 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_302_n N_A_702_21#_c_784_n 0.00782494f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_283_n N_A_702_21#_c_777_n 0.0448021f $X=5.415 $Y=1.655 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_285_n N_A_702_21#_c_777_n 0.00932877f $X=5.5 $Y=0.81 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_302_n N_SET_B_c_882_n 0.00261058f $X=5.645 $Y=1.825 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_283_n N_SET_B_c_886_n 0.00404989f $X=5.415 $Y=1.655 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_284_n N_SET_B_c_886_n 0.0343911f $X=6.37 $Y=0.81 $X2=0 $Y2=0
cc_358 N_A_27_47#_c_285_n N_SET_B_c_886_n 0.00603182f $X=5.5 $Y=0.81 $X2=0 $Y2=0
cc_359 N_A_27_47#_c_286_n N_SET_B_c_886_n 0.0189103f $X=6.56 $Y=0.81 $X2=0 $Y2=0
cc_360 N_A_27_47#_c_302_n N_A_506_47#_c_1022_n 0.0023633f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_292_n N_A_506_47#_c_1014_n 0.0031094f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_283_n N_A_506_47#_c_1014_n 0.00474618f $X=5.415 $Y=1.655
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_284_n N_A_506_47#_c_1014_n 0.0102775f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_285_n N_A_506_47#_c_1014_n 0.00679842f $X=5.5 $Y=0.81 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_292_n N_A_506_47#_c_1024_n 0.024165f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_301_n N_A_506_47#_c_1024_n 0.00202479f $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_367 N_A_27_47#_c_302_n N_A_506_47#_c_1024_n 0.00251704f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_c_292_n N_A_506_47#_c_1025_n 0.0361774f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_302_n N_A_506_47#_c_1025_n 0.00220794f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_284_n N_A_506_47#_c_1015_n 0.00416353f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_291_n N_A_506_47#_c_1042_n 0.0124798f $X=2.96 $Y=1.99 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_299_n N_A_506_47#_c_1042_n 0.00261149f $X=2.585 $Y=1.825
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_302_n N_A_506_47#_c_1042_n 0.00443131f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_304_n N_A_506_47#_c_1042_n 0.0193114f $X=2.965 $Y=1.74 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_276_n N_A_506_47#_c_1046_n 0.00335745f $X=2.455 $Y=0.705
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_281_n N_A_506_47#_c_1046_n 0.0070258f $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_282_n N_A_506_47#_c_1046_n 9.58359e-19 $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_291_n N_A_506_47#_c_1026_n 0.00861559f $X=2.96 $Y=1.99 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_281_n N_A_506_47#_c_1026_n 0.00628894f $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_445_p N_A_506_47#_c_1026_n 4.07831e-19 $X=2.875 $Y=1.825
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_302_n N_A_506_47#_c_1026_n 0.013911f $X=5.645 $Y=1.825 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_304_n N_A_506_47#_c_1026_n 0.0285215f $X=2.965 $Y=1.74 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_302_n N_A_506_47#_c_1018_n 0.00512083f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_281_n N_A_506_47#_c_1019_n 0.00597075f $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_385 N_A_27_47#_c_302_n N_A_506_47#_c_1019_n 0.00458729f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_302_n N_A_506_47#_c_1020_n 0.00296278f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_c_283_n N_A_506_47#_c_1021_n 0.00786821f $X=5.415 $Y=1.655
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_302_n N_A_506_47#_c_1021_n 0.00148193f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_389 N_A_27_47#_c_286_n N_A_1288_261#_c_1172_n 4.44985e-19 $X=6.56 $Y=0.81
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_c_288_n N_A_1288_261#_c_1172_n 0.0180537f $X=6.645 $Y=0.93
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_277_n N_A_1288_261#_M1034_g 0.0628903f $X=6.645 $Y=0.765
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_c_286_n N_A_1288_261#_M1034_g 8.58205e-19 $X=6.56 $Y=0.81
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_292_n N_A_1126_413#_c_1267_n 0.00794725f $X=5.54 $Y=1.99
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_300_n N_A_1126_413#_c_1267_n 0.00109575f $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_301_n N_A_1126_413#_c_1267_n 0.0183376f $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_c_302_n N_A_1126_413#_c_1267_n 0.00152637f $X=5.645 $Y=1.825
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_292_n N_A_1126_413#_c_1260_n 5.01151e-19 $X=5.54 $Y=1.99
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_c_283_n N_A_1126_413#_c_1260_n 0.00507933f $X=5.415 $Y=1.655
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_300_n N_A_1126_413#_c_1260_n 0.00742868f $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_301_n N_A_1126_413#_c_1260_n 0.0212476f $X=5.79 $Y=1.825
+ $X2=0 $Y2=0
cc_401 N_A_27_47#_c_277_n N_A_1126_413#_c_1275_n 0.0104344f $X=6.645 $Y=0.765
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_284_n N_A_1126_413#_c_1275_n 0.00680222f $X=6.37 $Y=0.81
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_286_n N_A_1126_413#_c_1275_n 0.0150149f $X=6.56 $Y=0.81
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_c_288_n N_A_1126_413#_c_1275_n 8.69648e-19 $X=6.645 $Y=0.93
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_284_n N_A_1126_413#_c_1249_n 0.00259385f $X=6.37 $Y=0.81
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_286_n N_A_1126_413#_c_1249_n 0.0210672f $X=6.56 $Y=0.81
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_288_n N_A_1126_413#_c_1249_n 0.00278641f $X=6.645 $Y=0.93
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_284_n N_A_1126_413#_c_1250_n 0.00719613f $X=6.37 $Y=0.81
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_277_n N_A_1126_413#_c_1251_n 0.00248785f $X=6.645 $Y=0.765
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_286_n N_A_1126_413#_c_1251_n 0.0220255f $X=6.56 $Y=0.81
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_288_n N_A_1126_413#_c_1251_n 0.00157366f $X=6.645 $Y=0.93
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_c_292_n N_A_1126_413#_c_1264_n 0.00102409f $X=5.54 $Y=1.99
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_402_p N_VPWR_M1007_d 0.00171205f $X=0.775 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_414 N_A_27_47#_c_290_n N_VPWR_c_1533_n 0.00859878f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_293_n N_VPWR_c_1533_n 0.00629408f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_402_p N_VPWR_c_1533_n 0.0135522f $X=0.775 $Y=1.795 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_297_n N_VPWR_c_1533_n 0.0246493f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_418 N_A_27_47#_c_298_n N_VPWR_c_1533_n 0.0014373f $X=0.895 $Y=1.825 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_290_n N_VPWR_c_1534_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_290_n N_VPWR_c_1535_n 0.00191848f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_299_n N_VPWR_c_1535_n 0.0016741f $X=2.585 $Y=1.825 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_293_n N_VPWR_c_1544_n 0.00180073f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_297_n N_VPWR_c_1544_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_424 N_A_27_47#_c_291_n N_VPWR_c_1545_n 0.00440543f $X=2.96 $Y=1.99 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_c_292_n N_VPWR_c_1547_n 0.00510448f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_c_301_n N_VPWR_c_1547_n 0.0032218f $X=5.79 $Y=1.825 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_c_290_n N_VPWR_c_1532_n 0.00665316f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_291_n N_VPWR_c_1532_n 0.00645014f $X=2.96 $Y=1.99 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_c_292_n N_VPWR_c_1532_n 0.00671662f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_c_293_n N_VPWR_c_1532_n 0.00426237f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_c_402_p N_VPWR_c_1532_n 5.98513e-19 $X=0.775 $Y=1.795 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_c_297_n N_VPWR_c_1532_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_c_298_n N_VPWR_c_1532_n 0.244302f $X=0.895 $Y=1.825 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_301_n N_VPWR_c_1532_n 0.00309512f $X=5.79 $Y=1.825 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_c_304_n N_VPWR_c_1532_n 0.0018449f $X=2.965 $Y=1.74 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_302_n N_VPWR_c_1554_n 0.00143103f $X=5.645 $Y=1.825 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_292_n N_VPWR_c_1555_n 0.00179407f $X=5.54 $Y=1.99 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_c_302_n N_VPWR_c_1555_n 0.0013893f $X=5.645 $Y=1.825 $X2=0
+ $Y2=0
cc_439 N_A_27_47#_c_299_n N_A_409_329#_M1019_d 8.84929e-19 $X=2.585 $Y=1.825
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_276_n N_A_409_329#_c_1733_n 0.00230176f $X=2.455 $Y=0.705
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_281_n N_A_409_329#_c_1733_n 0.00719598f $X=2.585 $Y=0.87
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_c_299_n N_A_409_329#_c_1735_n 0.021266f $X=2.585 $Y=1.825
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_c_299_n N_A_409_329#_c_1731_n 0.0157331f $X=2.585 $Y=1.825
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_276_n N_A_409_329#_c_1737_n 0.00409202f $X=2.455 $Y=0.705
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_299_n N_A_409_329#_c_1738_n 0.010951f $X=2.585 $Y=1.825
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_304_n N_A_409_329#_c_1738_n 0.00841982f $X=2.965 $Y=1.74
+ $X2=0 $Y2=0
cc_447 N_A_27_47#_c_278_n N_VGND_M1025_d 0.00227127f $X=0.66 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_448 N_A_27_47#_M1002_g N_VGND_c_1884_n 0.00585385f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_M1002_g N_VGND_c_1885_n 0.0030195f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_284_n N_VGND_c_1886_n 0.00194189f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_285_n N_VGND_c_1886_n 0.0129707f $X=5.5 $Y=0.81 $X2=0 $Y2=0
cc_452 N_A_27_47#_c_517_p N_VGND_c_1892_n 0.00725596f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_c_278_n N_VGND_c_1892_n 0.00244154f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_276_n N_VGND_c_1893_n 0.00556304f $X=2.455 $Y=0.705 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_281_n N_VGND_c_1893_n 0.00190868f $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_282_n N_VGND_c_1893_n 4.30307e-19 $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_M1025_s N_VGND_c_1898_n 0.00437169f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_M1002_g N_VGND_c_1898_n 0.0120602f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_276_n N_VGND_c_1898_n 0.00696803f $X=2.455 $Y=0.705 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_277_n N_VGND_c_1898_n 0.00537645f $X=6.645 $Y=0.765 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_517_p N_VGND_c_1898_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_278_n N_VGND_c_1898_n 0.00625251f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_281_n N_VGND_c_1898_n 0.00182252f $X=2.585 $Y=0.87 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_284_n N_VGND_c_1898_n 0.00729594f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_c_285_n N_VGND_c_1898_n 4.92512e-19 $X=5.5 $Y=0.81 $X2=0 $Y2=0
cc_466 N_A_27_47#_M1002_g N_VGND_c_1899_n 0.00176556f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_c_517_p N_VGND_c_1899_n 0.00895866f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_278_n N_VGND_c_1899_n 0.0228644f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_469 N_A_27_47#_c_287_n N_VGND_c_1899_n 6.84207e-19 $X=0.99 $Y=1.235 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_277_n N_VGND_c_1903_n 0.00368123f $X=6.645 $Y=0.765 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_284_n N_VGND_c_1903_n 0.00949562f $X=6.37 $Y=0.81 $X2=0
+ $Y2=0
cc_472 N_D_c_537_n N_A_211_363#_c_593_n 0.0105647f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_473 N_D_c_537_n N_A_211_363#_c_594_n 0.0114995f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_474 N_D_c_537_n N_A_211_363#_c_576_n 0.0123596f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_475 N_D_c_539_n N_A_211_363#_c_576_n 0.00343431f $X=1.955 $Y=1.17 $X2=0 $Y2=0
cc_476 N_D_c_537_n N_A_211_363#_c_582_n 0.00134388f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_477 N_D_M1017_g N_A_211_363#_c_582_n 0.00343113f $X=1.98 $Y=0.555 $X2=0 $Y2=0
cc_478 N_D_c_539_n N_A_211_363#_c_582_n 0.0140774f $X=1.955 $Y=1.17 $X2=0 $Y2=0
cc_479 N_D_c_537_n N_A_211_363#_c_592_n 0.00436322f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_480 N_D_M1017_g N_A_211_363#_c_592_n 0.0036787f $X=1.98 $Y=0.555 $X2=0 $Y2=0
cc_481 N_D_c_537_n N_VPWR_c_1535_n 0.0117702f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_482 N_D_c_537_n N_VPWR_c_1545_n 0.00470513f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_483 N_D_c_537_n N_VPWR_c_1532_n 0.00518371f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_484 N_D_c_537_n N_A_409_329#_c_1728_n 0.0196745f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_485 N_D_M1017_g N_A_409_329#_c_1728_n 0.00519391f $X=1.98 $Y=0.555 $X2=0
+ $Y2=0
cc_486 N_D_c_539_n N_A_409_329#_c_1728_n 0.0477681f $X=1.955 $Y=1.17 $X2=0 $Y2=0
cc_487 N_D_c_537_n N_A_409_329#_c_1733_n 0.00230232f $X=1.955 $Y=1.57 $X2=0
+ $Y2=0
cc_488 N_D_M1017_g N_A_409_329#_c_1733_n 0.012828f $X=1.98 $Y=0.555 $X2=0 $Y2=0
cc_489 N_D_c_539_n N_A_409_329#_c_1733_n 0.024373f $X=1.955 $Y=1.17 $X2=0 $Y2=0
cc_490 N_D_c_537_n N_A_409_329#_c_1735_n 0.0133332f $X=1.955 $Y=1.57 $X2=0 $Y2=0
cc_491 N_D_c_539_n N_A_409_329#_c_1735_n 0.0140214f $X=1.955 $Y=1.17 $X2=0 $Y2=0
cc_492 N_D_c_539_n N_A_409_329#_c_1738_n 0.0140554f $X=1.955 $Y=1.17 $X2=0 $Y2=0
cc_493 N_D_M1017_g N_VGND_c_1885_n 0.00482545f $X=1.98 $Y=0.555 $X2=0 $Y2=0
cc_494 N_D_M1017_g N_VGND_c_1893_n 0.00425094f $X=1.98 $Y=0.555 $X2=0 $Y2=0
cc_495 N_D_M1017_g N_VGND_c_1898_n 0.00685456f $X=1.98 $Y=0.555 $X2=0 $Y2=0
cc_496 N_A_211_363#_M1021_g N_A_702_21#_M1027_g 0.0246593f $X=3.105 $Y=0.415
+ $X2=0 $Y2=0
cc_497 N_A_211_363#_c_578_n N_A_702_21#_M1027_g 0.0115768f $X=3.105 $Y=1.245
+ $X2=0 $Y2=0
cc_498 N_A_211_363#_c_586_n N_A_702_21#_M1027_g 0.00698184f $X=3.24 $Y=0.805
+ $X2=0 $Y2=0
cc_499 N_A_211_363#_c_587_n N_A_702_21#_M1027_g 0.00189271f $X=3.24 $Y=0.805
+ $X2=0 $Y2=0
cc_500 N_A_211_363#_c_590_n N_A_702_21#_M1027_g 0.00125199f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_501 N_A_211_363#_c_591_n N_A_702_21#_M1027_g 0.0200904f $X=3.165 $Y=0.93
+ $X2=0 $Y2=0
cc_502 N_A_211_363#_c_590_n N_A_702_21#_c_780_n 6.57625e-19 $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_503 N_A_211_363#_c_590_n N_A_702_21#_c_781_n 0.00123565f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_504 N_A_211_363#_c_590_n N_A_702_21#_c_776_n 0.015874f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_505 N_A_211_363#_c_590_n N_A_702_21#_c_783_n 0.00100416f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_506 N_A_211_363#_c_590_n N_A_702_21#_c_777_n 0.00569788f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_507 N_A_211_363#_c_590_n N_SET_B_c_882_n 0.00130401f $X=5.665 $Y=1.195 $X2=0
+ $Y2=0
cc_508 N_A_211_363#_M1012_g N_SET_B_c_886_n 0.00283363f $X=6.115 $Y=0.445 $X2=0
+ $Y2=0
cc_509 N_A_211_363#_c_580_n N_SET_B_c_886_n 0.00242505f $X=5.97 $Y=1.26 $X2=0
+ $Y2=0
cc_510 N_A_211_363#_c_588_n N_SET_B_c_886_n 0.0265487f $X=5.81 $Y=1.195 $X2=0
+ $Y2=0
cc_511 N_A_211_363#_c_589_n N_SET_B_c_886_n 0.00114117f $X=5.81 $Y=1.195 $X2=0
+ $Y2=0
cc_512 N_A_211_363#_c_590_n N_SET_B_c_886_n 0.0918817f $X=5.665 $Y=1.195 $X2=0
+ $Y2=0
cc_513 N_A_211_363#_c_590_n N_SET_B_c_887_n 0.0262012f $X=5.665 $Y=1.195 $X2=0
+ $Y2=0
cc_514 N_A_211_363#_c_590_n N_SET_B_c_889_n 0.00449551f $X=5.665 $Y=1.195 $X2=0
+ $Y2=0
cc_515 N_A_211_363#_c_590_n N_SET_B_c_892_n 0.00996743f $X=5.665 $Y=1.195 $X2=0
+ $Y2=0
cc_516 N_A_211_363#_c_590_n N_A_506_47#_c_1013_n 0.0032089f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_517 N_A_211_363#_c_580_n N_A_506_47#_c_1014_n 0.00912806f $X=5.97 $Y=1.26
+ $X2=0 $Y2=0
cc_518 N_A_211_363#_c_589_n N_A_506_47#_c_1014_n 3.19592e-19 $X=5.81 $Y=1.195
+ $X2=0 $Y2=0
cc_519 N_A_211_363#_c_590_n N_A_506_47#_c_1014_n 0.00138939f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_520 N_A_211_363#_M1012_g N_A_506_47#_c_1015_n 0.0412678f $X=6.115 $Y=0.445
+ $X2=0 $Y2=0
cc_521 N_A_211_363#_c_594_n N_A_506_47#_c_1042_n 0.00459362f $X=2.49 $Y=1.99
+ $X2=0 $Y2=0
cc_522 N_A_211_363#_M1021_g N_A_506_47#_c_1046_n 0.0120266f $X=3.105 $Y=0.415
+ $X2=0 $Y2=0
cc_523 N_A_211_363#_c_582_n N_A_506_47#_c_1046_n 0.00591552f $X=3.095 $Y=0.85
+ $X2=0 $Y2=0
cc_524 N_A_211_363#_c_586_n N_A_506_47#_c_1046_n 0.00205557f $X=3.24 $Y=0.805
+ $X2=0 $Y2=0
cc_525 N_A_211_363#_c_587_n N_A_506_47#_c_1046_n 0.0218855f $X=3.24 $Y=0.805
+ $X2=0 $Y2=0
cc_526 N_A_211_363#_c_591_n N_A_506_47#_c_1046_n 5.24271e-19 $X=3.165 $Y=0.93
+ $X2=0 $Y2=0
cc_527 N_A_211_363#_c_593_n N_A_506_47#_c_1026_n 8.38684e-19 $X=2.49 $Y=1.89
+ $X2=0 $Y2=0
cc_528 N_A_211_363#_c_584_n N_A_506_47#_c_1026_n 3.06581e-19 $X=3.385 $Y=1.19
+ $X2=0 $Y2=0
cc_529 N_A_211_363#_M1021_g N_A_506_47#_c_1017_n 0.00118384f $X=3.105 $Y=0.415
+ $X2=0 $Y2=0
cc_530 N_A_211_363#_c_578_n N_A_506_47#_c_1017_n 0.00109256f $X=3.105 $Y=1.245
+ $X2=0 $Y2=0
cc_531 N_A_211_363#_c_586_n N_A_506_47#_c_1017_n 0.0149193f $X=3.24 $Y=0.805
+ $X2=0 $Y2=0
cc_532 N_A_211_363#_c_587_n N_A_506_47#_c_1017_n 0.0244314f $X=3.24 $Y=0.805
+ $X2=0 $Y2=0
cc_533 N_A_211_363#_c_590_n N_A_506_47#_c_1017_n 0.0205647f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_534 N_A_211_363#_c_591_n N_A_506_47#_c_1017_n 7.7085e-19 $X=3.165 $Y=0.93
+ $X2=0 $Y2=0
cc_535 N_A_211_363#_c_590_n N_A_506_47#_c_1018_n 0.0226579f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_536 N_A_211_363#_c_578_n N_A_506_47#_c_1019_n 0.00242434f $X=3.105 $Y=1.245
+ $X2=0 $Y2=0
cc_537 N_A_211_363#_c_584_n N_A_506_47#_c_1019_n 0.00466397f $X=3.385 $Y=1.19
+ $X2=0 $Y2=0
cc_538 N_A_211_363#_c_587_n N_A_506_47#_c_1019_n 0.00439529f $X=3.24 $Y=0.805
+ $X2=0 $Y2=0
cc_539 N_A_211_363#_c_590_n N_A_506_47#_c_1019_n 0.0108475f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_540 N_A_211_363#_c_591_n N_A_506_47#_c_1019_n 5.43524e-19 $X=3.165 $Y=0.93
+ $X2=0 $Y2=0
cc_541 N_A_211_363#_c_590_n N_A_506_47#_c_1020_n 0.0119084f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_542 N_A_211_363#_c_580_n N_A_506_47#_c_1021_n 0.00408857f $X=5.97 $Y=1.26
+ $X2=0 $Y2=0
cc_543 N_A_211_363#_c_590_n N_A_506_47#_c_1021_n 0.00509204f $X=5.665 $Y=1.195
+ $X2=0 $Y2=0
cc_544 N_A_211_363#_c_598_n N_A_1288_261#_c_1172_n 0.0350643f $X=6.13 $Y=1.99
+ $X2=0 $Y2=0
cc_545 N_A_211_363#_c_581_n N_A_1288_261#_c_1172_n 0.0431735f $X=5.97 $Y=1.125
+ $X2=0 $Y2=0
cc_546 N_A_211_363#_c_598_n N_A_1126_413#_c_1267_n 0.00702778f $X=6.13 $Y=1.99
+ $X2=0 $Y2=0
cc_547 N_A_211_363#_c_597_n N_A_1126_413#_c_1260_n 0.011905f $X=6.13 $Y=1.89
+ $X2=0 $Y2=0
cc_548 N_A_211_363#_c_598_n N_A_1126_413#_c_1260_n 5.64786e-19 $X=6.13 $Y=1.99
+ $X2=0 $Y2=0
cc_549 N_A_211_363#_c_581_n N_A_1126_413#_c_1260_n 0.00126981f $X=5.97 $Y=1.125
+ $X2=0 $Y2=0
cc_550 N_A_211_363#_c_589_n N_A_1126_413#_c_1260_n 0.00505459f $X=5.81 $Y=1.195
+ $X2=0 $Y2=0
cc_551 N_A_211_363#_c_581_n N_A_1126_413#_c_1250_n 0.010381f $X=5.97 $Y=1.125
+ $X2=0 $Y2=0
cc_552 N_A_211_363#_c_588_n N_A_1126_413#_c_1250_n 0.00214482f $X=5.81 $Y=1.195
+ $X2=0 $Y2=0
cc_553 N_A_211_363#_c_589_n N_A_1126_413#_c_1250_n 0.0122615f $X=5.81 $Y=1.195
+ $X2=0 $Y2=0
cc_554 N_A_211_363#_c_598_n N_A_1126_413#_c_1262_n 2.46208e-19 $X=6.13 $Y=1.99
+ $X2=0 $Y2=0
cc_555 N_A_211_363#_c_598_n N_A_1126_413#_c_1264_n 0.0149113f $X=6.13 $Y=1.99
+ $X2=0 $Y2=0
cc_556 N_A_211_363#_c_592_n N_VPWR_c_1533_n 0.0206383f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_557 N_A_211_363#_c_592_n N_VPWR_c_1534_n 0.015988f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_558 N_A_211_363#_c_594_n N_VPWR_c_1535_n 0.0010427f $X=2.49 $Y=1.99 $X2=0
+ $Y2=0
cc_559 N_A_211_363#_c_592_n N_VPWR_c_1535_n 0.0226553f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_560 N_A_211_363#_c_594_n N_VPWR_c_1545_n 0.00621307f $X=2.49 $Y=1.99 $X2=0
+ $Y2=0
cc_561 N_A_211_363#_c_598_n N_VPWR_c_1547_n 0.00445421f $X=6.13 $Y=1.99 $X2=0
+ $Y2=0
cc_562 N_A_211_363#_c_594_n N_VPWR_c_1532_n 0.00724577f $X=2.49 $Y=1.99 $X2=0
+ $Y2=0
cc_563 N_A_211_363#_c_598_n N_VPWR_c_1532_n 0.00628429f $X=6.13 $Y=1.99 $X2=0
+ $Y2=0
cc_564 N_A_211_363#_c_592_n N_VPWR_c_1532_n 0.00409094f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_565 N_A_211_363#_c_598_n N_VPWR_c_1556_n 0.00199481f $X=6.13 $Y=1.99 $X2=0
+ $Y2=0
cc_566 N_A_211_363#_c_582_n N_A_409_329#_M1017_d 4.25819e-19 $X=3.095 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_567 N_A_211_363#_c_582_n N_A_409_329#_c_1728_n 0.0148354f $X=3.095 $Y=0.85
+ $X2=0 $Y2=0
cc_568 N_A_211_363#_c_592_n N_A_409_329#_c_1728_n 0.0682158f $X=1.2 $Y=0.51
+ $X2=0 $Y2=0
cc_569 N_A_211_363#_c_582_n N_A_409_329#_c_1733_n 0.0214599f $X=3.095 $Y=0.85
+ $X2=0 $Y2=0
cc_570 N_A_211_363#_c_587_n N_A_409_329#_c_1733_n 0.00191581f $X=3.24 $Y=0.805
+ $X2=0 $Y2=0
cc_571 N_A_211_363#_c_582_n N_A_409_329#_c_1729_n 0.00435851f $X=3.095 $Y=0.85
+ $X2=0 $Y2=0
cc_572 N_A_211_363#_c_585_n N_A_409_329#_c_1729_n 0.00280684f $X=1.395 $Y=0.805
+ $X2=0 $Y2=0
cc_573 N_A_211_363#_c_592_n N_A_409_329#_c_1729_n 0.0131564f $X=1.2 $Y=0.51
+ $X2=0 $Y2=0
cc_574 N_A_211_363#_c_592_n N_A_409_329#_c_1731_n 0.0115156f $X=1.2 $Y=0.51
+ $X2=0 $Y2=0
cc_575 N_A_211_363#_c_593_n N_A_409_329#_c_1738_n 0.00147341f $X=2.49 $Y=1.89
+ $X2=0 $Y2=0
cc_576 N_A_211_363#_c_594_n N_A_409_329#_c_1738_n 0.00891072f $X=2.49 $Y=1.99
+ $X2=0 $Y2=0
cc_577 N_A_211_363#_c_585_n N_VGND_c_1884_n 5.1806e-19 $X=1.395 $Y=0.805 $X2=0
+ $Y2=0
cc_578 N_A_211_363#_c_592_n N_VGND_c_1884_n 0.00978627f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_579 N_A_211_363#_c_582_n N_VGND_c_1885_n 0.00124768f $X=3.095 $Y=0.85 $X2=0
+ $Y2=0
cc_580 N_A_211_363#_c_592_n N_VGND_c_1885_n 0.00823833f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_581 N_A_211_363#_M1021_g N_VGND_c_1893_n 0.00359964f $X=3.105 $Y=0.415 $X2=0
+ $Y2=0
cc_582 N_A_211_363#_M1002_d N_VGND_c_1898_n 0.0031895f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_583 N_A_211_363#_M1021_g N_VGND_c_1898_n 0.00584151f $X=3.105 $Y=0.415 $X2=0
+ $Y2=0
cc_584 N_A_211_363#_M1012_g N_VGND_c_1898_n 0.00595652f $X=6.115 $Y=0.445 $X2=0
+ $Y2=0
cc_585 N_A_211_363#_c_582_n N_VGND_c_1898_n 0.079188f $X=3.095 $Y=0.85 $X2=0
+ $Y2=0
cc_586 N_A_211_363#_c_585_n N_VGND_c_1898_n 0.0161996f $X=1.395 $Y=0.805 $X2=0
+ $Y2=0
cc_587 N_A_211_363#_c_586_n N_VGND_c_1898_n 0.0163517f $X=3.24 $Y=0.805 $X2=0
+ $Y2=0
cc_588 N_A_211_363#_c_592_n N_VGND_c_1898_n 0.00355424f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_589 N_A_211_363#_M1012_g N_VGND_c_1903_n 0.00437852f $X=6.115 $Y=0.445 $X2=0
+ $Y2=0
cc_590 N_A_211_363#_c_587_n A_636_47# 0.00109504f $X=3.24 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_591 N_A_702_21#_M1027_g N_SET_B_c_882_n 0.0119034f $X=3.585 $Y=0.445 $X2=0
+ $Y2=0
cc_592 N_A_702_21#_c_779_n N_SET_B_c_882_n 0.020463f $X=3.61 $Y=1.99 $X2=0 $Y2=0
cc_593 N_A_702_21#_c_780_n N_SET_B_c_882_n 0.00517985f $X=4.34 $Y=1.96 $X2=0
+ $Y2=0
cc_594 N_A_702_21#_c_783_n N_SET_B_c_882_n 0.00575143f $X=3.695 $Y=1.74 $X2=0
+ $Y2=0
cc_595 N_A_702_21#_c_779_n N_SET_B_c_894_n 0.0156789f $X=3.61 $Y=1.99 $X2=0
+ $Y2=0
cc_596 N_A_702_21#_c_780_n N_SET_B_c_894_n 0.0117591f $X=4.34 $Y=1.96 $X2=0
+ $Y2=0
cc_597 N_A_702_21#_M1027_g N_SET_B_M1026_g 0.0101173f $X=3.585 $Y=0.445 $X2=0
+ $Y2=0
cc_598 N_A_702_21#_c_777_n N_SET_B_c_886_n 0.0201744f $X=4.95 $Y=1.065 $X2=0
+ $Y2=0
cc_599 N_A_702_21#_c_777_n N_SET_B_c_887_n 6.43658e-19 $X=4.95 $Y=1.065 $X2=0
+ $Y2=0
cc_600 N_A_702_21#_M1027_g N_SET_B_c_889_n 0.0148962f $X=3.585 $Y=0.445 $X2=0
+ $Y2=0
cc_601 N_A_702_21#_c_776_n N_SET_B_c_889_n 6.99938e-19 $X=5.025 $Y=1.835 $X2=0
+ $Y2=0
cc_602 N_A_702_21#_c_777_n N_SET_B_c_889_n 2.45403e-19 $X=4.95 $Y=1.065 $X2=0
+ $Y2=0
cc_603 N_A_702_21#_M1027_g N_SET_B_c_892_n 0.00109852f $X=3.585 $Y=0.445 $X2=0
+ $Y2=0
cc_604 N_A_702_21#_c_777_n N_SET_B_c_892_n 0.015565f $X=4.95 $Y=1.065 $X2=0
+ $Y2=0
cc_605 N_A_702_21#_c_775_n N_A_506_47#_c_1012_n 0.00666987f $X=4.875 $Y=0.46
+ $X2=0 $Y2=0
cc_606 N_A_702_21#_c_776_n N_A_506_47#_c_1013_n 0.00252146f $X=5.025 $Y=1.835
+ $X2=0 $Y2=0
cc_607 N_A_702_21#_c_777_n N_A_506_47#_c_1013_n 0.00155564f $X=4.95 $Y=1.065
+ $X2=0 $Y2=0
cc_608 N_A_702_21#_c_781_n N_A_506_47#_c_1022_n 0.00453598f $X=4.94 $Y=1.96
+ $X2=0 $Y2=0
cc_609 N_A_702_21#_c_776_n N_A_506_47#_c_1022_n 0.00536992f $X=5.025 $Y=1.835
+ $X2=0 $Y2=0
cc_610 N_A_702_21#_c_781_n N_A_506_47#_c_1023_n 0.0115381f $X=4.94 $Y=1.96 $X2=0
+ $Y2=0
cc_611 N_A_702_21#_c_777_n N_A_506_47#_c_1014_n 0.0186016f $X=4.95 $Y=1.065
+ $X2=0 $Y2=0
cc_612 N_A_702_21#_c_781_n N_A_506_47#_c_1024_n 0.00131795f $X=4.94 $Y=1.96
+ $X2=0 $Y2=0
cc_613 N_A_702_21#_c_776_n N_A_506_47#_c_1024_n 0.00573895f $X=5.025 $Y=1.835
+ $X2=0 $Y2=0
cc_614 N_A_702_21#_c_781_n N_A_506_47#_c_1025_n 0.00770758f $X=4.94 $Y=1.96
+ $X2=0 $Y2=0
cc_615 N_A_702_21#_c_775_n N_A_506_47#_c_1015_n 0.00360556f $X=4.875 $Y=0.46
+ $X2=0 $Y2=0
cc_616 N_A_702_21#_c_779_n N_A_506_47#_c_1042_n 0.0022141f $X=3.61 $Y=1.99 $X2=0
+ $Y2=0
cc_617 N_A_702_21#_M1027_g N_A_506_47#_c_1046_n 0.00918626f $X=3.585 $Y=0.445
+ $X2=0 $Y2=0
cc_618 N_A_702_21#_M1027_g N_A_506_47#_c_1026_n 0.0103777f $X=3.585 $Y=0.445
+ $X2=0 $Y2=0
cc_619 N_A_702_21#_c_779_n N_A_506_47#_c_1026_n 0.00506348f $X=3.61 $Y=1.99
+ $X2=0 $Y2=0
cc_620 N_A_702_21#_c_783_n N_A_506_47#_c_1026_n 0.0370423f $X=3.695 $Y=1.74
+ $X2=0 $Y2=0
cc_621 N_A_702_21#_M1027_g N_A_506_47#_c_1017_n 0.0224362f $X=3.585 $Y=0.445
+ $X2=0 $Y2=0
cc_622 N_A_702_21#_c_780_n N_A_506_47#_c_1018_n 0.00979352f $X=4.34 $Y=1.96
+ $X2=0 $Y2=0
cc_623 N_A_702_21#_c_784_n N_A_506_47#_c_1018_n 0.00337624f $X=4.425 $Y=1.96
+ $X2=0 $Y2=0
cc_624 N_A_702_21#_M1027_g N_A_506_47#_c_1019_n 0.0100438f $X=3.585 $Y=0.445
+ $X2=0 $Y2=0
cc_625 N_A_702_21#_c_779_n N_A_506_47#_c_1019_n 0.00154583f $X=3.61 $Y=1.99
+ $X2=0 $Y2=0
cc_626 N_A_702_21#_c_783_n N_A_506_47#_c_1019_n 0.0205102f $X=3.695 $Y=1.74
+ $X2=0 $Y2=0
cc_627 N_A_702_21#_c_781_n N_A_506_47#_c_1020_n 0.00979462f $X=4.94 $Y=1.96
+ $X2=0 $Y2=0
cc_628 N_A_702_21#_c_776_n N_A_506_47#_c_1020_n 0.0232412f $X=5.025 $Y=1.835
+ $X2=0 $Y2=0
cc_629 N_A_702_21#_c_784_n N_A_506_47#_c_1020_n 0.00169427f $X=4.425 $Y=1.96
+ $X2=0 $Y2=0
cc_630 N_A_702_21#_c_781_n N_A_506_47#_c_1021_n 0.0029883f $X=4.94 $Y=1.96 $X2=0
+ $Y2=0
cc_631 N_A_702_21#_c_776_n N_A_506_47#_c_1021_n 0.0147229f $X=5.025 $Y=1.835
+ $X2=0 $Y2=0
cc_632 N_A_702_21#_c_777_n N_A_506_47#_c_1021_n 0.00411714f $X=4.95 $Y=1.065
+ $X2=0 $Y2=0
cc_633 N_A_702_21#_c_780_n N_VPWR_M1010_d 0.00142293f $X=4.34 $Y=1.96 $X2=0
+ $Y2=0
cc_634 N_A_702_21#_c_783_n N_VPWR_M1010_d 0.00165019f $X=3.695 $Y=1.74 $X2=0
+ $Y2=0
cc_635 N_A_702_21#_c_781_n N_VPWR_M1022_d 0.00182383f $X=4.94 $Y=1.96 $X2=0
+ $Y2=0
cc_636 N_A_702_21#_c_779_n N_VPWR_c_1545_n 0.0063127f $X=3.61 $Y=1.99 $X2=0
+ $Y2=0
cc_637 N_A_702_21#_c_783_n N_VPWR_c_1545_n 0.00186206f $X=3.695 $Y=1.74 $X2=0
+ $Y2=0
cc_638 N_A_702_21#_c_780_n N_VPWR_c_1546_n 0.00343021f $X=4.34 $Y=1.96 $X2=0
+ $Y2=0
cc_639 N_A_702_21#_c_858_p N_VPWR_c_1546_n 0.00733616f $X=4.425 $Y=2.21 $X2=0
+ $Y2=0
cc_640 N_A_702_21#_c_781_n N_VPWR_c_1546_n 0.00242429f $X=4.94 $Y=1.96 $X2=0
+ $Y2=0
cc_641 N_A_702_21#_c_781_n N_VPWR_c_1547_n 8.98216e-19 $X=4.94 $Y=1.96 $X2=0
+ $Y2=0
cc_642 N_A_702_21#_M1031_d N_VPWR_c_1532_n 0.00219951f $X=4.28 $Y=2.065 $X2=0
+ $Y2=0
cc_643 N_A_702_21#_c_779_n N_VPWR_c_1532_n 0.00765353f $X=3.61 $Y=1.99 $X2=0
+ $Y2=0
cc_644 N_A_702_21#_c_780_n N_VPWR_c_1532_n 0.00308649f $X=4.34 $Y=1.96 $X2=0
+ $Y2=0
cc_645 N_A_702_21#_c_858_p N_VPWR_c_1532_n 0.00288476f $X=4.425 $Y=2.21 $X2=0
+ $Y2=0
cc_646 N_A_702_21#_c_781_n N_VPWR_c_1532_n 0.00359426f $X=4.94 $Y=1.96 $X2=0
+ $Y2=0
cc_647 N_A_702_21#_c_783_n N_VPWR_c_1532_n 0.00197316f $X=3.695 $Y=1.74 $X2=0
+ $Y2=0
cc_648 N_A_702_21#_c_779_n N_VPWR_c_1554_n 0.00394773f $X=3.61 $Y=1.99 $X2=0
+ $Y2=0
cc_649 N_A_702_21#_c_780_n N_VPWR_c_1554_n 0.0102658f $X=4.34 $Y=1.96 $X2=0
+ $Y2=0
cc_650 N_A_702_21#_c_858_p N_VPWR_c_1554_n 0.00709892f $X=4.425 $Y=2.21 $X2=0
+ $Y2=0
cc_651 N_A_702_21#_c_783_n N_VPWR_c_1554_n 0.011698f $X=3.695 $Y=1.74 $X2=0
+ $Y2=0
cc_652 N_A_702_21#_c_858_p N_VPWR_c_1555_n 0.00895861f $X=4.425 $Y=2.21 $X2=0
+ $Y2=0
cc_653 N_A_702_21#_c_781_n N_VPWR_c_1555_n 0.0190229f $X=4.94 $Y=1.96 $X2=0
+ $Y2=0
cc_654 N_A_702_21#_c_775_n N_VGND_c_1886_n 0.0189546f $X=4.875 $Y=0.46 $X2=0
+ $Y2=0
cc_655 N_A_702_21#_M1027_g N_VGND_c_1893_n 0.0035977f $X=3.585 $Y=0.445 $X2=0
+ $Y2=0
cc_656 N_A_702_21#_c_775_n N_VGND_c_1894_n 0.00939086f $X=4.875 $Y=0.46 $X2=0
+ $Y2=0
cc_657 N_A_702_21#_c_777_n N_VGND_c_1894_n 0.00253654f $X=4.95 $Y=1.065 $X2=0
+ $Y2=0
cc_658 N_A_702_21#_M1030_d N_VGND_c_1898_n 0.00294605f $X=4.69 $Y=0.235 $X2=0
+ $Y2=0
cc_659 N_A_702_21#_M1027_g N_VGND_c_1898_n 0.00598452f $X=3.585 $Y=0.445 $X2=0
+ $Y2=0
cc_660 N_A_702_21#_c_775_n N_VGND_c_1898_n 0.00302049f $X=4.875 $Y=0.46 $X2=0
+ $Y2=0
cc_661 N_A_702_21#_c_777_n N_VGND_c_1898_n 0.00193724f $X=4.95 $Y=1.065 $X2=0
+ $Y2=0
cc_662 N_A_702_21#_M1027_g N_VGND_c_1901_n 0.00386585f $X=3.585 $Y=0.445 $X2=0
+ $Y2=0
cc_663 N_SET_B_M1026_g N_A_506_47#_c_1012_n 0.0271604f $X=4.255 $Y=0.445 $X2=0
+ $Y2=0
cc_664 N_SET_B_c_886_n N_A_506_47#_c_1013_n 0.00136929f $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_665 N_SET_B_c_889_n N_A_506_47#_c_1013_n 0.0148276f $X=4.19 $Y=0.98 $X2=0
+ $Y2=0
cc_666 N_SET_B_c_882_n N_A_506_47#_c_1022_n 0.0102791f $X=4.19 $Y=1.89 $X2=0
+ $Y2=0
cc_667 N_SET_B_c_894_n N_A_506_47#_c_1023_n 0.023055f $X=4.19 $Y=1.99 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_886_n N_A_506_47#_c_1014_n 0.00391536f $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_669 N_SET_B_c_886_n N_A_506_47#_c_1016_n 0.00446783f $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_670 N_SET_B_c_889_n N_A_506_47#_c_1016_n 0.0271604f $X=4.19 $Y=0.98 $X2=0
+ $Y2=0
cc_671 N_SET_B_c_892_n N_A_506_47#_c_1016_n 0.00309199f $X=4.365 $Y=0.85 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_882_n N_A_506_47#_c_1017_n 0.0010852f $X=4.19 $Y=1.89 $X2=0
+ $Y2=0
cc_673 N_SET_B_M1026_g N_A_506_47#_c_1017_n 0.00372275f $X=4.255 $Y=0.445 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_887_n N_A_506_47#_c_1017_n 8.97856e-19 $X=4.51 $Y=0.85 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_889_n N_A_506_47#_c_1017_n 0.00236863f $X=4.19 $Y=0.98 $X2=0
+ $Y2=0
cc_676 N_SET_B_c_892_n N_A_506_47#_c_1017_n 0.0262735f $X=4.365 $Y=0.85 $X2=0
+ $Y2=0
cc_677 N_SET_B_c_882_n N_A_506_47#_c_1018_n 0.0128663f $X=4.19 $Y=1.89 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_887_n N_A_506_47#_c_1018_n 2.49951e-19 $X=4.51 $Y=0.85 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_889_n N_A_506_47#_c_1018_n 0.00307815f $X=4.19 $Y=0.98 $X2=0
+ $Y2=0
cc_680 N_SET_B_c_892_n N_A_506_47#_c_1018_n 0.0362166f $X=4.365 $Y=0.85 $X2=0
+ $Y2=0
cc_681 N_SET_B_c_882_n N_A_506_47#_c_1020_n 0.00370432f $X=4.19 $Y=1.89 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_886_n N_A_506_47#_c_1020_n 0.00340769f $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_892_n N_A_506_47#_c_1020_n 0.00265163f $X=4.365 $Y=0.85 $X2=0
+ $Y2=0
cc_684 N_SET_B_c_882_n N_A_506_47#_c_1021_n 0.0207524f $X=4.19 $Y=1.89 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_886_n N_A_506_47#_c_1021_n 2.76699e-19 $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_895_n N_A_1288_261#_c_1172_n 0.00291216f $X=7.53 $Y=1.89 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_885_n N_A_1288_261#_c_1172_n 0.00482334f $X=7.52 $Y=1.535 $X2=0
+ $Y2=0
cc_688 N_SET_B_M1037_g N_A_1288_261#_M1034_g 0.0649482f $X=7.365 $Y=0.445 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_885_n N_A_1288_261#_M1034_g 0.0117891f $X=7.52 $Y=1.535 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_891_n N_A_1288_261#_M1034_g 0.00102512f $X=7.425 $Y=0.98 $X2=0
+ $Y2=0
cc_691 N_SET_B_c_888_n N_A_1288_261#_c_1174_n 0.00138899f $X=7.59 $Y=0.85 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_891_n N_A_1288_261#_c_1174_n 0.00815269f $X=7.425 $Y=0.98 $X2=0
+ $Y2=0
cc_693 N_SET_B_c_895_n N_A_1288_261#_c_1178_n 0.0117802f $X=7.53 $Y=1.89 $X2=0
+ $Y2=0
cc_694 N_SET_B_c_898_n N_A_1288_261#_c_1178_n 0.00902936f $X=7.52 $Y=1.685 $X2=0
+ $Y2=0
cc_695 N_SET_B_c_896_n N_A_1126_413#_c_1254_n 0.0129863f $X=7.53 $Y=1.99 $X2=0
+ $Y2=0
cc_696 N_SET_B_c_898_n N_A_1126_413#_c_1254_n 0.0153499f $X=7.52 $Y=1.685 $X2=0
+ $Y2=0
cc_697 N_SET_B_M1037_g N_A_1126_413#_M1028_g 0.0125249f $X=7.365 $Y=0.445 $X2=0
+ $Y2=0
cc_698 N_SET_B_c_890_n N_A_1126_413#_M1028_g 0.00745739f $X=7.425 $Y=0.98 $X2=0
+ $Y2=0
cc_699 N_SET_B_c_891_n N_A_1126_413#_M1028_g 0.00435751f $X=7.425 $Y=0.98 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_885_n N_A_1126_413#_c_1246_n 0.00474887f $X=7.52 $Y=1.535 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_898_n N_A_1126_413#_c_1246_n 0.00161253f $X=7.52 $Y=1.685 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_890_n N_A_1126_413#_c_1246_n 0.0224328f $X=7.425 $Y=0.98 $X2=0
+ $Y2=0
cc_703 N_SET_B_c_886_n N_A_1126_413#_c_1275_n 0.00677694f $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_704 N_SET_B_c_886_n N_A_1126_413#_c_1249_n 0.0109187f $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_886_n N_A_1126_413#_c_1250_n 0.00493969f $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_896_n N_A_1126_413#_c_1262_n 0.00481616f $X=7.53 $Y=1.99 $X2=0
+ $Y2=0
cc_707 N_SET_B_M1037_g N_A_1126_413#_c_1251_n 0.00278604f $X=7.365 $Y=0.445
+ $X2=0 $Y2=0
cc_708 N_SET_B_c_885_n N_A_1126_413#_c_1251_n 0.00159228f $X=7.52 $Y=1.535 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_886_n N_A_1126_413#_c_1251_n 0.0180658f $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_710 N_SET_B_c_888_n N_A_1126_413#_c_1251_n 4.39597e-19 $X=7.59 $Y=0.85 $X2=0
+ $Y2=0
cc_711 N_SET_B_c_890_n N_A_1126_413#_c_1251_n 0.00157366f $X=7.425 $Y=0.98 $X2=0
+ $Y2=0
cc_712 N_SET_B_c_891_n N_A_1126_413#_c_1251_n 0.0252903f $X=7.425 $Y=0.98 $X2=0
+ $Y2=0
cc_713 N_SET_B_c_885_n N_A_1126_413#_c_1252_n 0.0013797f $X=7.52 $Y=1.535 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_885_n N_A_1126_413#_c_1253_n 0.0123274f $X=7.52 $Y=1.535 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_898_n N_A_1126_413#_c_1253_n 5.27224e-19 $X=7.52 $Y=1.685 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_886_n N_A_1126_413#_c_1253_n 0.00766354f $X=7.445 $Y=0.85 $X2=0
+ $Y2=0
cc_717 N_SET_B_c_888_n N_A_1126_413#_c_1253_n 0.00171194f $X=7.59 $Y=0.85 $X2=0
+ $Y2=0
cc_718 N_SET_B_c_890_n N_A_1126_413#_c_1253_n 0.00347176f $X=7.425 $Y=0.98 $X2=0
+ $Y2=0
cc_719 N_SET_B_c_891_n N_A_1126_413#_c_1253_n 0.0344844f $X=7.425 $Y=0.98 $X2=0
+ $Y2=0
cc_720 N_SET_B_c_896_n N_VPWR_c_1536_n 0.010162f $X=7.53 $Y=1.99 $X2=0 $Y2=0
cc_721 N_SET_B_c_896_n N_VPWR_c_1540_n 0.00742396f $X=7.53 $Y=1.99 $X2=0 $Y2=0
cc_722 N_SET_B_c_894_n N_VPWR_c_1546_n 0.0048505f $X=4.19 $Y=1.99 $X2=0 $Y2=0
cc_723 N_SET_B_c_894_n N_VPWR_c_1532_n 0.00518398f $X=4.19 $Y=1.99 $X2=0 $Y2=0
cc_724 N_SET_B_c_896_n N_VPWR_c_1532_n 0.0147625f $X=7.53 $Y=1.99 $X2=0 $Y2=0
cc_725 N_SET_B_c_894_n N_VPWR_c_1554_n 0.0103343f $X=4.19 $Y=1.99 $X2=0 $Y2=0
cc_726 N_SET_B_c_894_n N_VPWR_c_1555_n 7.74208e-19 $X=4.19 $Y=1.99 $X2=0 $Y2=0
cc_727 N_SET_B_c_896_n N_VPWR_c_1556_n 0.00497911f $X=7.53 $Y=1.99 $X2=0 $Y2=0
cc_728 N_SET_B_c_891_n N_VGND_M1037_d 0.00117915f $X=7.425 $Y=0.98 $X2=0 $Y2=0
cc_729 N_SET_B_c_886_n N_VGND_c_1886_n 0.00733061f $X=7.445 $Y=0.85 $X2=0 $Y2=0
cc_730 N_SET_B_c_892_n N_VGND_c_1894_n 0.00213925f $X=4.365 $Y=0.85 $X2=0 $Y2=0
cc_731 N_SET_B_M1037_g N_VGND_c_1898_n 0.00141612f $X=7.365 $Y=0.445 $X2=0 $Y2=0
cc_732 N_SET_B_c_886_n N_VGND_c_1898_n 0.136054f $X=7.445 $Y=0.85 $X2=0 $Y2=0
cc_733 N_SET_B_c_887_n N_VGND_c_1898_n 0.0154019f $X=4.51 $Y=0.85 $X2=0 $Y2=0
cc_734 N_SET_B_c_888_n N_VGND_c_1898_n 0.0131415f $X=7.59 $Y=0.85 $X2=0 $Y2=0
cc_735 N_SET_B_c_891_n N_VGND_c_1898_n 0.0013061f $X=7.425 $Y=0.98 $X2=0 $Y2=0
cc_736 N_SET_B_c_892_n N_VGND_c_1898_n 0.00237941f $X=4.365 $Y=0.85 $X2=0 $Y2=0
cc_737 N_SET_B_M1026_g N_VGND_c_1901_n 0.013844f $X=4.255 $Y=0.445 $X2=0 $Y2=0
cc_738 N_SET_B_c_887_n N_VGND_c_1901_n 0.00153265f $X=4.51 $Y=0.85 $X2=0 $Y2=0
cc_739 N_SET_B_c_889_n N_VGND_c_1901_n 0.00134756f $X=4.19 $Y=0.98 $X2=0 $Y2=0
cc_740 N_SET_B_c_892_n N_VGND_c_1901_n 0.0251483f $X=4.365 $Y=0.85 $X2=0 $Y2=0
cc_741 N_SET_B_M1037_g N_VGND_c_1903_n 8.70124e-19 $X=7.365 $Y=0.445 $X2=0 $Y2=0
cc_742 N_SET_B_c_891_n N_VGND_c_1903_n 8.77612e-19 $X=7.425 $Y=0.98 $X2=0 $Y2=0
cc_743 N_SET_B_M1037_g N_VGND_c_1904_n 0.0226474f $X=7.365 $Y=0.445 $X2=0 $Y2=0
cc_744 N_SET_B_c_886_n N_VGND_c_1904_n 5.4944e-19 $X=7.445 $Y=0.85 $X2=0 $Y2=0
cc_745 N_SET_B_c_888_n N_VGND_c_1904_n 0.00154076f $X=7.59 $Y=0.85 $X2=0 $Y2=0
cc_746 N_SET_B_c_890_n N_VGND_c_1904_n 9.26709e-19 $X=7.425 $Y=0.98 $X2=0 $Y2=0
cc_747 N_SET_B_c_891_n N_VGND_c_1904_n 0.0312846f $X=7.425 $Y=0.98 $X2=0 $Y2=0
cc_748 N_A_506_47#_c_1025_n N_A_1126_413#_c_1267_n 9.38727e-19 $X=5.13 $Y=1.99
+ $X2=0 $Y2=0
cc_749 N_A_506_47#_c_1042_n N_VPWR_c_1545_n 0.0425549f $X=3.27 $Y=2.335 $X2=0
+ $Y2=0
cc_750 N_A_506_47#_c_1023_n N_VPWR_c_1546_n 0.00315013f $X=4.66 $Y=1.99 $X2=0
+ $Y2=0
cc_751 N_A_506_47#_c_1025_n N_VPWR_c_1547_n 0.00591633f $X=5.13 $Y=1.99 $X2=0
+ $Y2=0
cc_752 N_A_506_47#_M1033_d N_VPWR_c_1532_n 0.00192288f $X=2.58 $Y=2.065 $X2=0
+ $Y2=0
cc_753 N_A_506_47#_c_1023_n N_VPWR_c_1532_n 0.00358098f $X=4.66 $Y=1.99 $X2=0
+ $Y2=0
cc_754 N_A_506_47#_c_1025_n N_VPWR_c_1532_n 0.00554886f $X=5.13 $Y=1.99 $X2=0
+ $Y2=0
cc_755 N_A_506_47#_c_1042_n N_VPWR_c_1532_n 0.0149757f $X=3.27 $Y=2.335 $X2=0
+ $Y2=0
cc_756 N_A_506_47#_c_1023_n N_VPWR_c_1554_n 6.83681e-19 $X=4.66 $Y=1.99 $X2=0
+ $Y2=0
cc_757 N_A_506_47#_c_1023_n N_VPWR_c_1555_n 0.0101587f $X=4.66 $Y=1.99 $X2=0
+ $Y2=0
cc_758 N_A_506_47#_c_1025_n N_VPWR_c_1555_n 0.00901789f $X=5.13 $Y=1.99 $X2=0
+ $Y2=0
cc_759 N_A_506_47#_c_1046_n N_A_409_329#_c_1737_n 0.00758237f $X=3.52 $Y=0.365
+ $X2=0 $Y2=0
cc_760 N_A_506_47#_c_1042_n N_A_409_329#_c_1738_n 0.0102747f $X=3.27 $Y=2.335
+ $X2=0 $Y2=0
cc_761 N_A_506_47#_c_1042_n A_610_413# 0.00898626f $X=3.27 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_762 N_A_506_47#_c_1026_n A_610_413# 0.0058128f $X=3.355 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_763 N_A_506_47#_c_1046_n N_VGND_M1027_d 0.00216229f $X=3.52 $Y=0.365 $X2=0
+ $Y2=0
cc_764 N_A_506_47#_c_1017_n N_VGND_M1027_d 0.00251036f $X=3.63 $Y=1.23 $X2=0
+ $Y2=0
cc_765 N_A_506_47#_c_1012_n N_VGND_c_1886_n 0.00394489f $X=4.615 $Y=0.735 $X2=0
+ $Y2=0
cc_766 N_A_506_47#_c_1014_n N_VGND_c_1886_n 0.00913201f $X=5.63 $Y=0.825 $X2=0
+ $Y2=0
cc_767 N_A_506_47#_c_1015_n N_VGND_c_1886_n 0.00901822f $X=5.705 $Y=0.735 $X2=0
+ $Y2=0
cc_768 N_A_506_47#_c_1046_n N_VGND_c_1893_n 0.0613943f $X=3.52 $Y=0.365 $X2=0
+ $Y2=0
cc_769 N_A_506_47#_c_1012_n N_VGND_c_1894_n 0.00585385f $X=4.615 $Y=0.735 $X2=0
+ $Y2=0
cc_770 N_A_506_47#_c_1014_n N_VGND_c_1894_n 0.00163052f $X=5.63 $Y=0.825 $X2=0
+ $Y2=0
cc_771 N_A_506_47#_M1003_d N_VGND_c_1898_n 0.0035796f $X=2.53 $Y=0.235 $X2=0
+ $Y2=0
cc_772 N_A_506_47#_c_1012_n N_VGND_c_1898_n 0.00768024f $X=4.615 $Y=0.735 $X2=0
+ $Y2=0
cc_773 N_A_506_47#_c_1014_n N_VGND_c_1898_n 5.56212e-19 $X=5.63 $Y=0.825 $X2=0
+ $Y2=0
cc_774 N_A_506_47#_c_1015_n N_VGND_c_1898_n 0.00700878f $X=5.705 $Y=0.735 $X2=0
+ $Y2=0
cc_775 N_A_506_47#_c_1046_n N_VGND_c_1898_n 0.024944f $X=3.52 $Y=0.365 $X2=0
+ $Y2=0
cc_776 N_A_506_47#_c_1012_n N_VGND_c_1901_n 0.00304708f $X=4.615 $Y=0.735 $X2=0
+ $Y2=0
cc_777 N_A_506_47#_c_1046_n N_VGND_c_1901_n 0.0174415f $X=3.52 $Y=0.365 $X2=0
+ $Y2=0
cc_778 N_A_506_47#_c_1017_n N_VGND_c_1901_n 0.00475551f $X=3.63 $Y=1.23 $X2=0
+ $Y2=0
cc_779 N_A_506_47#_c_1015_n N_VGND_c_1903_n 0.00437852f $X=5.705 $Y=0.735 $X2=0
+ $Y2=0
cc_780 N_A_506_47#_c_1046_n A_636_47# 0.00625113f $X=3.52 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_781 N_A_1288_261#_c_1178_n N_A_1126_413#_c_1254_n 0.0156189f $X=8.21 $Y=1.67
+ $X2=0 $Y2=0
cc_782 N_A_1288_261#_c_1174_n N_A_1126_413#_M1028_g 0.0107516f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_783 N_A_1288_261#_c_1174_n N_A_1126_413#_c_1245_n 0.0267728f $X=8.445
+ $Y=1.575 $X2=0 $Y2=0
cc_784 N_A_1288_261#_c_1175_n N_A_1126_413#_c_1245_n 0.00339526f $X=8.445
+ $Y=0.515 $X2=0 $Y2=0
cc_785 N_A_1288_261#_c_1178_n N_A_1126_413#_c_1245_n 0.0071742f $X=8.21 $Y=1.67
+ $X2=0 $Y2=0
cc_786 N_A_1288_261#_c_1179_n N_A_1126_413#_c_1245_n 0.00109088f $X=8.445
+ $Y=1.67 $X2=0 $Y2=0
cc_787 N_A_1288_261#_c_1174_n N_A_1126_413#_c_1246_n 0.00519959f $X=8.445
+ $Y=1.575 $X2=0 $Y2=0
cc_788 N_A_1288_261#_c_1178_n N_A_1126_413#_c_1246_n 0.00382811f $X=8.21 $Y=1.67
+ $X2=0 $Y2=0
cc_789 N_A_1288_261#_c_1174_n N_A_1126_413#_c_1257_n 6.49825e-19 $X=8.445
+ $Y=1.575 $X2=0 $Y2=0
cc_790 N_A_1288_261#_c_1179_n N_A_1126_413#_c_1257_n 9.05513e-19 $X=8.445
+ $Y=1.67 $X2=0 $Y2=0
cc_791 N_A_1288_261#_c_1205_p N_A_1126_413#_c_1258_n 0.00120203f $X=8.295
+ $Y=1.87 $X2=0 $Y2=0
cc_792 N_A_1288_261#_c_1174_n N_A_1126_413#_M1006_g 7.06846e-19 $X=8.445
+ $Y=1.575 $X2=0 $Y2=0
cc_793 N_A_1288_261#_c_1172_n N_A_1126_413#_c_1260_n 0.00848051f $X=6.54 $Y=1.99
+ $X2=0 $Y2=0
cc_794 N_A_1288_261#_c_1178_n N_A_1126_413#_c_1260_n 0.0135877f $X=8.21 $Y=1.67
+ $X2=0 $Y2=0
cc_795 N_A_1288_261#_M1034_g N_A_1126_413#_c_1275_n 0.00578747f $X=7.005
+ $Y=0.445 $X2=0 $Y2=0
cc_796 N_A_1288_261#_c_1172_n N_A_1126_413#_c_1249_n 0.0153888f $X=6.54 $Y=1.99
+ $X2=0 $Y2=0
cc_797 N_A_1288_261#_c_1178_n N_A_1126_413#_c_1249_n 0.0315564f $X=8.21 $Y=1.67
+ $X2=0 $Y2=0
cc_798 N_A_1288_261#_c_1172_n N_A_1126_413#_c_1262_n 0.0185082f $X=6.54 $Y=1.99
+ $X2=0 $Y2=0
cc_799 N_A_1288_261#_c_1178_n N_A_1126_413#_c_1262_n 0.0688065f $X=8.21 $Y=1.67
+ $X2=0 $Y2=0
cc_800 N_A_1288_261#_M1034_g N_A_1126_413#_c_1251_n 0.01482f $X=7.005 $Y=0.445
+ $X2=0 $Y2=0
cc_801 N_A_1288_261#_c_1172_n N_A_1126_413#_c_1263_n 0.00296227f $X=6.54 $Y=1.99
+ $X2=0 $Y2=0
cc_802 N_A_1288_261#_c_1172_n N_A_1126_413#_c_1264_n 0.0047082f $X=6.54 $Y=1.99
+ $X2=0 $Y2=0
cc_803 N_A_1288_261#_c_1172_n N_A_1126_413#_c_1345_n 0.0041236f $X=6.54 $Y=1.99
+ $X2=0 $Y2=0
cc_804 N_A_1288_261#_M1034_g N_A_1126_413#_c_1345_n 0.00355592f $X=7.005
+ $Y=0.445 $X2=0 $Y2=0
cc_805 N_A_1288_261#_c_1178_n N_A_1126_413#_c_1345_n 0.0136304f $X=8.21 $Y=1.67
+ $X2=0 $Y2=0
cc_806 N_A_1288_261#_c_1174_n N_A_1126_413#_c_1252_n 0.0174138f $X=8.445
+ $Y=1.575 $X2=0 $Y2=0
cc_807 N_A_1288_261#_c_1178_n N_A_1126_413#_c_1253_n 0.0777752f $X=8.21 $Y=1.67
+ $X2=0 $Y2=0
cc_808 N_A_1288_261#_c_1174_n N_A_1738_47#_c_1412_n 0.0283443f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_809 N_A_1288_261#_c_1175_n N_A_1738_47#_c_1412_n 0.0254199f $X=8.445 $Y=0.515
+ $X2=0 $Y2=0
cc_810 N_A_1288_261#_c_1205_p N_A_1738_47#_c_1421_n 0.0257384f $X=8.295 $Y=1.87
+ $X2=0 $Y2=0
cc_811 N_A_1288_261#_c_1205_p N_A_1738_47#_c_1422_n 0.00670345f $X=8.295 $Y=1.87
+ $X2=0 $Y2=0
cc_812 N_A_1288_261#_c_1174_n N_A_1738_47#_c_1422_n 0.021487f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_813 N_A_1288_261#_c_1179_n N_A_1738_47#_c_1422_n 0.0155746f $X=8.445 $Y=1.67
+ $X2=0 $Y2=0
cc_814 N_A_1288_261#_c_1174_n N_A_1738_47#_c_1414_n 0.0165785f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_815 N_A_1288_261#_c_1178_n N_VPWR_M1000_d 0.00253127f $X=8.21 $Y=1.67 $X2=0
+ $Y2=0
cc_816 N_A_1288_261#_c_1205_p N_VPWR_c_1536_n 0.0317496f $X=8.295 $Y=1.87 $X2=0
+ $Y2=0
cc_817 N_A_1288_261#_c_1178_n N_VPWR_c_1536_n 0.0191712f $X=8.21 $Y=1.67 $X2=0
+ $Y2=0
cc_818 N_A_1288_261#_c_1172_n N_VPWR_c_1547_n 5.99585e-19 $X=6.54 $Y=1.99 $X2=0
+ $Y2=0
cc_819 N_A_1288_261#_c_1205_p N_VPWR_c_1548_n 0.00739842f $X=8.295 $Y=1.87 $X2=0
+ $Y2=0
cc_820 N_A_1288_261#_M1023_d N_VPWR_c_1532_n 0.00577926f $X=8.15 $Y=1.645 $X2=0
+ $Y2=0
cc_821 N_A_1288_261#_c_1172_n N_VPWR_c_1532_n 0.00125542f $X=6.54 $Y=1.99 $X2=0
+ $Y2=0
cc_822 N_A_1288_261#_c_1205_p N_VPWR_c_1532_n 0.00614354f $X=8.295 $Y=1.87 $X2=0
+ $Y2=0
cc_823 N_A_1288_261#_c_1172_n N_VPWR_c_1556_n 0.0171834f $X=6.54 $Y=1.99 $X2=0
+ $Y2=0
cc_824 N_A_1288_261#_c_1175_n N_VGND_c_1890_n 0.0140151f $X=8.445 $Y=0.515 $X2=0
+ $Y2=0
cc_825 N_A_1288_261#_M1028_d N_VGND_c_1898_n 0.00391384f $X=8.16 $Y=0.235 $X2=0
+ $Y2=0
cc_826 N_A_1288_261#_M1034_g N_VGND_c_1898_n 0.00495706f $X=7.005 $Y=0.445 $X2=0
+ $Y2=0
cc_827 N_A_1288_261#_c_1175_n N_VGND_c_1898_n 0.0121445f $X=8.445 $Y=0.515 $X2=0
+ $Y2=0
cc_828 N_A_1288_261#_M1034_g N_VGND_c_1903_n 0.00367922f $X=7.005 $Y=0.445 $X2=0
+ $Y2=0
cc_829 N_A_1288_261#_M1034_g N_VGND_c_1904_n 0.00217209f $X=7.005 $Y=0.445 $X2=0
+ $Y2=0
cc_830 N_A_1126_413#_M1006_g N_A_1738_47#_M1001_g 0.0189791f $X=9.075 $Y=0.445
+ $X2=0 $Y2=0
cc_831 N_A_1126_413#_c_1258_n N_A_1738_47#_c_1416_n 0.0151315f $X=9.05 $Y=1.77
+ $X2=0 $Y2=0
cc_832 N_A_1126_413#_c_1248_n N_A_1738_47#_c_1416_n 0.0129816f $X=9.05 $Y=1.26
+ $X2=0 $Y2=0
cc_833 N_A_1126_413#_M1006_g N_A_1738_47#_c_1412_n 0.0168506f $X=9.075 $Y=0.445
+ $X2=0 $Y2=0
cc_834 N_A_1126_413#_M1006_g N_A_1738_47#_c_1413_n 0.00861898f $X=9.075 $Y=0.445
+ $X2=0 $Y2=0
cc_835 N_A_1126_413#_c_1248_n N_A_1738_47#_c_1413_n 0.0129394f $X=9.05 $Y=1.26
+ $X2=0 $Y2=0
cc_836 N_A_1126_413#_c_1254_n N_A_1738_47#_c_1421_n 0.00144689f $X=8.06 $Y=1.57
+ $X2=0 $Y2=0
cc_837 N_A_1126_413#_c_1245_n N_A_1738_47#_c_1421_n 0.00240579f $X=8.95 $Y=1.26
+ $X2=0 $Y2=0
cc_838 N_A_1126_413#_c_1258_n N_A_1738_47#_c_1421_n 0.00606783f $X=9.05 $Y=1.77
+ $X2=0 $Y2=0
cc_839 N_A_1126_413#_c_1254_n N_A_1738_47#_c_1422_n 4.30877e-19 $X=8.06 $Y=1.57
+ $X2=0 $Y2=0
cc_840 N_A_1126_413#_c_1245_n N_A_1738_47#_c_1422_n 0.0105805f $X=8.95 $Y=1.26
+ $X2=0 $Y2=0
cc_841 N_A_1126_413#_c_1257_n N_A_1738_47#_c_1422_n 0.00939457f $X=9.05 $Y=1.67
+ $X2=0 $Y2=0
cc_842 N_A_1126_413#_c_1258_n N_A_1738_47#_c_1422_n 0.00760246f $X=9.05 $Y=1.77
+ $X2=0 $Y2=0
cc_843 N_A_1126_413#_c_1248_n N_A_1738_47#_c_1422_n 0.00295914f $X=9.05 $Y=1.26
+ $X2=0 $Y2=0
cc_844 N_A_1126_413#_c_1245_n N_A_1738_47#_c_1414_n 0.0108298f $X=8.95 $Y=1.26
+ $X2=0 $Y2=0
cc_845 N_A_1126_413#_c_1248_n N_A_1738_47#_c_1414_n 5.08488e-19 $X=9.05 $Y=1.26
+ $X2=0 $Y2=0
cc_846 N_A_1126_413#_c_1248_n N_A_1738_47#_c_1415_n 0.0189791f $X=9.05 $Y=1.26
+ $X2=0 $Y2=0
cc_847 N_A_1126_413#_c_1262_n N_VPWR_M1011_d 0.00226245f $X=7.14 $Y=2 $X2=0
+ $Y2=0
cc_848 N_A_1126_413#_c_1254_n N_VPWR_c_1536_n 0.0190345f $X=8.06 $Y=1.57 $X2=0
+ $Y2=0
cc_849 N_A_1126_413#_c_1262_n N_VPWR_c_1536_n 0.0075203f $X=7.14 $Y=2 $X2=0
+ $Y2=0
cc_850 N_A_1126_413#_c_1263_n N_VPWR_c_1536_n 0.0139175f $X=7.295 $Y=2.21 $X2=0
+ $Y2=0
cc_851 N_A_1126_413#_c_1258_n N_VPWR_c_1537_n 0.00650857f $X=9.05 $Y=1.77 $X2=0
+ $Y2=0
cc_852 N_A_1126_413#_c_1262_n N_VPWR_c_1540_n 0.0036467f $X=7.14 $Y=2 $X2=0
+ $Y2=0
cc_853 N_A_1126_413#_c_1263_n N_VPWR_c_1540_n 0.0103119f $X=7.295 $Y=2.21 $X2=0
+ $Y2=0
cc_854 N_A_1126_413#_c_1267_n N_VPWR_c_1547_n 0.0224673f $X=6.07 $Y=2.29 $X2=0
+ $Y2=0
cc_855 N_A_1126_413#_c_1262_n N_VPWR_c_1547_n 0.00268786f $X=7.14 $Y=2 $X2=0
+ $Y2=0
cc_856 N_A_1126_413#_c_1264_n N_VPWR_c_1547_n 0.00983468f $X=6.18 $Y=2 $X2=0
+ $Y2=0
cc_857 N_A_1126_413#_c_1254_n N_VPWR_c_1548_n 0.00427505f $X=8.06 $Y=1.57 $X2=0
+ $Y2=0
cc_858 N_A_1126_413#_c_1258_n N_VPWR_c_1548_n 0.00674661f $X=9.05 $Y=1.77 $X2=0
+ $Y2=0
cc_859 N_A_1126_413#_M1035_d N_VPWR_c_1532_n 0.00289852f $X=5.63 $Y=2.065 $X2=0
+ $Y2=0
cc_860 N_A_1126_413#_M1000_s N_VPWR_c_1532_n 0.00413719f $X=7.17 $Y=2.065 $X2=0
+ $Y2=0
cc_861 N_A_1126_413#_c_1254_n N_VPWR_c_1532_n 0.00873932f $X=8.06 $Y=1.57 $X2=0
+ $Y2=0
cc_862 N_A_1126_413#_c_1258_n N_VPWR_c_1532_n 0.0133366f $X=9.05 $Y=1.77 $X2=0
+ $Y2=0
cc_863 N_A_1126_413#_c_1267_n N_VPWR_c_1532_n 0.0108989f $X=6.07 $Y=2.29 $X2=0
+ $Y2=0
cc_864 N_A_1126_413#_c_1262_n N_VPWR_c_1532_n 0.0127539f $X=7.14 $Y=2 $X2=0
+ $Y2=0
cc_865 N_A_1126_413#_c_1263_n N_VPWR_c_1532_n 0.0086238f $X=7.295 $Y=2.21 $X2=0
+ $Y2=0
cc_866 N_A_1126_413#_c_1264_n N_VPWR_c_1532_n 0.00748335f $X=6.18 $Y=2 $X2=0
+ $Y2=0
cc_867 N_A_1126_413#_c_1267_n N_VPWR_c_1555_n 0.00518401f $X=6.07 $Y=2.29 $X2=0
+ $Y2=0
cc_868 N_A_1126_413#_c_1262_n N_VPWR_c_1556_n 0.030653f $X=7.14 $Y=2 $X2=0 $Y2=0
cc_869 N_A_1126_413#_c_1263_n N_VPWR_c_1556_n 0.00894969f $X=7.295 $Y=2.21 $X2=0
+ $Y2=0
cc_870 N_A_1126_413#_c_1264_n N_VPWR_c_1556_n 0.0118413f $X=6.18 $Y=2 $X2=0
+ $Y2=0
cc_871 N_A_1126_413#_c_1262_n A_1244_413# 0.00184128f $X=7.14 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_872 N_A_1126_413#_c_1264_n A_1244_413# 0.00358395f $X=6.18 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_873 N_A_1126_413#_c_1275_n N_VGND_c_1886_n 0.00548171f $X=6.92 $Y=0.39 $X2=0
+ $Y2=0
cc_874 N_A_1126_413#_M1006_g N_VGND_c_1887_n 0.00297294f $X=9.075 $Y=0.445 $X2=0
+ $Y2=0
cc_875 N_A_1126_413#_M1028_g N_VGND_c_1890_n 0.00505556f $X=8.085 $Y=0.505 $X2=0
+ $Y2=0
cc_876 N_A_1126_413#_M1006_g N_VGND_c_1890_n 0.00585385f $X=9.075 $Y=0.445 $X2=0
+ $Y2=0
cc_877 N_A_1126_413#_M1012_d N_VGND_c_1898_n 0.00252861f $X=6.19 $Y=0.235 $X2=0
+ $Y2=0
cc_878 N_A_1126_413#_M1028_g N_VGND_c_1898_n 0.00991048f $X=8.085 $Y=0.505 $X2=0
+ $Y2=0
cc_879 N_A_1126_413#_M1006_g N_VGND_c_1898_n 0.0121216f $X=9.075 $Y=0.445 $X2=0
+ $Y2=0
cc_880 N_A_1126_413#_c_1275_n N_VGND_c_1898_n 0.0143646f $X=6.92 $Y=0.39 $X2=0
+ $Y2=0
cc_881 N_A_1126_413#_c_1275_n N_VGND_c_1903_n 0.0385814f $X=6.92 $Y=0.39 $X2=0
+ $Y2=0
cc_882 N_A_1126_413#_M1028_g N_VGND_c_1904_n 0.019957f $X=8.085 $Y=0.505 $X2=0
+ $Y2=0
cc_883 N_A_1126_413#_c_1246_n N_VGND_c_1904_n 0.00340309f $X=8.16 $Y=1.26 $X2=0
+ $Y2=0
cc_884 N_A_1126_413#_c_1252_n N_VGND_c_1904_n 0.00614106f $X=7.955 $Y=1.26 $X2=0
+ $Y2=0
cc_885 N_A_1126_413#_c_1253_n N_VGND_c_1904_n 2.87913e-19 $X=7.79 $Y=1.29 $X2=0
+ $Y2=0
cc_886 N_A_1126_413#_c_1275_n A_1344_47# 0.00244121f $X=6.92 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_887 N_A_1738_47#_c_1421_n N_VPWR_c_1536_n 0.00150527f $X=8.815 $Y=2 $X2=0
+ $Y2=0
cc_888 N_A_1738_47#_c_1416_n N_VPWR_c_1537_n 0.0154386f $X=9.575 $Y=1.41 $X2=0
+ $Y2=0
cc_889 N_A_1738_47#_c_1417_n N_VPWR_c_1537_n 7.64428e-19 $X=10.045 $Y=1.41 $X2=0
+ $Y2=0
cc_890 N_A_1738_47#_c_1413_n N_VPWR_c_1537_n 0.0111295f $X=11.2 $Y=1.16 $X2=0
+ $Y2=0
cc_891 N_A_1738_47#_c_1422_n N_VPWR_c_1537_n 0.0188541f $X=8.815 $Y=1.915 $X2=0
+ $Y2=0
cc_892 N_A_1738_47#_c_1417_n N_VPWR_c_1538_n 0.00293525f $X=10.045 $Y=1.41 $X2=0
+ $Y2=0
cc_893 N_A_1738_47#_c_1418_n N_VPWR_c_1538_n 0.00313746f $X=10.515 $Y=1.41 $X2=0
+ $Y2=0
cc_894 N_A_1738_47#_c_1418_n N_VPWR_c_1539_n 6.95418e-19 $X=10.515 $Y=1.41 $X2=0
+ $Y2=0
cc_895 N_A_1738_47#_c_1419_n N_VPWR_c_1539_n 0.0123478f $X=10.985 $Y=1.41 $X2=0
+ $Y2=0
cc_896 N_A_1738_47#_c_1420_n N_VPWR_c_1539_n 0.0176915f $X=11.455 $Y=1.41 $X2=0
+ $Y2=0
cc_897 N_A_1738_47#_c_1416_n N_VPWR_c_1542_n 0.0046653f $X=9.575 $Y=1.41 $X2=0
+ $Y2=0
cc_898 N_A_1738_47#_c_1417_n N_VPWR_c_1542_n 0.00643255f $X=10.045 $Y=1.41 $X2=0
+ $Y2=0
cc_899 N_A_1738_47#_c_1421_n N_VPWR_c_1548_n 0.0166846f $X=8.815 $Y=2 $X2=0
+ $Y2=0
cc_900 N_A_1738_47#_c_1418_n N_VPWR_c_1549_n 0.00702461f $X=10.515 $Y=1.41 $X2=0
+ $Y2=0
cc_901 N_A_1738_47#_c_1419_n N_VPWR_c_1549_n 0.00622633f $X=10.985 $Y=1.41 $X2=0
+ $Y2=0
cc_902 N_A_1738_47#_c_1420_n N_VPWR_c_1550_n 0.00427505f $X=11.455 $Y=1.41 $X2=0
+ $Y2=0
cc_903 N_A_1738_47#_M1009_s N_VPWR_c_1532_n 0.00219849f $X=8.69 $Y=1.845 $X2=0
+ $Y2=0
cc_904 N_A_1738_47#_c_1416_n N_VPWR_c_1532_n 0.00802193f $X=9.575 $Y=1.41 $X2=0
+ $Y2=0
cc_905 N_A_1738_47#_c_1417_n N_VPWR_c_1532_n 0.0111474f $X=10.045 $Y=1.41 $X2=0
+ $Y2=0
cc_906 N_A_1738_47#_c_1418_n N_VPWR_c_1532_n 0.0125271f $X=10.515 $Y=1.41 $X2=0
+ $Y2=0
cc_907 N_A_1738_47#_c_1419_n N_VPWR_c_1532_n 0.010479f $X=10.985 $Y=1.41 $X2=0
+ $Y2=0
cc_908 N_A_1738_47#_c_1420_n N_VPWR_c_1532_n 0.00836369f $X=11.455 $Y=1.41 $X2=0
+ $Y2=0
cc_909 N_A_1738_47#_c_1421_n N_VPWR_c_1532_n 0.0121973f $X=8.815 $Y=2 $X2=0
+ $Y2=0
cc_910 N_A_1738_47#_c_1417_n N_Q_c_1798_n 0.0124576f $X=10.045 $Y=1.41 $X2=0
+ $Y2=0
cc_911 N_A_1738_47#_c_1418_n N_Q_c_1798_n 0.0173289f $X=10.515 $Y=1.41 $X2=0
+ $Y2=0
cc_912 N_A_1738_47#_c_1413_n N_Q_c_1798_n 0.042778f $X=11.2 $Y=1.16 $X2=0 $Y2=0
cc_913 N_A_1738_47#_c_1415_n N_Q_c_1798_n 0.00866575f $X=11.455 $Y=1.217 $X2=0
+ $Y2=0
cc_914 N_A_1738_47#_c_1416_n N_Q_c_1799_n 0.00533245f $X=9.575 $Y=1.41 $X2=0
+ $Y2=0
cc_915 N_A_1738_47#_c_1417_n N_Q_c_1799_n 0.00271972f $X=10.045 $Y=1.41 $X2=0
+ $Y2=0
cc_916 N_A_1738_47#_c_1413_n N_Q_c_1799_n 0.0198063f $X=11.2 $Y=1.16 $X2=0 $Y2=0
cc_917 N_A_1738_47#_c_1415_n N_Q_c_1799_n 0.00573619f $X=11.455 $Y=1.217 $X2=0
+ $Y2=0
cc_918 N_A_1738_47#_M1015_g N_Q_c_1813_n 0.00600753f $X=10.02 $Y=0.56 $X2=0
+ $Y2=0
cc_919 N_A_1738_47#_M1016_g N_Q_c_1813_n 0.0101899f $X=10.49 $Y=0.56 $X2=0 $Y2=0
cc_920 N_A_1738_47#_c_1413_n N_Q_c_1813_n 0.0389951f $X=11.2 $Y=1.16 $X2=0 $Y2=0
cc_921 N_A_1738_47#_c_1415_n N_Q_c_1813_n 0.00334116f $X=11.455 $Y=1.217 $X2=0
+ $Y2=0
cc_922 N_A_1738_47#_M1001_g N_Q_c_1794_n 0.00469739f $X=9.55 $Y=0.56 $X2=0 $Y2=0
cc_923 N_A_1738_47#_M1015_g N_Q_c_1794_n 0.0030035f $X=10.02 $Y=0.56 $X2=0 $Y2=0
cc_924 N_A_1738_47#_c_1413_n N_Q_c_1794_n 0.0211685f $X=11.2 $Y=1.16 $X2=0 $Y2=0
cc_925 N_A_1738_47#_c_1415_n N_Q_c_1794_n 0.00300434f $X=11.455 $Y=1.217 $X2=0
+ $Y2=0
cc_926 N_A_1738_47#_M1016_g N_Q_c_1821_n 0.00276487f $X=10.49 $Y=0.56 $X2=0
+ $Y2=0
cc_927 N_A_1738_47#_c_1418_n N_Q_c_1822_n 0.00447353f $X=10.515 $Y=1.41 $X2=0
+ $Y2=0
cc_928 N_A_1738_47#_c_1419_n N_Q_c_1822_n 0.0060715f $X=10.985 $Y=1.41 $X2=0
+ $Y2=0
cc_929 N_A_1738_47#_M1018_g N_Q_c_1824_n 0.0114403f $X=10.96 $Y=0.56 $X2=0 $Y2=0
cc_930 N_A_1738_47#_M1039_g N_Q_c_1824_n 0.0129206f $X=11.48 $Y=0.56 $X2=0 $Y2=0
cc_931 N_A_1738_47#_c_1413_n N_Q_c_1824_n 0.0368992f $X=11.2 $Y=1.16 $X2=0 $Y2=0
cc_932 N_A_1738_47#_c_1415_n N_Q_c_1824_n 0.00423509f $X=11.455 $Y=1.217 $X2=0
+ $Y2=0
cc_933 N_A_1738_47#_c_1419_n N_Q_c_1800_n 0.0167909f $X=10.985 $Y=1.41 $X2=0
+ $Y2=0
cc_934 N_A_1738_47#_c_1420_n N_Q_c_1800_n 0.0177208f $X=11.455 $Y=1.41 $X2=0
+ $Y2=0
cc_935 N_A_1738_47#_c_1413_n N_Q_c_1800_n 0.0387812f $X=11.2 $Y=1.16 $X2=0 $Y2=0
cc_936 N_A_1738_47#_c_1415_n N_Q_c_1800_n 0.0088244f $X=11.455 $Y=1.217 $X2=0
+ $Y2=0
cc_937 N_A_1738_47#_c_1413_n N_Q_c_1795_n 0.0132393f $X=11.2 $Y=1.16 $X2=0 $Y2=0
cc_938 N_A_1738_47#_c_1415_n N_Q_c_1795_n 0.00300434f $X=11.455 $Y=1.217 $X2=0
+ $Y2=0
cc_939 N_A_1738_47#_c_1413_n N_Q_c_1801_n 0.0125866f $X=11.2 $Y=1.16 $X2=0 $Y2=0
cc_940 N_A_1738_47#_c_1415_n N_Q_c_1801_n 0.00404574f $X=11.455 $Y=1.217 $X2=0
+ $Y2=0
cc_941 N_A_1738_47#_M1001_g Q 0.00548163f $X=9.55 $Y=0.56 $X2=0 $Y2=0
cc_942 N_A_1738_47#_M1015_g Q 0.0101751f $X=10.02 $Y=0.56 $X2=0 $Y2=0
cc_943 N_A_1738_47#_M1016_g Q 5.11689e-19 $X=10.49 $Y=0.56 $X2=0 $Y2=0
cc_944 N_A_1738_47#_c_1416_n Q 0.00674155f $X=9.575 $Y=1.41 $X2=0 $Y2=0
cc_945 N_A_1738_47#_c_1417_n Q 0.0127992f $X=10.045 $Y=1.41 $X2=0 $Y2=0
cc_946 N_A_1738_47#_c_1418_n Q 7.03855e-19 $X=10.515 $Y=1.41 $X2=0 $Y2=0
cc_947 N_A_1738_47#_c_1420_n Q 0.00241889f $X=11.455 $Y=1.41 $X2=0 $Y2=0
cc_948 N_A_1738_47#_M1039_g Q 0.019644f $X=11.48 $Y=0.56 $X2=0 $Y2=0
cc_949 N_A_1738_47#_c_1413_n Q 0.0179162f $X=11.2 $Y=1.16 $X2=0 $Y2=0
cc_950 N_A_1738_47#_c_1420_n Q 0.0077888f $X=11.455 $Y=1.41 $X2=0 $Y2=0
cc_951 N_A_1738_47#_M1001_g N_VGND_c_1887_n 0.00317478f $X=9.55 $Y=0.56 $X2=0
+ $Y2=0
cc_952 N_A_1738_47#_c_1413_n N_VGND_c_1887_n 0.00932312f $X=11.2 $Y=1.16 $X2=0
+ $Y2=0
cc_953 N_A_1738_47#_M1015_g N_VGND_c_1888_n 0.00404444f $X=10.02 $Y=0.56 $X2=0
+ $Y2=0
cc_954 N_A_1738_47#_M1016_g N_VGND_c_1888_n 0.0106106f $X=10.49 $Y=0.56 $X2=0
+ $Y2=0
cc_955 N_A_1738_47#_M1018_g N_VGND_c_1888_n 6.59605e-19 $X=10.96 $Y=0.56 $X2=0
+ $Y2=0
cc_956 N_A_1738_47#_M1018_g N_VGND_c_1889_n 0.00170602f $X=10.96 $Y=0.56 $X2=0
+ $Y2=0
cc_957 N_A_1738_47#_M1039_g N_VGND_c_1889_n 0.00976765f $X=11.48 $Y=0.56 $X2=0
+ $Y2=0
cc_958 N_A_1738_47#_c_1412_n N_VGND_c_1890_n 0.0102481f $X=8.815 $Y=0.51 $X2=0
+ $Y2=0
cc_959 N_A_1738_47#_M1001_g N_VGND_c_1895_n 0.00583607f $X=9.55 $Y=0.56 $X2=0
+ $Y2=0
cc_960 N_A_1738_47#_M1015_g N_VGND_c_1895_n 0.00397068f $X=10.02 $Y=0.56 $X2=0
+ $Y2=0
cc_961 N_A_1738_47#_M1016_g N_VGND_c_1896_n 0.00202909f $X=10.49 $Y=0.56 $X2=0
+ $Y2=0
cc_962 N_A_1738_47#_M1018_g N_VGND_c_1896_n 0.00436487f $X=10.96 $Y=0.56 $X2=0
+ $Y2=0
cc_963 N_A_1738_47#_M1039_g N_VGND_c_1897_n 0.00348405f $X=11.48 $Y=0.56 $X2=0
+ $Y2=0
cc_964 N_A_1738_47#_M1006_s N_VGND_c_1898_n 0.00474476f $X=8.69 $Y=0.235 $X2=0
+ $Y2=0
cc_965 N_A_1738_47#_M1001_g N_VGND_c_1898_n 0.0107689f $X=9.55 $Y=0.56 $X2=0
+ $Y2=0
cc_966 N_A_1738_47#_M1015_g N_VGND_c_1898_n 0.00584827f $X=10.02 $Y=0.56 $X2=0
+ $Y2=0
cc_967 N_A_1738_47#_M1016_g N_VGND_c_1898_n 0.00285823f $X=10.49 $Y=0.56 $X2=0
+ $Y2=0
cc_968 N_A_1738_47#_M1018_g N_VGND_c_1898_n 0.00620533f $X=10.96 $Y=0.56 $X2=0
+ $Y2=0
cc_969 N_A_1738_47#_M1039_g N_VGND_c_1898_n 0.00514632f $X=11.48 $Y=0.56 $X2=0
+ $Y2=0
cc_970 N_A_1738_47#_c_1412_n N_VGND_c_1898_n 0.00910216f $X=8.815 $Y=0.51 $X2=0
+ $Y2=0
cc_971 N_VPWR_c_1532_n N_A_409_329#_M1019_d 0.00346917f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_972 N_VPWR_M1019_s N_A_409_329#_c_1728_n 0.00246474f $X=1.595 $Y=1.645 $X2=0
+ $Y2=0
cc_973 N_VPWR_M1019_s N_A_409_329#_c_1735_n 0.00519643f $X=1.595 $Y=1.645 $X2=0
+ $Y2=0
cc_974 N_VPWR_c_1535_n N_A_409_329#_c_1735_n 0.00884569f $X=1.72 $Y=2.22 $X2=0
+ $Y2=0
cc_975 N_VPWR_c_1545_n N_A_409_329#_c_1735_n 0.00242894f $X=3.73 $Y=2.72 $X2=0
+ $Y2=0
cc_976 N_VPWR_c_1532_n N_A_409_329#_c_1735_n 0.00243543f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_977 N_VPWR_M1019_s N_A_409_329#_c_1731_n 0.00197378f $X=1.595 $Y=1.645 $X2=0
+ $Y2=0
cc_978 N_VPWR_c_1534_n N_A_409_329#_c_1731_n 3.86777e-19 $X=1.555 $Y=2.72 $X2=0
+ $Y2=0
cc_979 N_VPWR_c_1535_n N_A_409_329#_c_1731_n 0.0114817f $X=1.72 $Y=2.22 $X2=0
+ $Y2=0
cc_980 N_VPWR_c_1532_n N_A_409_329#_c_1731_n 7.1462e-19 $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_981 N_VPWR_c_1535_n N_A_409_329#_c_1738_n 0.0199789f $X=1.72 $Y=2.22 $X2=0
+ $Y2=0
cc_982 N_VPWR_c_1545_n N_A_409_329#_c_1738_n 0.011801f $X=3.73 $Y=2.72 $X2=0
+ $Y2=0
cc_983 N_VPWR_c_1532_n N_A_409_329#_c_1738_n 0.00307944f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_984 N_VPWR_c_1532_n A_610_413# 0.00374905f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_985 N_VPWR_c_1532_n A_1044_413# 0.00271936f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_986 N_VPWR_c_1532_n A_1244_413# 0.00243108f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_987 N_VPWR_c_1532_n N_Q_M1004_d 0.00444633f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_988 N_VPWR_c_1532_n N_Q_M1014_d 0.00656398f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_989 N_VPWR_c_1532_n N_Q_M1038_d 0.00430086f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_990 N_VPWR_M1008_s N_Q_c_1798_n 0.00187091f $X=10.135 $Y=1.485 $X2=0 $Y2=0
cc_991 N_VPWR_c_1538_n N_Q_c_1798_n 0.0143191f $X=10.28 $Y=2.16 $X2=0 $Y2=0
cc_992 N_VPWR_c_1539_n N_Q_c_1822_n 0.0400915f $X=11.22 $Y=2.02 $X2=0 $Y2=0
cc_993 N_VPWR_c_1549_n N_Q_c_1822_n 0.0118139f $X=11.055 $Y=2.72 $X2=0 $Y2=0
cc_994 N_VPWR_c_1532_n N_Q_c_1822_n 0.00646998f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_995 N_VPWR_M1036_s N_Q_c_1800_n 0.00187091f $X=11.075 $Y=1.485 $X2=0 $Y2=0
cc_996 N_VPWR_c_1539_n N_Q_c_1800_n 0.0210225f $X=11.22 $Y=2.02 $X2=0 $Y2=0
cc_997 N_VPWR_c_1537_n Q 0.0463319f $X=9.34 $Y=2 $X2=0 $Y2=0
cc_998 N_VPWR_c_1542_n Q 0.0167766f $X=10.165 $Y=2.72 $X2=0 $Y2=0
cc_999 N_VPWR_c_1532_n Q 0.0101428f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1000 N_VPWR_c_1539_n Q 0.0503882f $X=11.22 $Y=2.02 $X2=0 $Y2=0
cc_1001 N_VPWR_c_1550_n Q 0.0178516f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1002 N_VPWR_c_1532_n Q 0.00974347f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1003 N_A_409_329#_c_1728_n N_VGND_M1017_s 0.00109524f $X=1.615 $Y=1.795 $X2=0
+ $Y2=0
cc_1004 N_A_409_329#_c_1733_n N_VGND_M1017_s 0.00426381f $X=2.105 $Y=0.73 $X2=0
+ $Y2=0
cc_1005 N_A_409_329#_c_1729_n N_VGND_M1017_s 0.00222201f $X=1.7 $Y=0.73 $X2=0
+ $Y2=0
cc_1006 N_A_409_329#_c_1729_n N_VGND_c_1884_n 4.97798e-19 $X=1.7 $Y=0.73 $X2=0
+ $Y2=0
cc_1007 N_A_409_329#_c_1733_n N_VGND_c_1885_n 0.0105025f $X=2.105 $Y=0.73 $X2=0
+ $Y2=0
cc_1008 N_A_409_329#_c_1729_n N_VGND_c_1885_n 0.0114461f $X=1.7 $Y=0.73 $X2=0
+ $Y2=0
cc_1009 N_A_409_329#_c_1733_n N_VGND_c_1893_n 0.00314004f $X=2.105 $Y=0.73 $X2=0
+ $Y2=0
cc_1010 N_A_409_329#_c_1737_n N_VGND_c_1893_n 0.00861358f $X=2.19 $Y=0.47 $X2=0
+ $Y2=0
cc_1011 N_A_409_329#_M1017_d N_VGND_c_1898_n 0.00308719f $X=2.055 $Y=0.235 $X2=0
+ $Y2=0
cc_1012 N_A_409_329#_c_1733_n N_VGND_c_1898_n 0.00286993f $X=2.105 $Y=0.73 $X2=0
+ $Y2=0
cc_1013 N_A_409_329#_c_1729_n N_VGND_c_1898_n 8.52239e-19 $X=1.7 $Y=0.73 $X2=0
+ $Y2=0
cc_1014 N_A_409_329#_c_1737_n N_VGND_c_1898_n 0.00295275f $X=2.19 $Y=0.47 $X2=0
+ $Y2=0
cc_1015 N_Q_c_1813_n N_VGND_M1015_s 0.00435938f $X=10.665 $Y=0.8 $X2=0 $Y2=0
cc_1016 N_Q_c_1824_n N_VGND_M1018_s 0.00501873f $X=11.605 $Y=0.8 $X2=0 $Y2=0
cc_1017 Q N_VGND_c_1887_n 0.017029f $X=9.8 $Y=0.425 $X2=0 $Y2=0
cc_1018 N_Q_c_1813_n N_VGND_c_1888_n 0.01838f $X=10.665 $Y=0.8 $X2=0 $Y2=0
cc_1019 N_Q_c_1821_n N_VGND_c_1888_n 0.020522f $X=10.75 $Y=0.715 $X2=0 $Y2=0
cc_1020 Q N_VGND_c_1888_n 0.0214241f $X=9.8 $Y=0.425 $X2=0 $Y2=0
cc_1021 N_Q_c_1824_n N_VGND_c_1889_n 0.0220641f $X=11.605 $Y=0.8 $X2=0 $Y2=0
cc_1022 N_Q_c_1813_n N_VGND_c_1895_n 0.00203275f $X=10.665 $Y=0.8 $X2=0 $Y2=0
cc_1023 Q N_VGND_c_1895_n 0.017563f $X=9.8 $Y=0.425 $X2=0 $Y2=0
cc_1024 N_Q_c_1813_n N_VGND_c_1896_n 0.00202593f $X=10.665 $Y=0.8 $X2=0 $Y2=0
cc_1025 N_Q_c_1821_n N_VGND_c_1896_n 0.010834f $X=10.75 $Y=0.715 $X2=0 $Y2=0
cc_1026 N_Q_c_1824_n N_VGND_c_1896_n 0.00259521f $X=11.605 $Y=0.8 $X2=0 $Y2=0
cc_1027 N_Q_c_1824_n N_VGND_c_1897_n 0.0020257f $X=11.605 $Y=0.8 $X2=0 $Y2=0
cc_1028 Q N_VGND_c_1897_n 0.0165824f $X=11.645 $Y=0.425 $X2=0 $Y2=0
cc_1029 N_Q_M1001_d N_VGND_c_1898_n 0.00607858f $X=9.625 $Y=0.235 $X2=0 $Y2=0
cc_1030 N_Q_M1016_d N_VGND_c_1898_n 0.00329764f $X=10.565 $Y=0.235 $X2=0 $Y2=0
cc_1031 N_Q_M1039_d N_VGND_c_1898_n 0.00233692f $X=11.555 $Y=0.235 $X2=0 $Y2=0
cc_1032 N_Q_c_1813_n N_VGND_c_1898_n 0.00949269f $X=10.665 $Y=0.8 $X2=0 $Y2=0
cc_1033 N_Q_c_1821_n N_VGND_c_1898_n 0.00642326f $X=10.75 $Y=0.715 $X2=0 $Y2=0
cc_1034 N_Q_c_1824_n N_VGND_c_1898_n 0.0104497f $X=11.605 $Y=0.8 $X2=0 $Y2=0
cc_1035 Q N_VGND_c_1898_n 0.0110301f $X=9.8 $Y=0.425 $X2=0 $Y2=0
cc_1036 Q N_VGND_c_1898_n 0.00969741f $X=11.645 $Y=0.425 $X2=0 $Y2=0
cc_1037 N_VGND_c_1898_n A_636_47# 0.00226374f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1038 N_VGND_c_1898_n A_866_47# 0.0017066f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1039 N_VGND_c_1898_n A_1156_47# 0.0024588f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1040 N_VGND_c_1898_n A_1344_47# 0.00140476f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1041 N_VGND_c_1898_n A_1416_47# 0.00279792f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
