* File: sky130_fd_sc_hdll__or3b_4.pex.spice
* Created: Wed Sep  2 08:49:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR3B_4%C_N 2 3 5 8 10 11 19
c32 19 0 1.20913e-19 $X=0.52 $Y=1.16
c33 8 0 1.38818e-19 $X=0.52 $Y=0.445
r34 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r35 15 18 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.495 $Y2=1.16
r36 10 11 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.16
+ $X2=0.255 $Y2=1.53
r37 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r38 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r39 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r40 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.725
+ $X2=0.495 $Y2=2.01
r41 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.625 $X2=0.495
+ $Y2=1.725
r42 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r43 1 2 99.4732 $w=2e-07 $l=3e-07 $layer=POLY_cond $X=0.495 $Y=1.325 $X2=0.495
+ $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_4%A_186_21# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 43 44 45 50 55 64
c127 45 0 1.91481e-19 $X=2.615 $Y=0.74
c128 19 0 9.42572e-20 $X=1.5 $Y=1.41
c129 13 0 1.43265e-20 $X=1.03 $Y=1.41
r130 64 65 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.44 $Y=1.202
+ $X2=2.465 $Y2=1.202
r131 61 62 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.945 $Y=1.202
+ $X2=1.97 $Y2=1.202
r132 58 59 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.475 $Y=1.202
+ $X2=1.5 $Y2=1.202
r133 57 58 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=1.03 $Y=1.202
+ $X2=1.475 $Y2=1.202
r134 56 57 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.005 $Y=1.202
+ $X2=1.03 $Y2=1.202
r135 54 55 74.9313 $w=2.03e-07 $l=1.385e-06 $layer=LI1_cond $X=4.352 $Y=0.825
+ $X2=4.352 $Y2=2.21
r136 50 55 6.82152 $w=2.15e-07 $l=1.49543e-07 $layer=LI1_cond $X=4.25 $Y=2.317
+ $X2=4.352 $Y2=2.21
r137 50 52 5.62821 $w=2.13e-07 $l=1.05e-07 $layer=LI1_cond $X=4.25 $Y=2.317
+ $X2=4.145 $Y2=2.317
r138 47 49 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.145 $Y=0.74
+ $X2=4.145 $Y2=0.74
r139 45 47 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.615 $Y=0.74
+ $X2=3.145 $Y2=0.74
r140 44 54 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=4.25 $Y=0.74
+ $X2=4.352 $Y2=0.825
r141 44 49 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.25 $Y=0.74
+ $X2=4.145 $Y2=0.74
r142 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.53 $Y=0.825
+ $X2=2.615 $Y2=0.74
r143 42 43 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.53 $Y=0.825
+ $X2=2.53 $Y2=1.075
r144 41 64 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=2.405 $Y=1.202
+ $X2=2.44 $Y2=1.202
r145 41 62 56.3629 $w=3.72e-07 $l=4.35e-07 $layer=POLY_cond $X=2.405 $Y=1.202
+ $X2=1.97 $Y2=1.202
r146 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.405
+ $Y=1.16 $X2=2.405 $Y2=1.16
r147 37 61 41.4624 $w=3.72e-07 $l=3.2e-07 $layer=POLY_cond $X=1.625 $Y=1.202
+ $X2=1.945 $Y2=1.202
r148 37 59 16.1962 $w=3.72e-07 $l=1.25e-07 $layer=POLY_cond $X=1.625 $Y=1.202
+ $X2=1.5 $Y2=1.202
r149 36 40 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.625 $Y=1.16
+ $X2=2.405 $Y2=1.16
r150 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.16 $X2=1.625 $Y2=1.16
r151 34 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=1.16
+ $X2=2.53 $Y2=1.075
r152 34 40 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.445 $Y=1.16
+ $X2=2.405 $Y2=1.16
r153 31 65 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.465 $Y=0.995
+ $X2=2.465 $Y2=1.202
r154 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.465 $Y=0.995
+ $X2=2.465 $Y2=0.56
r155 28 64 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.44 $Y=1.41
+ $X2=2.44 $Y2=1.202
r156 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.44 $Y=1.41
+ $X2=2.44 $Y2=1.985
r157 25 62 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.97 $Y=1.41
+ $X2=1.97 $Y2=1.202
r158 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.97 $Y=1.41
+ $X2=1.97 $Y2=1.985
r159 22 61 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.945 $Y=0.995
+ $X2=1.945 $Y2=1.202
r160 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.945 $Y=0.995
+ $X2=1.945 $Y2=0.56
r161 19 59 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.5 $Y2=1.202
r162 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.5 $Y2=1.985
r163 16 58 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=1.202
r164 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=0.56
r165 13 57 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.202
r166 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.985
r167 10 56 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=1.202
r168 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.56
r169 3 52 600 $w=1.7e-07 $l=8.79517e-07 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=1.485 $X2=4.145 $Y2=2.295
r170 2 49 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=3.96
+ $Y=0.235 $X2=4.145 $Y2=0.74
r171 1 47 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.235 $X2=3.145 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_4%A 1 3 4 6 7 11
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.885
+ $Y=1.16 $X2=2.885 $Y2=1.16
r36 7 11 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.955 $Y=1.53
+ $X2=2.955 $Y2=1.16
r37 4 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=2.935 $Y=0.995
+ $X2=2.91 $Y2=1.16
r38 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.935 $Y=0.995
+ $X2=2.935 $Y2=0.56
r39 1 10 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.91 $Y=1.41
+ $X2=2.91 $Y2=1.16
r40 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.91 $Y=1.41 $X2=2.91
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_4%B 1 3 4 6 7 8
r28 7 8 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.45 $Y=1.16 $X2=3.45
+ $Y2=1.53
r29 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=1.16 $X2=3.415 $Y2=1.16
r30 4 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.44 $Y2=1.16
r31 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.38 $Y=1.41 $X2=3.38
+ $Y2=1.985
r32 1 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.355 $Y=0.995
+ $X2=3.44 $Y2=1.16
r33 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.355 $Y=0.995
+ $X2=3.355 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_4%A_27_47# 1 2 7 9 10 12 15 17 18 19 22 23 27
+ 32 34
c92 32 0 1.43265e-20 $X=0.26 $Y=1.975
c93 19 0 1.20913e-19 $X=0.645 $Y=1.925
r94 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.945
+ $Y=1.16 $X2=3.945 $Y2=1.16
r95 25 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.945 $Y=1.87
+ $X2=3.945 $Y2=1.16
r96 24 34 4.50329 $w=2e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.815 $Y=1.955
+ $X2=0.73 $Y2=1.925
r97 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.86 $Y=1.955
+ $X2=3.945 $Y2=1.87
r98 23 24 198.658 $w=1.68e-07 $l=3.045e-06 $layer=LI1_cond $X=3.86 $Y=1.955
+ $X2=0.815 $Y2=1.955
r99 22 34 1.93381 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.73 $Y=1.81
+ $X2=0.73 $Y2=1.925
r100 21 22 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=0.73 $Y=0.905
+ $X2=0.73 $Y2=1.81
r101 20 32 1.45362 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.925
+ $X2=0.215 $Y2=1.925
r102 19 34 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.645 $Y=1.925
+ $X2=0.73 $Y2=1.925
r103 19 20 15.0319 $w=2.28e-07 $l=3e-07 $layer=LI1_cond $X=0.645 $Y=1.925
+ $X2=0.345 $Y2=1.925
r104 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.73 $Y2=0.905
r105 17 18 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.345 $Y2=0.82
r106 13 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.735
+ $X2=0.345 $Y2=0.82
r107 13 15 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=0.215 $Y=0.735
+ $X2=0.215 $Y2=0.455
r108 10 28 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=3.91 $Y=1.41
+ $X2=3.97 $Y2=1.16
r109 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.91 $Y=1.41
+ $X2=3.91 $Y2=1.985
r110 7 28 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.885 $Y=0.995
+ $X2=3.97 $Y2=1.16
r111 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.885 $Y=0.995
+ $X2=3.885 $Y2=0.56
r112 2 32 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.8 $X2=0.26 $Y2=1.975
r113 1 15 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_4%VPWR 1 2 3 12 16 18 22 24 26 31 41 42 45 48
+ 51
r65 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r66 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r67 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r70 39 42 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r71 39 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 38 41 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r73 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r74 36 51 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=2.65 $Y2=2.72
r75 36 38 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=2.99 $Y2=2.72
r76 35 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 35 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r79 32 45 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.96 $Y=2.72 $X2=0.78
+ $Y2=2.72
r80 32 34 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.96 $Y=2.72
+ $X2=1.15 $Y2=2.72
r81 31 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.52 $Y=2.72 $X2=1.71
+ $Y2=2.72
r82 31 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.52 $Y=2.72 $X2=1.15
+ $Y2=2.72
r83 26 45 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.78
+ $Y2=2.72
r84 26 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r85 24 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r87 20 51 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=2.635
+ $X2=2.65 $Y2=2.72
r88 20 22 10.0469 $w=3.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.65 $Y=2.635
+ $X2=2.65 $Y2=2.295
r89 19 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.9 $Y=2.72 $X2=1.71
+ $Y2=2.72
r90 18 51 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=2.65 $Y2=2.72
r91 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=1.9 $Y2=2.72
r92 14 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=2.635
+ $X2=1.71 $Y2=2.72
r93 14 16 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.71 $Y=2.635
+ $X2=1.71 $Y2=2.295
r94 10 45 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=2.635
+ $X2=0.78 $Y2=2.72
r95 10 12 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.78 $Y=2.635
+ $X2=0.78 $Y2=2.295
r96 3 22 600 $w=1.7e-07 $l=8.79517e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.485 $X2=2.675 $Y2=2.295
r97 2 16 600 $w=1.7e-07 $l=8.79517e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.485 $X2=1.735 $Y2=2.295
r98 1 12 600 $w=1.7e-07 $l=5.90741e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.8 $X2=0.795 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_4%X 1 2 3 4 15 18 19 23 25 29 34
c59 25 0 1.38818e-19 $X=1.22 $Y=0.82
c60 18 0 9.42572e-20 $X=1.14 $Y=1.415
r61 29 34 3.03274 $w=2.83e-07 $l=7.5e-08 $layer=LI1_cond $X=2.205 $Y=1.557
+ $X2=2.28 $Y2=1.557
r62 26 29 37.8082 $w=2.83e-07 $l=9.35e-07 $layer=LI1_cond $X=1.27 $Y=1.557
+ $X2=2.205 $Y2=1.557
r63 26 28 3.26681 $w=2.85e-07 $l=1.3e-07 $layer=LI1_cond $X=1.27 $Y=1.557
+ $X2=1.14 $Y2=1.557
r64 21 23 15.4476 $w=2.33e-07 $l=3.15e-07 $layer=LI1_cond $X=2.122 $Y=0.735
+ $X2=2.122 $Y2=0.42
r65 20 25 3.9231 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.43 $Y=0.82 $X2=1.22
+ $Y2=0.82
r66 19 21 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.005 $Y=0.82
+ $X2=2.122 $Y2=0.735
r67 19 20 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.005 $Y=0.82
+ $X2=1.43 $Y2=0.82
r68 18 28 3.56836 $w=2.6e-07 $l=1.42e-07 $layer=LI1_cond $X=1.14 $Y=1.415
+ $X2=1.14 $Y2=1.557
r69 17 25 2.80976 $w=3.4e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.14 $Y=0.905
+ $X2=1.22 $Y2=0.82
r70 17 18 22.6056 $w=2.58e-07 $l=5.1e-07 $layer=LI1_cond $X=1.14 $Y=0.905
+ $X2=1.14 $Y2=1.415
r71 13 25 2.80976 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.735
+ $X2=1.22 $Y2=0.82
r72 13 15 9.3293 $w=4.18e-07 $l=3.4e-07 $layer=LI1_cond $X=1.22 $Y=0.735
+ $X2=1.22 $Y2=0.395
r73 4 29 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=2.06
+ $Y=1.485 $X2=2.205 $Y2=1.615
r74 3 28 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.615
r75 2 23 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.235 $X2=2.155 $Y2=0.42
r76 1 15 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=1.08
+ $Y=0.235 $X2=1.265 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_4%VGND 1 2 3 4 17 21 23 27 29 31 32 33 41 42
+ 45 48 52 58
c73 3 0 1.91481e-19 $X=2.54 $Y=0.235
r74 52 55 10.4768 $w=4.38e-07 $l=4e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.62
+ $Y2=0.4
r75 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r76 49 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r77 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r78 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r79 42 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r80 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r81 39 52 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=3.62
+ $Y2=0
r82 39 41 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=4.37
+ $Y2=0
r83 38 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r84 38 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r85 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r86 35 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=0 $X2=0.755
+ $Y2=0
r87 35 37 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.84 $Y=0 $X2=1.61
+ $Y2=0
r88 33 46 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r89 33 58 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r90 31 37 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.61
+ $Y2=0
r91 31 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.735
+ $Y2=0
r92 30 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.84 $Y=0 $X2=2.65
+ $Y2=0
r93 29 52 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.62
+ $Y2=0
r94 29 30 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=2.84
+ $Y2=0
r95 25 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=0.085
+ $X2=2.65 $Y2=0
r96 25 27 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.65 $Y=0.085
+ $X2=2.65 $Y2=0.4
r97 24 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.82 $Y=0 $X2=1.735
+ $Y2=0
r98 23 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.65
+ $Y2=0
r99 23 24 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=1.82
+ $Y2=0
r100 19 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0
r101 19 21 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0.4
r102 15 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r103 15 17 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.4
r104 4 55 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.235 $X2=3.615 $Y2=0.4
r105 3 27 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.54
+ $Y=0.235 $X2=2.675 $Y2=0.4
r106 2 21 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.235 $X2=1.735 $Y2=0.4
r107 1 17 182 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.755 $Y2=0.4
.ends

