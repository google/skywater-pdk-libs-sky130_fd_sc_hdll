* File: sky130_fd_sc_hdll__xnor3_4.pex.spice
* Created: Wed Sep  2 08:54:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%A_101_21# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 32 33 35 36 38 40 42 43 45 47 49 55 63
c142 13 0 1.63304e-19 $X=1.05 $Y=0.995
r143 62 63 5.91008 $w=3.67e-07 $l=4.5e-08 $layer=POLY_cond $X=2 $Y=1.202
+ $X2=2.045 $Y2=1.202
r144 61 62 55.8174 $w=3.67e-07 $l=4.25e-07 $layer=POLY_cond $X=1.575 $Y=1.202
+ $X2=2 $Y2=1.202
r145 60 61 5.91008 $w=3.67e-07 $l=4.5e-08 $layer=POLY_cond $X=1.53 $Y=1.202
+ $X2=1.575 $Y2=1.202
r146 59 60 59.7575 $w=3.67e-07 $l=4.55e-07 $layer=POLY_cond $X=1.075 $Y=1.202
+ $X2=1.53 $Y2=1.202
r147 58 59 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.05 $Y=1.202
+ $X2=1.075 $Y2=1.202
r148 57 58 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=0.605 $Y=1.202
+ $X2=1.05 $Y2=1.202
r149 56 57 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.58 $Y=1.202
+ $X2=0.605 $Y2=1.202
r150 54 63 9.19346 $w=3.67e-07 $l=7e-08 $layer=POLY_cond $X=2.115 $Y=1.202
+ $X2=2.045 $Y2=1.202
r151 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=1.16 $X2=2.115 $Y2=1.16
r152 51 53 19.3167 $w=2.4e-07 $l=3.8e-07 $layer=LI1_cond $X=2.157 $Y=0.78
+ $X2=2.157 $Y2=1.16
r153 47 55 11.3723 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=3.9 $Y=0.355 $X2=3.7
+ $Y2=0.355
r154 47 49 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=3.9 $Y=0.355
+ $X2=4.02 $Y2=0.355
r155 43 45 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=2.85 $Y=2.32
+ $X2=3.945 $Y2=2.32
r156 42 55 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=2.735 $Y=0.34
+ $X2=3.7 $Y2=0.34
r157 40 43 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.74 $Y=2.235
+ $X2=2.85 $Y2=2.32
r158 39 40 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=2.74 $Y=2.045
+ $X2=2.74 $Y2=2.235
r159 37 42 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.625 $Y=0.425
+ $X2=2.735 $Y2=0.34
r160 37 38 14.1436 $w=2.18e-07 $l=2.7e-07 $layer=LI1_cond $X=2.625 $Y=0.425
+ $X2=2.625 $Y2=0.695
r161 35 39 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.63 $Y=1.96
+ $X2=2.74 $Y2=2.045
r162 35 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.63 $Y=1.96
+ $X2=2.285 $Y2=1.96
r163 34 51 2.75731 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.285 $Y=0.78
+ $X2=2.157 $Y2=0.78
r164 33 38 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.515 $Y=0.78
+ $X2=2.625 $Y2=0.695
r165 33 34 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.515 $Y=0.78
+ $X2=2.285 $Y2=0.78
r166 32 36 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.175 $Y=1.875
+ $X2=2.285 $Y2=1.96
r167 31 53 8.49444 $w=2.4e-07 $l=1.73767e-07 $layer=LI1_cond $X=2.175 $Y=1.325
+ $X2=2.157 $Y2=1.16
r168 31 32 28.8111 $w=2.18e-07 $l=5.5e-07 $layer=LI1_cond $X=2.175 $Y=1.325
+ $X2=2.175 $Y2=1.875
r169 28 63 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.045 $Y=1.41
+ $X2=2.045 $Y2=1.202
r170 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.045 $Y=1.41
+ $X2=2.045 $Y2=1.985
r171 25 62 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2 $Y=0.995 $X2=2
+ $Y2=1.202
r172 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2 $Y=0.995 $X2=2
+ $Y2=0.56
r173 22 61 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.575 $Y=1.41
+ $X2=1.575 $Y2=1.202
r174 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.575 $Y=1.41
+ $X2=1.575 $Y2=1.985
r175 19 60 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=1.202
r176 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=0.56
r177 16 59 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.075 $Y=1.41
+ $X2=1.075 $Y2=1.202
r178 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.075 $Y=1.41
+ $X2=1.075 $Y2=1.985
r179 13 58 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.05 $Y=0.995
+ $X2=1.05 $Y2=1.202
r180 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.05 $Y=0.995
+ $X2=1.05 $Y2=0.56
r181 10 57 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.605 $Y=1.41
+ $X2=0.605 $Y2=1.202
r182 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.605 $Y=1.41
+ $X2=0.605 $Y2=1.985
r183 7 56 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.58 $Y2=1.202
r184 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.58 $Y2=0.56
r185 2 45 600 $w=1.7e-07 $l=7.64068e-07 $layer=licon1_PDIFF $count=1 $X=3.8
+ $Y=1.625 $X2=3.945 $Y2=2.32
r186 1 49 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.245 $X2=4.02 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%C 1 3 7 8 10 11 13 15 18 19 23 25
c60 1 0 1.70967e-19 $X=2.585 $Y=0.995
r61 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.545
+ $Y=1.16 $X2=3.545 $Y2=1.16
r62 19 23 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.455 $Y=1.2 $X2=3.545
+ $Y2=1.2
r63 19 25 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.455 $Y=1.2 $X2=3.45
+ $Y2=1.2
r64 18 22 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.61 $Y=1.16
+ $X2=3.545 $Y2=1.16
r65 14 22 146.009 $w=3.3e-07 $l=8.35e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=3.545 $Y2=1.16
r66 14 15 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=2.61 $Y2=1.202
r67 11 18 39.7875 $w=2.42e-07 $l=1.9182e-07 $layer=POLY_cond $X=3.8 $Y=0.995
+ $X2=3.742 $Y2=1.16
r68 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.8 $Y=0.995 $X2=3.8
+ $Y2=0.565
r69 8 18 80.9439 $w=2.42e-07 $l=4.05685e-07 $layer=POLY_cond $X=3.71 $Y=1.55
+ $X2=3.742 $Y2=1.16
r70 8 10 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=3.71 $Y=1.55 $X2=3.71
+ $Y2=2.045
r71 4 15 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=2.61 $Y=1.41
+ $X2=2.61 $Y2=1.202
r72 4 7 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.61 $Y=1.41 $X2=2.61
+ $Y2=1.805
r73 1 15 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=2.585 $Y=0.995
+ $X2=2.61 $Y2=1.202
r74 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.585 $Y=0.995
+ $X2=2.585 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%A_532_93# 1 2 7 9 10 12 13 18 20 23 24 28
r72 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.22
+ $Y=1.16 $X2=4.22 $Y2=1.16
r73 25 28 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.115 $Y=1.16
+ $X2=4.22 $Y2=1.16
r74 22 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.115 $Y=1.325
+ $X2=4.115 $Y2=1.16
r75 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.115 $Y=1.325
+ $X2=4.115 $Y2=1.535
r76 21 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=1.62
+ $X2=2.99 $Y2=1.62
r77 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.03 $Y=1.62
+ $X2=4.115 $Y2=1.535
r78 20 21 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.03 $Y=1.62
+ $X2=3.075 $Y2=1.62
r79 16 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=1.535
+ $X2=2.99 $Y2=1.62
r80 16 18 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.99 $Y=1.535
+ $X2=2.99 $Y2=0.76
r81 13 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=1.62
+ $X2=2.99 $Y2=1.62
r82 13 15 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=2.905 $Y=1.62 $X2=2.845
+ $Y2=1.62
r83 10 29 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=4.33 $Y=0.995
+ $X2=4.245 $Y2=1.16
r84 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.33 $Y=0.995
+ $X2=4.33 $Y2=0.565
r85 7 29 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=4.245 $Y=1.41
+ $X2=4.245 $Y2=1.16
r86 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=4.245 $Y=1.41
+ $X2=4.245 $Y2=1.905
r87 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.485 $X2=2.845 $Y2=1.62
r88 1 18 182 $w=1.7e-07 $l=4.54148e-07 $layer=licon1_NDIFF $count=1 $X=2.66
+ $Y=0.465 $X2=2.99 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%A_1089_297# 1 2 7 9 12 14 15 16 18 19 21
+ 22 23 27 35 37 38 39 40 47 49 50 58
c180 37 0 1.57566e-19 $X=7.025 $Y=0.85
c181 27 0 1.36535e-19 $X=5.75 $Y=1.58
c182 14 0 1.24749e-19 $X=8.85 $Y=1.28
r183 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.77
+ $Y=1.11 $X2=8.77 $Y2=1.11
r184 50 56 11.8358 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.7 $Y=0.85 $X2=8.7
+ $Y2=1.11
r185 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.65 $Y=0.85
+ $X2=8.65 $Y2=0.85
r186 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.17 $Y=0.85
+ $X2=7.17 $Y2=0.85
r187 42 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.69 $Y=0.85
+ $X2=5.69 $Y2=0.85
r188 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.315 $Y=0.85
+ $X2=7.17 $Y2=0.85
r189 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.505 $Y=0.85
+ $X2=8.65 $Y2=0.85
r190 39 40 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=8.505 $Y=0.85
+ $X2=7.315 $Y2=0.85
r191 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.835 $Y=0.85
+ $X2=5.69 $Y2=0.85
r192 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.025 $Y=0.85
+ $X2=7.17 $Y2=0.85
r193 37 38 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=7.025 $Y=0.85
+ $X2=5.835 $Y2=0.85
r194 35 47 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=7.15 $Y=0.995
+ $X2=7.15 $Y2=0.85
r195 31 35 6.28605 $w=2.73e-07 $l=1.5e-07 $layer=LI1_cond $X=7 $Y=1.132 $X2=7.15
+ $Y2=1.132
r196 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7 $Y=1.16
+ $X2=7 $Y2=1.16
r197 28 58 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=5.75 $Y=1.445
+ $X2=5.75 $Y2=0.74
r198 27 28 0.275955 $w=2.9e-07 $l=1.35e-07 $layer=LI1_cond $X=5.75 $Y=1.58
+ $X2=5.75 $Y2=1.445
r199 25 27 6.82929 $w=2.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.59 $Y=1.58
+ $X2=5.75 $Y2=1.58
r200 22 32 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=7.26 $Y=1.16 $X2=7
+ $Y2=1.16
r201 22 23 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=7.26 $Y=1.16
+ $X2=7.36 $Y2=1.202
r202 19 55 38.5432 $w=3.18e-07 $l=2.03101e-07 $layer=POLY_cond $X=8.88 $Y=0.945
+ $X2=8.795 $Y2=1.11
r203 19 21 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.88 $Y=0.945
+ $X2=8.88 $Y2=0.535
r204 16 18 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.85 $Y=1.57
+ $X2=8.85 $Y2=2.065
r205 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.85 $Y=1.47 $X2=8.85
+ $Y2=1.57
r206 14 55 32.3713 $w=3.18e-07 $l=1.95576e-07 $layer=POLY_cond $X=8.85 $Y=1.28
+ $X2=8.795 $Y2=1.11
r207 14 15 62.9997 $w=2e-07 $l=1.9e-07 $layer=POLY_cond $X=8.85 $Y=1.28 $X2=8.85
+ $Y2=1.47
r208 10 23 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=7.385 $Y=0.995
+ $X2=7.36 $Y2=1.202
r209 10 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.385 $Y=0.995
+ $X2=7.385 $Y2=0.455
r210 7 23 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=7.36 $Y=1.41
+ $X2=7.36 $Y2=1.202
r211 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=7.36 $Y=1.41
+ $X2=7.36 $Y2=1.805
r212 2 25 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.445
+ $Y=1.485 $X2=5.59 $Y2=1.63
r213 1 58 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=5.625
+ $Y=0.235 $X2=5.81 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%B 1 3 6 8 9 13 16 18 19 22 24 25 28 31 35
+ 36 38 39 42 45
c134 39 0 1.94872e-19 $X=8.445 $Y=1.445
r135 39 45 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=8.53 $Y=1.53
+ $X2=8.465 $Y2=1.53
r136 38 45 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.375 $Y=1.53
+ $X2=8.465 $Y2=1.53
r137 36 43 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.265 $Y=1.16
+ $X2=8.265 $Y2=1.325
r138 36 42 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.265 $Y=1.16
+ $X2=8.265 $Y2=0.995
r139 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.24
+ $Y=1.16 $X2=8.24 $Y2=1.16
r140 33 38 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=8.265 $Y=1.445
+ $X2=8.375 $Y2=1.53
r141 33 35 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=8.265 $Y=1.445
+ $X2=8.265 $Y2=1.16
r142 31 32 29.1618 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=6.555 $Y=1.16
+ $X2=6.555 $Y2=1.085
r143 26 28 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=8.285 $Y=2.415
+ $X2=8.285 $Y2=1.965
r144 25 28 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=8.285 $Y=1.57
+ $X2=8.285 $Y2=1.965
r145 24 25 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.285 $Y=1.47 $X2=8.285
+ $Y2=1.57
r146 24 43 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=8.285 $Y=1.47
+ $X2=8.285 $Y2=1.325
r147 22 42 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.18 $Y=0.565
+ $X2=8.18 $Y2=0.995
r148 18 26 27.2212 $w=1.5e-07 $l=1.67705e-07 $layer=POLY_cond $X=8.185 $Y=2.54
+ $X2=8.285 $Y2=2.415
r149 18 19 784.532 $w=1.5e-07 $l=1.53e-06 $layer=POLY_cond $X=8.185 $Y=2.54
+ $X2=6.655 $Y2=2.54
r150 16 32 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.58 $Y=0.565
+ $X2=6.58 $Y2=1.085
r151 11 19 27.2212 $w=1.5e-07 $l=1.36015e-07 $layer=POLY_cond $X=6.555 $Y=2.455
+ $X2=6.655 $Y2=2.54
r152 11 13 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=6.555 $Y=2.455
+ $X2=6.555 $Y2=1.905
r153 10 31 83.702 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=6.555 $Y=1.41
+ $X2=6.555 $Y2=1.16
r154 10 13 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=6.555 $Y=1.41
+ $X2=6.555 $Y2=1.905
r155 8 31 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=6.455 $Y=1.16
+ $X2=6.555 $Y2=1.16
r156 8 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=6.455 $Y=1.16
+ $X2=5.625 $Y2=1.16
r157 4 9 21.9219 $w=2.44e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.55 $Y=1.085
+ $X2=5.625 $Y2=1.16
r158 4 29 38.5205 $w=2.44e-07 $l=2.63847e-07 $layer=POLY_cond $X=5.55 $Y=1.085
+ $X2=5.355 $Y2=1.247
r159 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.55 $Y=1.085
+ $X2=5.55 $Y2=0.56
r160 1 29 9.95785 $w=1.8e-07 $l=1.63e-07 $layer=POLY_cond $X=5.355 $Y=1.41
+ $X2=5.355 $Y2=1.247
r161 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.355 $Y=1.41
+ $X2=5.355 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%A 1 3 4 6 7
c38 1 0 1.94872e-19 $X=9.405 $Y=1.41
r39 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.3 $Y=1.16
+ $X2=9.3 $Y2=1.16
r40 4 10 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=9.43 $Y=0.995
+ $X2=9.335 $Y2=1.16
r41 4 6 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=9.43 $Y=0.995 $X2=9.43
+ $Y2=0.555
r42 1 10 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=9.405 $Y=1.41
+ $X2=9.335 $Y2=1.16
r43 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.405 $Y=1.41
+ $X2=9.405 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%A_1207_297# 1 2 3 4 13 15 16 18 19 21 23
+ 27 28 29 30 37 38 41 44 45
c135 30 0 1.07404e-19 $X=9.79 $Y=1.495
c136 13 0 3.96944e-20 $X=9.875 $Y=1.41
r137 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.16 $Y=0.51
+ $X2=9.16 $Y2=0.51
r138 41 50 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=6.16 $Y=0.51
+ $X2=6.16 $Y2=1.94
r139 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.16 $Y=0.51
+ $X2=6.16 $Y2=0.51
r140 38 40 0.121883 $w=2.3e-07 $l=1.55e-07 $layer=MET1_cond $X=6.315 $Y=0.51
+ $X2=6.16 $Y2=0.51
r141 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.015 $Y=0.51
+ $X2=9.16 $Y2=0.51
r142 37 38 3.34158 $w=1.4e-07 $l=2.7e-06 $layer=MET1_cond $X=9.015 $Y=0.51
+ $X2=6.315 $Y2=0.51
r143 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.85
+ $Y=1.16 $X2=9.85 $Y2=1.16
r144 33 35 17.9567 $w=2.31e-07 $l=3.4e-07 $layer=LI1_cond $X=9.845 $Y=0.82
+ $X2=9.845 $Y2=1.16
r145 32 45 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=9.19 $Y=0.735
+ $X2=9.19 $Y2=0.51
r146 31 41 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=6.16 $Y=0.485
+ $X2=6.16 $Y2=0.51
r147 29 35 9.58904 $w=2.31e-07 $l=1.90526e-07 $layer=LI1_cond $X=9.79 $Y=1.325
+ $X2=9.845 $Y2=1.16
r148 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.79 $Y=1.325
+ $X2=9.79 $Y2=1.495
r149 28 32 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=9.335 $Y=0.82
+ $X2=9.19 $Y2=0.735
r150 27 33 2.5345 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=9.705 $Y=0.82
+ $X2=9.845 $Y2=0.82
r151 27 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.705 $Y=0.82
+ $X2=9.335 $Y2=0.82
r152 23 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=9.705 $Y=1.6
+ $X2=9.79 $Y2=1.495
r153 23 25 28.2554 $w=2.08e-07 $l=5.35e-07 $layer=LI1_cond $X=9.705 $Y=1.6
+ $X2=9.17 $Y2=1.6
r154 19 31 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.245 $Y=0.375
+ $X2=6.16 $Y2=0.485
r155 19 21 5.76222 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=6.245 $Y=0.375
+ $X2=6.355 $Y2=0.375
r156 16 36 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=9.9 $Y=0.995
+ $X2=9.875 $Y2=1.16
r157 16 18 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=9.9 $Y=0.995
+ $X2=9.9 $Y2=0.555
r158 13 36 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=9.875 $Y=1.41
+ $X2=9.875 $Y2=1.16
r159 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.875 $Y=1.41
+ $X2=9.875 $Y2=1.985
r160 4 25 600 $w=1.7e-07 $l=2.42178e-07 $layer=licon1_PDIFF $count=1 $X=8.94
+ $Y=1.645 $X2=9.17 $Y2=1.62
r161 3 50 600 $w=1.7e-07 $l=5.13712e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=1.485 $X2=6.16 $Y2=1.94
r162 2 45 182 $w=1.7e-07 $l=4.85747e-07 $layer=licon1_NDIFF $count=1 $X=8.955
+ $Y=0.235 $X2=9.17 $Y2=0.625
r163 1 21 182 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_NDIFF $count=1 $X=6.205
+ $Y=0.245 $X2=6.355 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%VPWR 1 2 3 4 5 18 24 28 32 36 39 40 41 42
+ 44 45 46 61 67 68 71 74
c117 5 0 1.07404e-19 $X=9.495 $Y=1.485
r118 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r119 68 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=9.43 $Y2=2.72
r120 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r121 65 67 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=9.81 $Y=2.72
+ $X2=10.35 $Y2=2.72
r122 64 78 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=9.43 $Y2=2.72
r123 63 64 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r124 61 65 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=9.617 $Y=2.72
+ $X2=9.81 $Y2=2.72
r125 61 78 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r126 61 74 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=9.617 $Y=2.72
+ $X2=9.617 $Y2=2.36
r127 61 63 269.77 $w=1.68e-07 $l=4.135e-06 $layer=LI1_cond $X=9.425 $Y=2.72
+ $X2=5.29 $Y2=2.72
r128 60 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r129 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r130 57 60 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r131 57 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r132 56 59 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r133 56 57 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r134 54 71 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.45 $Y=2.72
+ $X2=2.257 $Y2=2.72
r135 54 56 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.45 $Y=2.72 $X2=2.53
+ $Y2=2.72
r136 53 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r137 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r138 46 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r139 46 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r140 44 59 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=4.83 $Y2=2.72
r141 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=5.12 $Y2=2.72
r142 43 63 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.285 $Y=2.72
+ $X2=5.29 $Y2=2.72
r143 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=2.72
+ $X2=5.12 $Y2=2.72
r144 41 52 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.225 $Y=2.72
+ $X2=1.15 $Y2=2.72
r145 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=2.72
+ $X2=1.31 $Y2=2.72
r146 39 49 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.285 $Y=2.72
+ $X2=0.23 $Y2=2.72
r147 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=2.72
+ $X2=0.37 $Y2=2.72
r148 38 52 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r149 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.455 $Y=2.72
+ $X2=0.37 $Y2=2.72
r150 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=2.635
+ $X2=5.12 $Y2=2.72
r151 34 36 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.12 $Y=2.635
+ $X2=5.12 $Y2=2.32
r152 30 71 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.257 $Y=2.635
+ $X2=2.257 $Y2=2.72
r153 30 32 10.0278 $w=3.83e-07 $l=3.35e-07 $layer=LI1_cond $X=2.257 $Y=2.635
+ $X2=2.257 $Y2=2.3
r154 29 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.31 $Y2=2.72
r155 28 71 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=2.257 $Y2=2.72
r156 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=1.395 $Y2=2.72
r157 24 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.31 $Y=1.66
+ $X2=1.31 $Y2=2.34
r158 22 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=2.635
+ $X2=1.31 $Y2=2.72
r159 22 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.31 $Y=2.635
+ $X2=1.31 $Y2=2.34
r160 18 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.37 $Y=1.66
+ $X2=0.37 $Y2=2.34
r161 16 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.37 $Y=2.635
+ $X2=0.37 $Y2=2.72
r162 16 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.37 $Y=2.635
+ $X2=0.37 $Y2=2.34
r163 5 74 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=9.495
+ $Y=1.485 $X2=9.64 $Y2=2.36
r164 4 36 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.995
+ $Y=2.175 $X2=5.12 $Y2=2.32
r165 3 32 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=2.135
+ $Y=1.485 $X2=2.285 $Y2=2.3
r166 2 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.165
+ $Y=1.485 $X2=1.31 $Y2=2.34
r167 2 24 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.165
+ $Y=1.485 $X2=1.31 $Y2=1.66
r168 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.485 $X2=0.37 $Y2=2.34
r169 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.485 $X2=0.37 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%X 1 2 3 4 15 19 23 27 29 30 32 35
c44 27 0 1.63304e-19 $X=1.79 $Y=0.56
r45 32 39 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.73 $Y=1.87
+ $X2=1.73 $Y2=2.3
r46 32 35 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.73 $Y=1.87
+ $X2=1.73 $Y2=1.62
r47 30 35 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.73 $Y=1.605
+ $X2=1.73 $Y2=1.62
r48 30 31 16.5482 $w=3.3e-07 $l=4.45e-07 $layer=LI1_cond $X=1.73 $Y=1.605
+ $X2=1.73 $Y2=1.16
r49 25 31 15.3484 $w=3.1e-07 $l=3.94968e-07 $layer=LI1_cond $X=1.72 $Y=0.77
+ $X2=1.73 $Y2=1.16
r50 25 27 7.80687 $w=3.08e-07 $l=2.1e-07 $layer=LI1_cond $X=1.72 $Y=0.77
+ $X2=1.72 $Y2=0.56
r51 24 29 1.45028 $w=3.3e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=1.16
+ $X2=0.815 $Y2=1.16
r52 23 31 0.209703 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=1.16
+ $X2=1.73 $Y2=1.16
r53 23 24 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.565 $Y=1.16
+ $X2=1.005 $Y2=1.16
r54 19 21 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.815 $Y=1.66
+ $X2=0.815 $Y2=2.34
r55 17 29 5.0389 $w=3.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=1.325
+ $X2=0.815 $Y2=1.16
r56 17 19 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=1.325
+ $X2=0.815 $Y2=1.66
r57 13 29 5.0389 $w=3.4e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.775 $Y=0.995
+ $X2=0.815 $Y2=1.16
r58 13 15 16.7104 $w=2.98e-07 $l=4.35e-07 $layer=LI1_cond $X=0.775 $Y=0.995
+ $X2=0.775 $Y2=0.56
r59 4 39 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=1.485 $X2=1.81 $Y2=2.3
r60 4 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=1.485 $X2=1.81 $Y2=1.62
r61 3 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.695
+ $Y=1.485 $X2=0.84 $Y2=2.34
r62 3 19 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.695
+ $Y=1.485 $X2=0.84 $Y2=1.66
r63 2 27 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.235 $X2=1.79 $Y2=0.56
r64 1 15 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=0.655
+ $Y=0.235 $X2=0.84 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%A_657_325# 1 2 3 4 13 17 22 24 25 28 29 30
+ 32 35 39 43 45 48 50
c155 39 0 1.57566e-19 $X=6.79 $Y=0.545
c156 29 0 1.36535e-19 $X=6.415 $Y=2.36
r157 46 48 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.5 $Y=0.74
+ $X2=6.79 $Y2=0.74
r158 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.95 $Y=1.12
+ $X2=5.06 $Y2=1.12
r159 37 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.79 $Y=0.655
+ $X2=6.79 $Y2=0.74
r160 37 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.79 $Y=0.655
+ $X2=6.79 $Y2=0.545
r161 33 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.585 $Y=2.36
+ $X2=6.5 $Y2=2.36
r162 33 35 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=6.585 $Y=2.36
+ $X2=8.605 $Y2=2.36
r163 32 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=2.275 $X2=6.5
+ $Y2=2.36
r164 31 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=0.825
+ $X2=6.5 $Y2=0.74
r165 31 32 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=6.5 $Y=0.825
+ $X2=6.5 $Y2=2.275
r166 29 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.415 $Y=2.36
+ $X2=6.5 $Y2=2.36
r167 29 30 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=6.415 $Y=2.36
+ $X2=5.89 $Y2=2.36
r168 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.805 $Y=2.275
+ $X2=5.89 $Y2=2.36
r169 27 28 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.805 $Y=2.065
+ $X2=5.805 $Y2=2.275
r170 26 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=1.98
+ $X2=5.06 $Y2=1.98
r171 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.72 $Y=1.98
+ $X2=5.805 $Y2=2.065
r172 25 26 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.72 $Y=1.98
+ $X2=5.145 $Y2=1.98
r173 24 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=1.895
+ $X2=5.06 $Y2=1.98
r174 23 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=1.205
+ $X2=5.06 $Y2=1.12
r175 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.06 $Y=1.205
+ $X2=5.06 $Y2=1.895
r176 22 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=1.035
+ $X2=4.95 $Y2=1.12
r177 21 22 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.95 $Y=0.455
+ $X2=4.95 $Y2=1.035
r178 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.865 $Y=0.37
+ $X2=4.95 $Y2=0.455
r179 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.865 $Y=0.37
+ $X2=4.57 $Y2=0.37
r180 13 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.975 $Y=1.98
+ $X2=5.06 $Y2=1.98
r181 13 15 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=4.975 $Y=1.98
+ $X2=3.475 $Y2=1.98
r182 4 35 600 $w=1.7e-07 $l=8.21995e-07 $layer=licon1_PDIFF $count=1 $X=8.375
+ $Y=1.645 $X2=8.605 $Y2=2.36
r183 3 15 600 $w=1.7e-07 $l=4.39858e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.625 $X2=3.475 $Y2=1.98
r184 2 39 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.245 $X2=6.79 $Y2=0.545
r185 1 19 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=4.405
+ $Y=0.245 $X2=4.57 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%A_681_49# 1 2 3 4 13 16 17 19 21 24 26 27
+ 29 34 35 36 37 40 43
c135 29 0 1.24749e-19 $X=8.45 $Y=0.38
r136 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.17 $Y=1.53
+ $X2=7.17 $Y2=1.53
r137 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.72 $Y=1.53
+ $X2=4.72 $Y2=1.53
r138 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.865 $Y=1.53
+ $X2=4.72 $Y2=1.53
r139 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.025 $Y=1.53
+ $X2=7.17 $Y2=1.53
r140 36 37 2.67326 $w=1.4e-07 $l=2.16e-06 $layer=MET1_cond $X=7.025 $Y=1.53
+ $X2=4.865 $Y2=1.53
r141 32 34 10.6148 $w=2.78e-07 $l=2.15e-07 $layer=LI1_cond $X=3.54 $Y=0.765
+ $X2=3.755 $Y2=0.765
r142 27 35 11.5258 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=8.365 $Y=0.36
+ $X2=8.155 $Y2=0.36
r143 27 29 4.48918 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=8.365 $Y=0.36
+ $X2=8.45 $Y2=0.36
r144 26 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.645 $Y=0.34
+ $X2=8.155 $Y2=0.34
r145 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.56 $Y=0.425
+ $X2=7.645 $Y2=0.34
r146 23 24 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.56 $Y=0.425
+ $X2=7.56 $Y2=1.445
r147 22 44 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=7.23 $Y=1.53
+ $X2=7.022 $Y2=1.53
r148 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.475 $Y=1.53
+ $X2=7.56 $Y2=1.445
r149 21 22 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.475 $Y=1.53
+ $X2=7.23 $Y2=1.53
r150 17 44 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=7.022 $Y=1.615
+ $X2=7.022 $Y2=1.53
r151 17 19 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=7.022 $Y=1.615
+ $X2=7.022 $Y2=1.62
r152 16 40 8.59825 $w=3.35e-07 $l=1.55997e-07 $layer=LI1_cond $X=4.61 $Y=1.375
+ $X2=4.612 $Y2=1.53
r153 15 16 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.61 $Y=0.795
+ $X2=4.61 $Y2=1.375
r154 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.525 $Y=0.71
+ $X2=4.61 $Y2=0.795
r155 13 34 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.525 $Y=0.71
+ $X2=3.755 $Y2=0.71
r156 4 19 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=6.645
+ $Y=1.485 $X2=6.99 $Y2=1.62
r157 3 40 600 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=1.485 $X2=4.585 $Y2=1.61
r158 2 29 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=8.255
+ $Y=0.245 $X2=8.45 $Y2=0.38
r159 1 32 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.405
+ $Y=0.245 $X2=3.54 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%A_1490_297# 1 2 3 4 15 18 23 26 29 31 36
r66 34 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=10.11 $Y=0.42
+ $X2=10.24 $Y2=0.42
r67 28 29 17.0922 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=10.115 $Y=1.99
+ $X2=9.79 $Y2=1.99
r68 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=10.24 $Y=1.875
+ $X2=10.24 $Y2=1.99
r69 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.24 $Y=0.585
+ $X2=10.24 $Y2=0.42
r70 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=10.24 $Y=0.585
+ $X2=10.24 $Y2=1.875
r71 21 31 3.15669 $w=2.28e-07 $l=6.3e-08 $layer=LI1_cond $X=10.177 $Y=1.99
+ $X2=10.24 $Y2=1.99
r72 21 28 3.10659 $w=2.28e-07 $l=6.2e-08 $layer=LI1_cond $X=10.177 $Y=1.99
+ $X2=10.115 $Y2=1.99
r73 21 23 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=10.177 $Y=2.105
+ $X2=10.177 $Y2=2.3
r74 20 29 113.519 $w=1.68e-07 $l=1.74e-06 $layer=LI1_cond $X=8.05 $Y=2.02
+ $X2=9.79 $Y2=2.02
r75 18 20 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.985 $Y=2.02
+ $X2=8.05 $Y2=2.02
r76 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.9 $Y=1.935
+ $X2=7.985 $Y2=2.02
r77 13 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=7.9 $Y=1.935
+ $X2=7.9 $Y2=0.76
r78 4 28 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=9.965
+ $Y=1.485 $X2=10.115 $Y2=1.96
r79 4 23 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=9.965
+ $Y=1.485 $X2=10.115 $Y2=2.3
r80 3 20 600 $w=1.7e-07 $l=8.25227e-07 $layer=licon1_PDIFF $count=1 $X=7.45
+ $Y=1.485 $X2=8.05 $Y2=2.02
r81 2 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.975
+ $Y=0.235 $X2=10.11 $Y2=0.42
r82 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.245 $X2=7.9 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR3_4%VGND 1 2 3 4 5 18 22 24 28 32 36 39 40 41
+ 42 44 45 46 54 70 71 74 77
c127 71 0 1.70967e-19 $X=10.35 $Y=0
c128 36 0 3.96944e-20 $X=9.64 $Y=0.4
r129 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r130 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r131 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r132 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r133 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r134 65 68 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=9.43
+ $Y2=0
r135 65 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r136 64 67 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=9.43
+ $Y2=0
r137 64 65 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r138 62 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=0 $X2=5.29
+ $Y2=0
r139 62 64 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.375 $Y=0
+ $X2=5.75 $Y2=0
r140 61 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r141 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r142 58 61 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r143 58 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r144 57 60 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r145 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r146 55 74 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.195
+ $Y2=0
r147 55 57 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.345 $Y=0
+ $X2=2.53 $Y2=0
r148 54 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=0 $X2=5.29
+ $Y2=0
r149 54 60 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.205 $Y=0
+ $X2=4.83 $Y2=0
r150 53 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r151 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r152 46 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r153 46 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r154 44 67 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.555 $Y=0
+ $X2=9.43 $Y2=0
r155 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.555 $Y=0 $X2=9.64
+ $Y2=0
r156 43 70 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=9.725 $Y=0
+ $X2=10.35 $Y2=0
r157 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.725 $Y=0 $X2=9.64
+ $Y2=0
r158 41 52 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.15
+ $Y2=0
r159 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.31
+ $Y2=0
r160 39 49 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.23
+ $Y2=0
r161 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.37
+ $Y2=0
r162 38 52 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.455 $Y=0
+ $X2=1.15 $Y2=0
r163 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.37
+ $Y2=0
r164 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.64 $Y=0.085
+ $X2=9.64 $Y2=0
r165 34 36 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.64 $Y=0.085
+ $X2=9.64 $Y2=0.4
r166 30 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.29 $Y=0.085
+ $X2=5.29 $Y2=0
r167 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.29 $Y=0.085
+ $X2=5.29 $Y2=0.36
r168 26 74 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0
r169 26 28 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0.36
r170 25 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.31
+ $Y2=0
r171 24 74 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=2.195
+ $Y2=0
r172 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=1.395 $Y2=0
r173 20 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=0.085
+ $X2=1.31 $Y2=0
r174 20 22 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.31 $Y=0.085
+ $X2=1.31 $Y2=0.56
r175 16 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.37 $Y2=0
r176 16 18 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.37 $Y2=0.56
r177 5 36 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=9.505
+ $Y=0.235 $X2=9.64 $Y2=0.4
r178 4 32 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=5.135
+ $Y=0.235 $X2=5.29 $Y2=0.36
r179 3 28 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.235 $X2=2.26 $Y2=0.36
r180 2 22 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.31 $Y2=0.56
r181 1 18 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.56
.ends

