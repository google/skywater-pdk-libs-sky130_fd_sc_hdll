* File: sky130_fd_sc_hdll__a21o_8.spice
* Created: Wed Sep  2 08:17:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21o_8.pex.spice"
.subckt sky130_fd_sc_hdll__a21o_8  VNB VPB A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1000 A_297_47# N_A2_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65 AD=0.0845
+ AS=0.169 PD=0.91 PS=1.82 NRD=13.836 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75006.7
+ A=0.0975 P=1.6 MULT=1
MM1008 N_A_213_47#_M1008_d N_A1_M1008_g A_297_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.0845 PD=0.92 PS=0.91 NRD=0 NRS=13.836 M=1 R=4.33333 SA=75000.6
+ SB=75006.3 A=0.0975 P=1.6 MULT=1
MM1004 N_A_213_47#_M1008_d N_A1_M1004_g A_131_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.0845 PD=0.92 PS=0.91 NRD=0 NRS=13.836 M=1 R=4.33333 SA=75001
+ SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1014 A_131_47# N_A2_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65 AD=0.0845
+ AS=0.13975 PD=0.91 PS=1.08 NRD=13.836 NRS=13.836 M=1 R=4.33333 SA=75001.4
+ SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1016 N_A_213_47#_M1016_d N_B1_M1016_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.13975 PD=0.92 PS=1.08 NRD=0 NRS=13.836 M=1 R=4.33333 SA=75002
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1023 N_A_213_47#_M1016_d N_B1_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.28925 PD=0.92 PS=1.54 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.4
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_213_47#_M1001_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.28925 PD=0.92 PS=1.54 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75003.5 SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1002 N_X_M1001_d N_A_213_47#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.9
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_213_47#_M1006_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.4
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1006_d N_A_213_47#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.8
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1019 N_X_M1019_d N_A_213_47#_M1019_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.3
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1020 N_X_M1019_d N_A_213_47#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.8
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1022 N_X_M1022_d N_A_213_47#_M1022_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.3
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1026 N_X_M1022_d N_A_213_47#_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_A2_M1011_g N_A_27_297#_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1003 N_A_27_297#_M1003_d N_A1_M1003_g N_VPWR_M1011_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1024 N_A_27_297#_M1003_d N_A1_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1024_s N_A2_M1017_g N_A_27_297#_M1017_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1017_s N_B1_M1009_g N_A_213_47#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1012 N_A_27_297#_M1012_d N_B1_M1012_g N_A_213_47#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_X_M1005_d N_A_213_47#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1007 N_X_M1005_d N_A_213_47#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1013 N_X_M1013_d N_A_213_47#_M1013_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1015 N_X_M1013_d N_A_213_47#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1018 N_X_M1018_d N_A_213_47#_M1018_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1021 N_X_M1018_d N_A_213_47#_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1025 N_X_M1025_d N_A_213_47#_M1025_g N_VPWR_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1027 N_X_M1025_d N_A_213_47#_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=13.161 P=19.61
c_52 VNB 0 1.34369e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hdll__a21o_8.pxi.spice"
*
.ends
*
*
