* File: sky130_fd_sc_hdll__clkbuf_12.pex.spice
* Created: Thu Aug 27 19:01:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_12%A 1 3 6 10 12 14 15 17 20 24 26 28 29 40
c75 40 0 1.95681e-20 $X=1.88 $Y=1.155
c76 26 0 1.38915e-19 $X=1.905 $Y=1.41
r77 40 41 2.5803 $w=4.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.155
+ $X2=1.905 $Y2=1.155
r78 39 40 43.349 $w=4.67e-07 $l=4.2e-07 $layer=POLY_cond $X=1.46 $Y=1.155
+ $X2=1.88 $Y2=1.155
r79 38 39 2.5803 $w=4.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.155
+ $X2=1.46 $Y2=1.155
r80 36 38 28.8994 $w=4.67e-07 $l=2.8e-07 $layer=POLY_cond $X=1.155 $Y=1.155
+ $X2=1.435 $Y2=1.155
r81 34 36 19.6103 $w=4.67e-07 $l=1.9e-07 $layer=POLY_cond $X=0.965 $Y=1.155
+ $X2=1.155 $Y2=1.155
r82 33 34 2.5803 $w=4.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.155
+ $X2=0.965 $Y2=1.155
r83 32 33 43.349 $w=4.67e-07 $l=4.2e-07 $layer=POLY_cond $X=0.52 $Y=1.155
+ $X2=0.94 $Y2=1.155
r84 31 32 2.5803 $w=4.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.155
+ $X2=0.52 $Y2=1.155
r85 29 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.155
+ $Y=1.16 $X2=1.155 $Y2=1.16
r86 26 41 25.192 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.155
r87 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r88 22 40 29.6916 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.88 $Y=0.9
+ $X2=1.88 $Y2=1.155
r89 22 24 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.88 $Y=0.9
+ $X2=1.88 $Y2=0.445
r90 18 39 29.6916 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.46 $Y=0.9
+ $X2=1.46 $Y2=1.155
r91 18 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.46 $Y=0.9
+ $X2=1.46 $Y2=0.445
r92 15 38 25.192 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.155
r93 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r94 12 34 25.192 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.155
r95 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r96 8 33 29.6916 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.94 $Y=0.9 $X2=0.94
+ $Y2=1.155
r97 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.94 $Y=0.9 $X2=0.94
+ $Y2=0.445
r98 4 32 29.6916 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.52 $Y=0.9 $X2=0.52
+ $Y2=1.155
r99 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=0.9 $X2=0.52
+ $Y2=0.445
r100 1 31 25.192 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.155
r101 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_12%A_117_297# 1 2 3 4 13 15 18 22 24 26 27
+ 29 32 36 38 40 41 43 46 50 52 54 55 57 60 64 66 68 69 71 74 78 80 82 83 85 88
+ 92 94 96 97 99 103 105 106 107 111 114 116 119 126 131 132 134 159
c271 134 0 1.41094e-19 $X=1.67 $Y=1.62
c272 131 0 1.68289e-20 $X=1.67 $Y=0.81
c273 106 0 1.68289e-20 $X=0.865 $Y=0.81
c274 94 0 8.80852e-20 $X=7.545 $Y=1.41
r275 159 160 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=7.52 $Y=1.18
+ $X2=7.545 $Y2=1.18
r276 158 159 49.1359 $w=4.12e-07 $l=4.2e-07 $layer=POLY_cond $X=7.1 $Y=1.18
+ $X2=7.52 $Y2=1.18
r277 157 158 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=7.075 $Y=1.18
+ $X2=7.1 $Y2=1.18
r278 156 157 54.9854 $w=4.12e-07 $l=4.7e-07 $layer=POLY_cond $X=6.605 $Y=1.18
+ $X2=7.075 $Y2=1.18
r279 155 156 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=6.58 $Y=1.18
+ $X2=6.605 $Y2=1.18
r280 152 153 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=6.135 $Y=1.18
+ $X2=6.16 $Y2=1.18
r281 151 152 54.9854 $w=4.12e-07 $l=4.7e-07 $layer=POLY_cond $X=5.665 $Y=1.18
+ $X2=6.135 $Y2=1.18
r282 150 151 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=5.64 $Y=1.18
+ $X2=5.665 $Y2=1.18
r283 149 150 49.1359 $w=4.12e-07 $l=4.2e-07 $layer=POLY_cond $X=5.22 $Y=1.18
+ $X2=5.64 $Y2=1.18
r284 148 149 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=5.195 $Y=1.18
+ $X2=5.22 $Y2=1.18
r285 147 148 54.9854 $w=4.12e-07 $l=4.7e-07 $layer=POLY_cond $X=4.725 $Y=1.18
+ $X2=5.195 $Y2=1.18
r286 146 147 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.18
+ $X2=4.725 $Y2=1.18
r287 145 146 49.1359 $w=4.12e-07 $l=4.2e-07 $layer=POLY_cond $X=4.28 $Y=1.18
+ $X2=4.7 $Y2=1.18
r288 144 145 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=4.255 $Y=1.18
+ $X2=4.28 $Y2=1.18
r289 143 144 54.9854 $w=4.12e-07 $l=4.7e-07 $layer=POLY_cond $X=3.785 $Y=1.18
+ $X2=4.255 $Y2=1.18
r290 142 143 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.18
+ $X2=3.785 $Y2=1.18
r291 141 142 49.1359 $w=4.12e-07 $l=4.2e-07 $layer=POLY_cond $X=3.34 $Y=1.18
+ $X2=3.76 $Y2=1.18
r292 140 141 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=3.315 $Y=1.18
+ $X2=3.34 $Y2=1.18
r293 139 140 54.9854 $w=4.12e-07 $l=4.7e-07 $layer=POLY_cond $X=2.845 $Y=1.18
+ $X2=3.315 $Y2=1.18
r294 138 139 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.18
+ $X2=2.845 $Y2=1.18
r295 135 136 2.92476 $w=4.12e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.18
+ $X2=2.4 $Y2=1.18
r296 127 155 7.01942 $w=4.12e-07 $l=6e-08 $layer=POLY_cond $X=6.52 $Y=1.18
+ $X2=6.58 $Y2=1.18
r297 127 153 42.1165 $w=4.12e-07 $l=3.6e-07 $layer=POLY_cond $X=6.52 $Y=1.18
+ $X2=6.16 $Y2=1.18
r298 126 127 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=6.52
+ $Y=1.16 $X2=6.52 $Y2=1.16
r299 124 138 44.4563 $w=4.12e-07 $l=3.8e-07 $layer=POLY_cond $X=2.44 $Y=1.18
+ $X2=2.82 $Y2=1.18
r300 124 136 4.67961 $w=4.12e-07 $l=4e-08 $layer=POLY_cond $X=2.44 $Y=1.18
+ $X2=2.4 $Y2=1.18
r301 123 126 204.433 $w=2.28e-07 $l=4.08e-06 $layer=LI1_cond $X=2.44 $Y=1.19
+ $X2=6.52 $Y2=1.19
r302 123 124 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=2.44
+ $Y=1.16 $X2=2.44 $Y2=1.16
r303 121 132 1.92582 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=1.19
+ $X2=1.67 $Y2=1.19
r304 121 123 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.805 $Y=1.19
+ $X2=2.44 $Y2=1.19
r305 117 134 3.82129 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.57
r306 117 119 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=2.3
r307 116 134 3.82129 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.67 $Y=1.475
+ $X2=1.67 $Y2=1.57
r308 115 132 4.51169 $w=2.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.67 $Y=1.305
+ $X2=1.67 $Y2=1.19
r309 115 116 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.67 $Y=1.305
+ $X2=1.67 $Y2=1.475
r310 114 132 4.51169 $w=2.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.67 $Y=1.075
+ $X2=1.67 $Y2=1.19
r311 113 131 3.82129 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.67 $Y=0.905
+ $X2=1.67 $Y2=0.81
r312 113 114 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.67 $Y=0.905
+ $X2=1.67 $Y2=1.075
r313 109 131 3.82129 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.67 $Y=0.715
+ $X2=1.67 $Y2=0.81
r314 109 111 11.5244 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.67 $Y=0.715
+ $X2=1.67 $Y2=0.445
r315 108 130 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.57
+ $X2=0.73 $Y2=1.57
r316 107 134 2.63355 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=1.57
+ $X2=1.67 $Y2=1.57
r317 107 108 37.3589 $w=1.88e-07 $l=6.4e-07 $layer=LI1_cond $X=1.535 $Y=1.57
+ $X2=0.895 $Y2=1.57
r318 105 131 2.63355 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=0.81
+ $X2=1.67 $Y2=0.81
r319 105 106 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=0.81
+ $X2=0.865 $Y2=0.81
r320 101 106 7.08811 $w=1.9e-07 $l=1.7621e-07 $layer=LI1_cond $X=0.73 $Y=0.715
+ $X2=0.865 $Y2=0.81
r321 101 103 11.5244 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.73 $Y=0.715
+ $X2=0.73 $Y2=0.445
r322 97 130 2.73294 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.57
r323 97 99 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.3
r324 94 160 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.18
r325 94 96 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.985
r326 90 159 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=7.52 $Y=0.95
+ $X2=7.52 $Y2=1.18
r327 90 92 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.52 $Y=0.95
+ $X2=7.52 $Y2=0.445
r328 86 158 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=7.1 $Y=0.95
+ $X2=7.1 $Y2=1.18
r329 86 88 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.1 $Y=0.95
+ $X2=7.1 $Y2=0.445
r330 83 157 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.18
r331 83 85 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.985
r332 80 156 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.18
r333 80 82 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.985
r334 76 155 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.58 $Y=0.95
+ $X2=6.58 $Y2=1.18
r335 76 78 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.58 $Y=0.95
+ $X2=6.58 $Y2=0.445
r336 72 153 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.16 $Y=0.95
+ $X2=6.16 $Y2=1.18
r337 72 74 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.16 $Y=0.95
+ $X2=6.16 $Y2=0.445
r338 69 152 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.18
r339 69 71 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.985
r340 66 151 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.18
r341 66 68 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r342 62 150 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.64 $Y=0.95
+ $X2=5.64 $Y2=1.18
r343 62 64 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.64 $Y=0.95
+ $X2=5.64 $Y2=0.445
r344 58 149 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.22 $Y=0.95
+ $X2=5.22 $Y2=1.18
r345 58 60 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.22 $Y=0.95
+ $X2=5.22 $Y2=0.445
r346 55 148 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.18
r347 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r348 52 147 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.18
r349 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r350 48 146 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.7 $Y=0.95
+ $X2=4.7 $Y2=1.18
r351 48 50 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.7 $Y=0.95
+ $X2=4.7 $Y2=0.445
r352 44 145 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.28 $Y=0.95
+ $X2=4.28 $Y2=1.18
r353 44 46 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.28 $Y=0.95
+ $X2=4.28 $Y2=0.445
r354 41 144 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.18
r355 41 43 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r356 38 143 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.18
r357 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r358 34 142 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.76 $Y=0.95
+ $X2=3.76 $Y2=1.18
r359 34 36 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.76 $Y=0.95
+ $X2=3.76 $Y2=0.445
r360 30 141 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.34 $Y=0.95
+ $X2=3.34 $Y2=1.18
r361 30 32 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.34 $Y=0.95
+ $X2=3.34 $Y2=0.445
r362 27 140 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.18
r363 27 29 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r364 24 139 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.18
r365 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r366 20 138 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.82 $Y=0.95
+ $X2=2.82 $Y2=1.18
r367 20 22 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.82 $Y=0.95
+ $X2=2.82 $Y2=0.445
r368 16 136 26.5862 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.4 $Y=0.95
+ $X2=2.4 $Y2=1.18
r369 16 18 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.4 $Y=0.95
+ $X2=2.4 $Y2=0.445
r370 13 135 22.168 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.18
r371 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r372 4 134 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.62
r373 4 119 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.3
r374 3 130 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.62
r375 3 99 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.3
r376 2 111 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.445
r377 1 103 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_12%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 40 44 48
+ 50 54 56 60 62 66 70 74 79 80 82 83 84 86 91 104 105 111 114 117 120 123 126
r134 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r135 124 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r136 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r137 121 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r138 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r139 118 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r140 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r141 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r142 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r143 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r144 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r145 102 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r146 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r147 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r148 99 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.75 $Y2=2.72
r149 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r150 96 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=2.72
+ $X2=5.9 $Y2=2.72
r151 96 98 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.065 $Y=2.72
+ $X2=6.67 $Y2=2.72
r152 95 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r153 95 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r154 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r155 92 111 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.2 $Y2=2.72
r156 92 94 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.61 $Y2=2.72
r157 91 114 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=2.125 $Y2=2.72
r158 91 94 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=1.61 $Y2=2.72
r159 90 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r160 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r161 87 108 4.49698 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r162 87 89 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r163 86 111 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.2 $Y2=2.72
r164 86 89 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r165 84 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r166 84 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r167 82 101 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.615 $Y=2.72
+ $X2=7.59 $Y2=2.72
r168 82 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.615 $Y=2.72
+ $X2=7.78 $Y2=2.72
r169 81 104 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.945 $Y=2.72
+ $X2=8.05 $Y2=2.72
r170 81 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.945 $Y=2.72
+ $X2=7.78 $Y2=2.72
r171 79 98 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.67 $Y2=2.72
r172 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.84 $Y2=2.72
r173 78 101 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=7.005 $Y=2.72
+ $X2=7.59 $Y2=2.72
r174 78 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=2.72
+ $X2=6.84 $Y2=2.72
r175 74 77 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.78 $Y=1.63
+ $X2=7.78 $Y2=2.31
r176 72 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=2.72
r177 72 77 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=2.31
r178 68 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2.72
r179 68 70 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=1.96
r180 64 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2.72
r181 64 66 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=1.96
r182 63 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=2.72
+ $X2=4.96 $Y2=2.72
r183 62 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.9 $Y2=2.72
r184 62 63 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.125 $Y2=2.72
r185 58 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2.72
r186 58 60 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=1.96
r187 57 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.02 $Y2=2.72
r188 56 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.96 $Y2=2.72
r189 56 57 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.185 $Y2=2.72
r190 52 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r191 52 54 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=1.96
r192 51 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.08 $Y2=2.72
r193 50 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=4.02 $Y2=2.72
r194 50 51 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=3.245 $Y2=2.72
r195 46 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r196 46 48 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=1.96
r197 45 114 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.125 $Y2=2.72
r198 44 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=3.08 $Y2=2.72
r199 44 45 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=2.275 $Y2=2.72
r200 40 43 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=2.125 $Y=1.64
+ $X2=2.125 $Y2=2.32
r201 38 114 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=2.635
+ $X2=2.125 $Y2=2.72
r202 38 43 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=2.125 $Y=2.635
+ $X2=2.125 $Y2=2.32
r203 34 111 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r204 34 36 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r205 30 33 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=0.245 $Y=1.66
+ $X2=0.245 $Y2=2.34
r206 28 108 3.0207 $w=3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.197 $Y2=2.72
r207 28 33 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.245 $Y2=2.34
r208 9 77 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=2.31
r209 9 74 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=1.63
r210 8 70 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=1.96
r211 7 66 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=1.96
r212 6 60 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.96
r213 5 54 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.96
r214 4 48 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.96
r215 3 43 400 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.32
r216 3 40 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.64
r217 2 36 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r218 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r219 1 30 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_12%X 1 2 3 4 5 6 7 8 9 10 11 12 37 39 43 45
+ 46 47 51 55 57 59 63 67 69 71 75 79 81 83 87 91 93 95 99 103 107 109 110 112
+ 113 115 116 118 120 123 124
c197 123 0 1.41094e-19 $X=7.31 $Y=1.62
c198 46 0 1.95681e-20 $X=2.745 $Y=0.81
c199 37 0 5.08297e-20 $X=2.595 $Y=1.665
r200 121 124 7.0285 $w=4.83e-07 $l=2.85e-07 $layer=LI1_cond $X=7.202 $Y=1.475
+ $X2=7.202 $Y2=1.19
r201 121 123 2.82679 $w=3.77e-07 $l=9.5e-08 $layer=LI1_cond $X=7.202 $Y=1.475
+ $X2=7.202 $Y2=1.57
r202 119 124 7.0285 $w=4.83e-07 $l=2.85e-07 $layer=LI1_cond $X=7.202 $Y=0.905
+ $X2=7.202 $Y2=1.19
r203 119 120 2.82679 $w=3.77e-07 $l=9.5e-08 $layer=LI1_cond $X=7.202 $Y=0.905
+ $X2=7.202 $Y2=0.81
r204 101 123 2.82679 $w=3.77e-07 $l=1.48068e-07 $layer=LI1_cond $X=7.31 $Y=1.665
+ $X2=7.202 $Y2=1.57
r205 101 103 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.31 $Y=1.665
+ $X2=7.31 $Y2=2.3
r206 97 120 2.82679 $w=3.77e-07 $l=1.48068e-07 $layer=LI1_cond $X=7.31 $Y=0.715
+ $X2=7.202 $Y2=0.81
r207 97 99 11.5244 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.31 $Y=0.715
+ $X2=7.31 $Y2=0.445
r208 96 118 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=6.505 $Y=1.57
+ $X2=6.37 $Y2=1.57
r209 95 123 3.89798 $w=1.9e-07 $l=2.42e-07 $layer=LI1_cond $X=6.96 $Y=1.57
+ $X2=7.202 $Y2=1.57
r210 95 96 26.5598 $w=1.88e-07 $l=4.55e-07 $layer=LI1_cond $X=6.96 $Y=1.57
+ $X2=6.505 $Y2=1.57
r211 94 116 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=6.505 $Y=0.81
+ $X2=6.37 $Y2=0.81
r212 93 120 3.89798 $w=1.9e-07 $l=2.42e-07 $layer=LI1_cond $X=6.96 $Y=0.81
+ $X2=7.202 $Y2=0.81
r213 93 94 26.5598 $w=1.88e-07 $l=4.55e-07 $layer=LI1_cond $X=6.96 $Y=0.81
+ $X2=6.505 $Y2=0.81
r214 89 118 0.11353 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.37 $Y=1.665
+ $X2=6.37 $Y2=1.57
r215 89 91 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.37 $Y=1.665
+ $X2=6.37 $Y2=2.3
r216 85 116 0.11353 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.37 $Y=0.715
+ $X2=6.37 $Y2=0.81
r217 85 87 11.5244 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.37 $Y=0.715
+ $X2=6.37 $Y2=0.445
r218 84 115 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=5.565 $Y=1.57
+ $X2=5.43 $Y2=1.57
r219 83 118 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=6.235 $Y=1.57
+ $X2=6.37 $Y2=1.57
r220 83 84 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=6.235 $Y=1.57
+ $X2=5.565 $Y2=1.57
r221 82 113 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=5.565 $Y=0.81
+ $X2=5.43 $Y2=0.81
r222 81 116 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=6.235 $Y=0.81
+ $X2=6.37 $Y2=0.81
r223 81 82 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=6.235 $Y=0.81
+ $X2=5.565 $Y2=0.81
r224 77 115 0.11353 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.43 $Y=1.665
+ $X2=5.43 $Y2=1.57
r225 77 79 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.43 $Y=1.665
+ $X2=5.43 $Y2=2.3
r226 73 113 0.11353 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.43 $Y=0.715
+ $X2=5.43 $Y2=0.81
r227 73 75 11.5244 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.43 $Y=0.715
+ $X2=5.43 $Y2=0.445
r228 72 112 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=1.57
+ $X2=4.49 $Y2=1.57
r229 71 115 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=5.295 $Y=1.57
+ $X2=5.43 $Y2=1.57
r230 71 72 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=5.295 $Y=1.57
+ $X2=4.625 $Y2=1.57
r231 70 110 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=0.81
+ $X2=4.49 $Y2=0.81
r232 69 113 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=5.295 $Y=0.81
+ $X2=5.43 $Y2=0.81
r233 69 70 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=5.295 $Y=0.81
+ $X2=4.625 $Y2=0.81
r234 65 112 0.11353 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.49 $Y=1.665
+ $X2=4.49 $Y2=1.57
r235 65 67 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.49 $Y=1.665
+ $X2=4.49 $Y2=2.3
r236 61 110 0.11353 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.49 $Y=0.715
+ $X2=4.49 $Y2=0.81
r237 61 63 11.5244 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.49 $Y=0.715
+ $X2=4.49 $Y2=0.445
r238 60 109 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=1.57
+ $X2=3.55 $Y2=1.57
r239 59 112 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=1.57
+ $X2=4.49 $Y2=1.57
r240 59 60 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=1.57
+ $X2=3.685 $Y2=1.57
r241 58 107 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=0.81
+ $X2=3.55 $Y2=0.81
r242 57 110 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=0.81
+ $X2=4.49 $Y2=0.81
r243 57 58 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=0.81
+ $X2=3.685 $Y2=0.81
r244 53 109 0.11353 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=1.57
r245 53 55 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=2.3
r246 49 107 0.11353 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.55 $Y=0.715
+ $X2=3.55 $Y2=0.81
r247 49 51 11.5244 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.55 $Y=0.715
+ $X2=3.55 $Y2=0.445
r248 48 106 4.45288 $w=1.9e-07 $l=1.5e-07 $layer=LI1_cond $X=2.745 $Y=1.57
+ $X2=2.595 $Y2=1.57
r249 47 109 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=1.57
+ $X2=3.55 $Y2=1.57
r250 47 48 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=1.57
+ $X2=2.745 $Y2=1.57
r251 45 107 6.84645 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=0.81
+ $X2=3.55 $Y2=0.81
r252 45 46 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=0.81
+ $X2=2.745 $Y2=0.81
r253 41 46 7.08811 $w=1.9e-07 $l=1.7621e-07 $layer=LI1_cond $X=2.61 $Y=0.715
+ $X2=2.745 $Y2=0.81
r254 41 43 11.5244 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.61 $Y=0.715
+ $X2=2.61 $Y2=0.445
r255 37 106 2.82016 $w=3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.595 $Y=1.665
+ $X2=2.595 $Y2=1.57
r256 37 39 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=2.595 $Y=1.665
+ $X2=2.595 $Y2=2.3
r257 12 123 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=1.62
r258 12 103 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=2.3
r259 11 118 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=1.62
r260 11 91 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=2.3
r261 10 115 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.62
r262 10 79 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.3
r263 9 112 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.62
r264 9 67 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2.3
r265 8 109 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.62
r266 8 55 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.3
r267 7 106 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r268 7 39 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.3
r269 6 99 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=7.175
+ $Y=0.235 $X2=7.31 $Y2=0.445
r270 5 87 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.235 $X2=6.37 $Y2=0.445
r271 4 75 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.235 $X2=5.43 $Y2=0.445
r272 3 63 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.49 $Y2=0.445
r273 2 51 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.55 $Y2=0.445
r274 1 43 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_12%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 40 44
+ 46 50 52 56 58 62 66 70 73 74 76 77 78 80 85 98 99 105 108 111 114 117 120
r128 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r129 118 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r130 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r131 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r132 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r133 112 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r134 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r135 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r136 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r137 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r138 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r139 96 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.05
+ $Y2=0
r140 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r141 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r142 93 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=5.75 $Y2=0
r143 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r144 90 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=0 $X2=5.9
+ $Y2=0
r145 90 92 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.065 $Y=0
+ $X2=6.67 $Y2=0
r146 89 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.07 $Y2=0
r147 89 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=1.15 $Y2=0
r148 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r149 86 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.2
+ $Y2=0
r150 86 88 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r151 85 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=2.14 $Y2=0
r152 85 88 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=1.61 $Y2=0
r153 84 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.15 $Y2=0
r154 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r155 81 102 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r156 81 83 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r157 80 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r158 80 83 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r159 78 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r160 78 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r161 76 95 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.59
+ $Y2=0
r162 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.78
+ $Y2=0
r163 75 98 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.945 $Y=0
+ $X2=8.05 $Y2=0
r164 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.945 $Y=0 $X2=7.78
+ $Y2=0
r165 73 92 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.67
+ $Y2=0
r166 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.84
+ $Y2=0
r167 72 95 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=7.59 $Y2=0
r168 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=0 $X2=6.84
+ $Y2=0
r169 68 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.78 $Y=0.085
+ $X2=7.78 $Y2=0
r170 68 70 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=7.78 $Y=0.085
+ $X2=7.78 $Y2=0.445
r171 64 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0
r172 64 66 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0.445
r173 60 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0.085
+ $X2=5.9 $Y2=0
r174 60 62 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.9 $Y=0.085
+ $X2=5.9 $Y2=0.445
r175 59 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0
+ $X2=4.96 $Y2=0
r176 58 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.9
+ $Y2=0
r177 58 59 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=5.125 $Y2=0
r178 54 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r179 54 56 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.445
r180 53 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=4.02 $Y2=0
r181 52 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0
+ $X2=4.96 $Y2=0
r182 52 53 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.795 $Y=0
+ $X2=4.185 $Y2=0
r183 48 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r184 48 50 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.445
r185 47 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0
+ $X2=3.08 $Y2=0
r186 46 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0
+ $X2=4.02 $Y2=0
r187 46 47 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=0
+ $X2=3.245 $Y2=0
r188 42 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0
r189 42 44 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.445
r190 41 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.14 $Y2=0
r191 40 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0
+ $X2=3.08 $Y2=0
r192 40 41 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=0
+ $X2=2.305 $Y2=0
r193 36 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r194 36 38 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.445
r195 32 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0
r196 32 34 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.445
r197 28 102 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r198 28 30 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.445
r199 9 70 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=7.595
+ $Y=0.235 $X2=7.78 $Y2=0.445
r200 8 66 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.235 $X2=6.84 $Y2=0.445
r201 7 62 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=5.715
+ $Y=0.235 $X2=5.9 $Y2=0.445
r202 6 56 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.445
r203 5 50 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.445
r204 4 44 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.445
r205 3 38 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.445
r206 2 34 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.445
r207 1 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

