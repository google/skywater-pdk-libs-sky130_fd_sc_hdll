# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__bufbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__bufbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA  1.409500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  2.044400 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.480000 0.260000 3.860000 0.735000 ;
        RECT 3.480000 0.735000 7.240000 0.905000 ;
        RECT 3.480000 1.445000 7.240000 1.615000 ;
        RECT 3.480000 1.615000 3.860000 2.465000 ;
        RECT 4.420000 0.260000 4.800000 0.735000 ;
        RECT 4.420000 1.615000 4.800000 2.465000 ;
        RECT 5.360000 0.260000 5.740000 0.735000 ;
        RECT 5.360000 1.615000 5.740000 2.465000 ;
        RECT 6.300000 0.260000 6.680000 0.735000 ;
        RECT 6.300000 1.615000 6.680000 2.465000 ;
        RECT 6.860000 0.905000 7.240000 1.445000 ;
    END
  END X
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.260000 0.425000 0.735000 ;
      RECT 0.095000  0.735000 0.830000 0.905000 ;
      RECT 0.095000  1.445000 0.830000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.160000 ;
      RECT 0.645000  0.085000 0.815000 0.565000 ;
      RECT 0.645000  1.785000 0.815000 2.635000 ;
      RECT 0.660000  0.905000 0.830000 0.995000 ;
      RECT 0.660000  0.995000 1.140000 1.325000 ;
      RECT 0.660000  1.325000 0.830000 1.445000 ;
      RECT 1.050000  0.260000 1.480000 0.825000 ;
      RECT 1.050000  1.545000 1.480000 2.465000 ;
      RECT 1.310000  0.825000 1.480000 1.075000 ;
      RECT 1.310000  1.075000 2.920000 1.275000 ;
      RECT 1.310000  1.275000 1.480000 1.545000 ;
      RECT 1.650000  0.260000 1.980000 0.735000 ;
      RECT 1.650000  0.735000 3.310000 0.905000 ;
      RECT 1.650000  1.445000 3.310000 1.615000 ;
      RECT 1.650000  1.615000 1.980000 2.465000 ;
      RECT 2.200000  0.085000 2.370000 0.565000 ;
      RECT 2.200000  1.785000 2.370000 2.635000 ;
      RECT 2.540000  0.260000 2.920000 0.735000 ;
      RECT 2.540000  1.615000 2.920000 2.465000 ;
      RECT 3.140000  0.085000 3.310000 0.565000 ;
      RECT 3.140000  0.905000 3.310000 1.075000 ;
      RECT 3.140000  1.075000 5.910000 1.275000 ;
      RECT 3.140000  1.275000 3.310000 1.445000 ;
      RECT 3.140000  1.785000 3.310000 2.635000 ;
      RECT 4.080000  0.085000 4.250000 0.565000 ;
      RECT 4.080000  1.835000 4.250000 2.635000 ;
      RECT 5.020000  0.085000 5.190000 0.565000 ;
      RECT 5.020000  1.835000 5.190000 2.635000 ;
      RECT 5.960000  0.085000 6.130000 0.565000 ;
      RECT 5.960000  1.835000 6.130000 2.635000 ;
      RECT 6.900000  0.085000 7.070000 0.565000 ;
      RECT 6.900000  1.835000 7.070000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufbuf_8
END LIBRARY
