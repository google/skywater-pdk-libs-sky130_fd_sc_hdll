* File: sky130_fd_sc_hdll__einvp_4.pxi.spice
* Created: Wed Sep  2 08:31:47 2020
* 
x_PM_SKY130_FD_SC_HDLL__EINVP_4%TE N_TE_c_84_n N_TE_M1004_g N_TE_c_85_n
+ N_TE_M1013_g N_TE_c_86_n N_TE_c_87_n N_TE_M1000_g N_TE_c_88_n N_TE_c_89_n
+ N_TE_M1006_g N_TE_c_90_n N_TE_c_91_n N_TE_M1007_g N_TE_c_92_n N_TE_c_93_n
+ N_TE_M1010_g N_TE_c_94_n N_TE_c_95_n N_TE_c_96_n TE TE
+ PM_SKY130_FD_SC_HDLL__EINVP_4%TE
x_PM_SKY130_FD_SC_HDLL__EINVP_4%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1004_s
+ N_A_27_47#_c_171_n N_A_27_47#_M1003_g N_A_27_47#_c_172_n N_A_27_47#_c_173_n
+ N_A_27_47#_c_174_n N_A_27_47#_M1011_g N_A_27_47#_c_175_n N_A_27_47#_c_176_n
+ N_A_27_47#_M1015_g N_A_27_47#_c_177_n N_A_27_47#_c_178_n N_A_27_47#_M1016_g
+ N_A_27_47#_c_179_n N_A_27_47#_c_180_n N_A_27_47#_c_181_n N_A_27_47#_c_166_n
+ N_A_27_47#_c_182_n N_A_27_47#_c_167_n N_A_27_47#_c_168_n N_A_27_47#_c_183_n
+ N_A_27_47#_c_169_n N_A_27_47#_c_170_n N_A_27_47#_c_212_n
+ PM_SKY130_FD_SC_HDLL__EINVP_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EINVP_4%A N_A_c_281_n N_A_M1001_g N_A_c_287_n
+ N_A_M1005_g N_A_c_282_n N_A_M1002_g N_A_c_288_n N_A_M1012_g N_A_M1008_g
+ N_A_c_289_n N_A_M1014_g N_A_M1009_g N_A_c_290_n N_A_M1017_g A A A N_A_c_285_n
+ A A PM_SKY130_FD_SC_HDLL__EINVP_4%A
x_PM_SKY130_FD_SC_HDLL__EINVP_4%VPWR N_VPWR_M1004_d N_VPWR_M1003_d
+ N_VPWR_M1015_d N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_358_n
+ N_VPWR_c_359_n N_VPWR_c_360_n VPWR N_VPWR_c_361_n N_VPWR_c_362_n
+ N_VPWR_c_354_n N_VPWR_c_364_n N_VPWR_c_365_n
+ PM_SKY130_FD_SC_HDLL__EINVP_4%VPWR
x_PM_SKY130_FD_SC_HDLL__EINVP_4%A_235_309# N_A_235_309#_M1003_s
+ N_A_235_309#_M1011_s N_A_235_309#_M1016_s N_A_235_309#_M1012_d
+ N_A_235_309#_M1017_d N_A_235_309#_c_432_n N_A_235_309#_c_433_n
+ N_A_235_309#_c_429_n N_A_235_309#_c_444_n N_A_235_309#_c_446_n
+ N_A_235_309#_c_450_n N_A_235_309#_c_455_n N_A_235_309#_c_482_n
+ N_A_235_309#_c_492_p N_A_235_309#_c_430_n N_A_235_309#_c_431_n
+ N_A_235_309#_c_451_n N_A_235_309#_c_487_n
+ PM_SKY130_FD_SC_HDLL__EINVP_4%A_235_309#
x_PM_SKY130_FD_SC_HDLL__EINVP_4%Z N_Z_M1001_s N_Z_M1008_s N_Z_M1005_s
+ N_Z_M1014_s N_Z_c_501_n N_Z_c_503_n N_Z_c_504_n Z Z Z Z Z N_Z_c_531_n
+ PM_SKY130_FD_SC_HDLL__EINVP_4%Z
x_PM_SKY130_FD_SC_HDLL__EINVP_4%VGND N_VGND_M1013_d N_VGND_M1006_s
+ N_VGND_M1010_s N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n VGND
+ N_VGND_c_560_n N_VGND_c_561_n N_VGND_c_562_n N_VGND_c_563_n N_VGND_c_564_n
+ N_VGND_c_565_n N_VGND_c_566_n N_VGND_c_567_n
+ PM_SKY130_FD_SC_HDLL__EINVP_4%VGND
x_PM_SKY130_FD_SC_HDLL__EINVP_4%A_213_47# N_A_213_47#_M1000_d
+ N_A_213_47#_M1007_d N_A_213_47#_M1001_d N_A_213_47#_M1002_d
+ N_A_213_47#_M1009_d N_A_213_47#_c_638_n N_A_213_47#_c_640_n
+ N_A_213_47#_c_643_n N_A_213_47#_c_645_n N_A_213_47#_c_634_n
+ N_A_213_47#_c_635_n N_A_213_47#_c_636_n N_A_213_47#_c_637_n
+ N_A_213_47#_c_648_n PM_SKY130_FD_SC_HDLL__EINVP_4%A_213_47#
cc_1 VNB N_TE_c_84_n 0.0423276f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_TE_c_85_n 0.0187467f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.96
cc_3 VNB N_TE_c_86_n 0.0180867f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=1.035
cc_4 VNB N_TE_c_87_n 0.0152112f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.96
cc_5 VNB N_TE_c_88_n 0.0185436f $X=-0.19 $Y=-0.24 $X2=1.405 $Y2=1.035
cc_6 VNB N_TE_c_89_n 0.0147241f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.96
cc_7 VNB N_TE_c_90_n 0.0113615f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=1.035
cc_8 VNB N_TE_c_91_n 0.0150799f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.96
cc_9 VNB N_TE_c_92_n 0.0184719f $X=-0.19 $Y=-0.24 $X2=2.345 $Y2=1.035
cc_10 VNB N_TE_c_93_n 0.0184185f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.96
cc_11 VNB N_TE_c_94_n 0.00661167f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.035
cc_12 VNB N_TE_c_95_n 0.00446222f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=1.035
cc_13 VNB N_TE_c_96_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.035
cc_14 VNB TE 0.0134173f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_15 VNB N_A_27_47#_c_166_n 0.0156742f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_16 VNB N_A_27_47#_c_167_n 0.00759518f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_17 VNB N_A_27_47#_c_168_n 7.52914e-19 $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_18 VNB N_A_27_47#_c_169_n 0.00767716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_170_n 0.0303506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_c_281_n 0.0219887f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_21 VNB N_A_c_282_n 0.0160107f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=1.035
cc_22 VNB N_A_M1008_g 0.0184527f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.56
cc_23 VNB N_A_M1009_g 0.0241067f $X=-0.19 $Y=-0.24 $X2=2.345 $Y2=1.035
cc_24 VNB N_A_c_285_n 0.107082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB A 0.0171378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_354_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Z_c_501_n 0.01243f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.56
cc_28 VNB Z 0.00162933f $X=-0.19 $Y=-0.24 $X2=2.345 $Y2=1.035
cc_29 VNB N_VGND_c_557_n 0.00217014f $X=-0.19 $Y=-0.24 $X2=1.405 $Y2=1.035
cc_30 VNB N_VGND_c_558_n 0.00206247f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.56
cc_31 VNB N_VGND_c_559_n 0.00529888f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_32 VNB N_VGND_c_560_n 0.014319f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.96
cc_33 VNB N_VGND_c_561_n 0.0150315f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.035
cc_34 VNB N_VGND_c_562_n 0.0134472f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.035
cc_35 VNB N_VGND_c_563_n 0.0644327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_564_n 0.281286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_565_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_566_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_567_n 0.00592999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_213_47#_c_634_n 0.00681676f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.56
cc_41 VNB N_A_213_47#_c_635_n 0.00333696f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_42 VNB N_A_213_47#_c_636_n 0.00343604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_213_47#_c_637_n 0.0120805f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_44 VPB N_TE_c_84_n 0.0385781f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_45 VPB TE 0.0127325f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_46 VPB N_A_27_47#_c_171_n 0.0195251f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.035
cc_47 VPB N_A_27_47#_c_172_n 0.00987291f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_48 VPB N_A_27_47#_c_173_n 0.0100079f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_49 VPB N_A_27_47#_c_174_n 0.0160921f $X=-0.19 $Y=1.305 $X2=1.405 $Y2=1.035
cc_50 VPB N_A_27_47#_c_175_n 0.00987215f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.56
cc_51 VPB N_A_27_47#_c_176_n 0.0160921f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.035
cc_52 VPB N_A_27_47#_c_177_n 0.00851129f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_53 VPB N_A_27_47#_c_178_n 0.0165132f $X=-0.19 $Y=1.305 $X2=2.345 $Y2=1.035
cc_54 VPB N_A_27_47#_c_179_n 0.0046927f $X=-0.19 $Y=1.305 $X2=2.42 $Y2=0.56
cc_55 VPB N_A_27_47#_c_180_n 0.00597984f $X=-0.19 $Y=1.305 $X2=2.42 $Y2=0.56
cc_56 VPB N_A_27_47#_c_181_n 0.00949374f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.035
cc_57 VPB N_A_27_47#_c_182_n 0.0198657f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_58 VPB N_A_27_47#_c_183_n 0.0173558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_169_n 0.0158945f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_170_n 0.00108677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_c_287_n 0.0164945f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.96
cc_62 VPB N_A_c_288_n 0.015727f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_63 VPB N_A_c_289_n 0.0158638f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.035
cc_64 VPB N_A_c_290_n 0.0198539f $X=-0.19 $Y=1.305 $X2=2.42 $Y2=0.96
cc_65 VPB N_A_c_285_n 0.0441615f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_355_n 0.00773567f $X=-0.19 $Y=1.305 $X2=1.405 $Y2=1.035
cc_67 VPB N_VPWR_c_356_n 0.0185717f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.96
cc_68 VPB N_VPWR_c_357_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=1.555 $Y2=1.035
cc_69 VPB N_VPWR_c_358_n 4.12646e-19 $X=-0.19 $Y=1.305 $X2=2.345 $Y2=1.035
cc_70 VPB N_VPWR_c_359_n 0.0156737f $X=-0.19 $Y=1.305 $X2=2.42 $Y2=0.56
cc_71 VPB N_VPWR_c_360_n 0.00476819f $X=-0.19 $Y=1.305 $X2=2.42 $Y2=0.56
cc_72 VPB N_VPWR_c_361_n 0.0150576f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=1.035
cc_73 VPB N_VPWR_c_362_n 0.0622668f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_354_n 0.0562244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_364_n 0.00638089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_365_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_235_309#_c_429_n 0.00147984f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_78 VPB N_A_235_309#_c_430_n 0.00923042f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.16
cc_79 VPB N_A_235_309#_c_431_n 0.0407578f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_Z_c_503_n 0.00214625f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.96
cc_81 VPB N_Z_c_504_n 0.00176159f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_82 TE N_A_27_47#_M1004_s 0.00430377f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_83 N_TE_c_90_n N_A_27_47#_c_172_n 0.0172013f $X=1.875 $Y=1.035 $X2=0 $Y2=0
cc_84 N_TE_c_95_n N_A_27_47#_c_173_n 0.0172013f $X=1.48 $Y=1.035 $X2=0 $Y2=0
cc_85 N_TE_c_92_n N_A_27_47#_c_175_n 0.0172013f $X=2.345 $Y=1.035 $X2=0 $Y2=0
cc_86 N_TE_c_96_n N_A_27_47#_c_179_n 0.0172013f $X=1.95 $Y=1.035 $X2=0 $Y2=0
cc_87 N_TE_c_85_n N_A_27_47#_c_166_n 0.00442265f $X=0.52 $Y=0.96 $X2=0 $Y2=0
cc_88 N_TE_c_84_n N_A_27_47#_c_182_n 0.00707894f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_89 N_TE_c_84_n N_A_27_47#_c_167_n 0.00511687f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_TE_c_85_n N_A_27_47#_c_167_n 0.0127793f $X=0.52 $Y=0.96 $X2=0 $Y2=0
cc_91 N_TE_c_86_n N_A_27_47#_c_167_n 3.34655e-19 $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_92 N_TE_c_87_n N_A_27_47#_c_167_n 0.00168622f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_93 TE N_A_27_47#_c_167_n 0.0191066f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_94 N_TE_c_84_n N_A_27_47#_c_168_n 0.00162134f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_95 N_TE_c_85_n N_A_27_47#_c_168_n 0.00779754f $X=0.52 $Y=0.96 $X2=0 $Y2=0
cc_96 N_TE_c_86_n N_A_27_47#_c_168_n 0.00304781f $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_97 N_TE_c_87_n N_A_27_47#_c_168_n 0.00305026f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_98 N_TE_c_84_n N_A_27_47#_c_183_n 0.0427271f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_99 N_TE_c_86_n N_A_27_47#_c_183_n 5.728e-19 $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_100 TE N_A_27_47#_c_183_n 0.042355f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_101 N_TE_c_88_n N_A_27_47#_c_169_n 0.0157059f $X=1.405 $Y=1.035 $X2=0 $Y2=0
cc_102 N_TE_c_90_n N_A_27_47#_c_169_n 0.00963839f $X=1.875 $Y=1.035 $X2=0 $Y2=0
cc_103 N_TE_c_92_n N_A_27_47#_c_169_n 0.0158766f $X=2.345 $Y=1.035 $X2=0 $Y2=0
cc_104 N_TE_c_94_n N_A_27_47#_c_169_n 0.0107224f $X=0.99 $Y=1.035 $X2=0 $Y2=0
cc_105 N_TE_c_95_n N_A_27_47#_c_169_n 0.00538458f $X=1.48 $Y=1.035 $X2=0 $Y2=0
cc_106 N_TE_c_96_n N_A_27_47#_c_169_n 0.0051004f $X=1.95 $Y=1.035 $X2=0 $Y2=0
cc_107 N_TE_c_92_n N_A_27_47#_c_170_n 0.00670692f $X=2.345 $Y=1.035 $X2=0 $Y2=0
cc_108 N_TE_c_84_n N_A_27_47#_c_212_n 0.0130842f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_109 N_TE_c_86_n N_A_27_47#_c_212_n 0.0149982f $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_110 N_TE_c_94_n N_A_27_47#_c_212_n 8.40576e-19 $X=0.99 $Y=1.035 $X2=0 $Y2=0
cc_111 TE N_A_27_47#_c_212_n 0.025787f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_112 N_TE_c_84_n N_VPWR_c_355_n 0.0144429f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_113 N_TE_c_84_n N_VPWR_c_361_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_114 N_TE_c_84_n N_VPWR_c_354_n 0.0049402f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_115 N_TE_c_84_n N_A_235_309#_c_432_n 0.00532598f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_116 N_TE_c_90_n N_A_235_309#_c_433_n 2.0345e-19 $X=1.875 $Y=1.035 $X2=0 $Y2=0
cc_117 N_TE_c_84_n N_A_235_309#_c_429_n 6.86088e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_118 N_TE_c_88_n N_A_235_309#_c_429_n 0.00104058f $X=1.405 $Y=1.035 $X2=0
+ $Y2=0
cc_119 N_TE_c_85_n N_VGND_c_557_n 0.0115037f $X=0.52 $Y=0.96 $X2=0 $Y2=0
cc_120 N_TE_c_86_n N_VGND_c_557_n 0.00135012f $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_121 N_TE_c_87_n N_VGND_c_557_n 0.00165782f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_122 N_TE_c_87_n N_VGND_c_558_n 6.09064e-19 $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_123 N_TE_c_89_n N_VGND_c_558_n 0.00993809f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_124 N_TE_c_91_n N_VGND_c_558_n 0.00162962f $X=1.95 $Y=0.96 $X2=0 $Y2=0
cc_125 N_TE_c_91_n N_VGND_c_559_n 6.17073e-19 $X=1.95 $Y=0.96 $X2=0 $Y2=0
cc_126 N_TE_c_93_n N_VGND_c_559_n 0.0110376f $X=2.42 $Y=0.96 $X2=0 $Y2=0
cc_127 N_TE_c_85_n N_VGND_c_560_n 0.00199015f $X=0.52 $Y=0.96 $X2=0 $Y2=0
cc_128 N_TE_c_87_n N_VGND_c_561_n 0.00585385f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_129 N_TE_c_89_n N_VGND_c_561_n 0.00199015f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_130 N_TE_c_91_n N_VGND_c_562_n 0.00428022f $X=1.95 $Y=0.96 $X2=0 $Y2=0
cc_131 N_TE_c_93_n N_VGND_c_562_n 0.00199015f $X=2.42 $Y=0.96 $X2=0 $Y2=0
cc_132 N_TE_c_85_n N_VGND_c_564_n 0.00369362f $X=0.52 $Y=0.96 $X2=0 $Y2=0
cc_133 N_TE_c_87_n N_VGND_c_564_n 0.0108458f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_134 N_TE_c_89_n N_VGND_c_564_n 0.00283749f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_135 N_TE_c_91_n N_VGND_c_564_n 0.005943f $X=1.95 $Y=0.96 $X2=0 $Y2=0
cc_136 N_TE_c_93_n N_VGND_c_564_n 0.00278819f $X=2.42 $Y=0.96 $X2=0 $Y2=0
cc_137 N_TE_c_87_n N_A_213_47#_c_638_n 0.00452417f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_138 N_TE_c_89_n N_A_213_47#_c_638_n 0.00413033f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_139 N_TE_c_89_n N_A_213_47#_c_640_n 0.0103232f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_140 N_TE_c_90_n N_A_213_47#_c_640_n 0.00278658f $X=1.875 $Y=1.035 $X2=0 $Y2=0
cc_141 N_TE_c_91_n N_A_213_47#_c_640_n 0.0113106f $X=1.95 $Y=0.96 $X2=0 $Y2=0
cc_142 N_TE_c_87_n N_A_213_47#_c_643_n 0.00182133f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_143 N_TE_c_88_n N_A_213_47#_c_643_n 0.00310054f $X=1.405 $Y=1.035 $X2=0 $Y2=0
cc_144 N_TE_c_93_n N_A_213_47#_c_645_n 0.00411053f $X=2.42 $Y=0.96 $X2=0 $Y2=0
cc_145 N_TE_c_93_n N_A_213_47#_c_634_n 0.0123079f $X=2.42 $Y=0.96 $X2=0 $Y2=0
cc_146 N_TE_c_93_n N_A_213_47#_c_635_n 0.00365585f $X=2.42 $Y=0.96 $X2=0 $Y2=0
cc_147 N_TE_c_92_n N_A_213_47#_c_648_n 0.00268716f $X=2.345 $Y=1.035 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_178_n N_A_c_287_n 0.0146382f $X=2.945 $Y=1.47 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_181_n N_A_c_287_n 0.00254398f $X=2.885 $Y=1.395 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_169_n N_A_c_285_n 0.00354582f $X=2.86 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_170_n N_A_c_285_n 0.0158325f $X=2.86 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_183_n N_VPWR_M1004_d 0.00571933f $X=0.712 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_153 N_A_27_47#_c_171_n N_VPWR_c_355_n 0.00320248f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_c_182_n N_VPWR_c_355_n 0.0263462f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_183_n N_VPWR_c_355_n 0.0276039f $X=0.712 $Y=1.785 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_171_n N_VPWR_c_356_n 0.00622633f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_171_n N_VPWR_c_357_n 0.0128003f $X=1.535 $Y=1.47 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_174_n N_VPWR_c_357_n 0.0111045f $X=2.005 $Y=1.47 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_176_n N_VPWR_c_357_n 6.18043e-19 $X=2.475 $Y=1.47 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_174_n N_VPWR_c_358_n 6.19581e-19 $X=2.005 $Y=1.47 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_176_n N_VPWR_c_358_n 0.0111045f $X=2.475 $Y=1.47 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_178_n N_VPWR_c_358_n 0.0146227f $X=2.945 $Y=1.47 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_174_n N_VPWR_c_359_n 0.00622633f $X=2.005 $Y=1.47 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_176_n N_VPWR_c_359_n 0.00622633f $X=2.475 $Y=1.47 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_182_n N_VPWR_c_361_n 0.0178308f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_178_n N_VPWR_c_362_n 0.00505556f $X=2.945 $Y=1.47 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_M1004_s N_VPWR_c_354_n 0.00252291f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_171_n N_VPWR_c_354_n 0.0118107f $X=1.535 $Y=1.47 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_174_n N_VPWR_c_354_n 0.0104011f $X=2.005 $Y=1.47 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_176_n N_VPWR_c_354_n 0.0104011f $X=2.475 $Y=1.47 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_178_n N_VPWR_c_354_n 0.00870867f $X=2.945 $Y=1.47 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_182_n N_VPWR_c_354_n 0.00986266f $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_183_n N_VPWR_c_354_n 0.00695765f $X=0.712 $Y=1.785 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_171_n N_A_235_309#_c_432_n 0.0124981f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_183_n N_A_235_309#_c_432_n 0.014384f $X=0.712 $Y=1.785 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_171_n N_A_235_309#_c_433_n 0.018301f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_172_n N_A_235_309#_c_433_n 0.0024163f $X=1.915 $Y=1.395
+ $X2=0 $Y2=0
cc_178 N_A_27_47#_c_174_n N_A_235_309#_c_433_n 0.0170681f $X=2.005 $Y=1.47 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_169_n N_A_235_309#_c_433_n 0.0375096f $X=2.86 $Y=1.16 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_183_n N_A_235_309#_c_429_n 0.0113703f $X=0.712 $Y=1.785
+ $X2=0 $Y2=0
cc_181 N_A_27_47#_c_169_n N_A_235_309#_c_429_n 0.0146313f $X=2.86 $Y=1.16 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_174_n N_A_235_309#_c_444_n 0.00546277f $X=2.005 $Y=1.47
+ $X2=0 $Y2=0
cc_183 N_A_27_47#_c_176_n N_A_235_309#_c_444_n 0.00546277f $X=2.475 $Y=1.47
+ $X2=0 $Y2=0
cc_184 N_A_27_47#_c_176_n N_A_235_309#_c_446_n 0.0171405f $X=2.475 $Y=1.47 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_177_n N_A_235_309#_c_446_n 0.00262074f $X=2.725 $Y=1.395
+ $X2=0 $Y2=0
cc_186 N_A_27_47#_c_178_n N_A_235_309#_c_446_n 0.0161333f $X=2.945 $Y=1.47 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_169_n N_A_235_309#_c_446_n 0.051295f $X=2.86 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_178_n N_A_235_309#_c_450_n 0.00469508f $X=2.945 $Y=1.47
+ $X2=0 $Y2=0
cc_189 N_A_27_47#_c_175_n N_A_235_309#_c_451_n 0.0025662f $X=2.385 $Y=1.395
+ $X2=0 $Y2=0
cc_190 N_A_27_47#_c_169_n N_A_235_309#_c_451_n 0.0111227f $X=2.86 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_181_n Z 6.98272e-19 $X=2.885 $Y=1.395 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_169_n Z 0.0286243f $X=2.86 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_170_n Z 2.3221e-19 $X=2.86 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_178_n Z 4.6355e-19 $X=2.945 $Y=1.47 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_167_n N_VGND_M1013_d 0.00326346f $X=0.622 $Y=0.825 $X2=-0.19
+ $Y2=-0.24
cc_196 N_A_27_47#_c_168_n N_VGND_M1013_d 9.97407e-19 $X=0.622 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_197 N_A_27_47#_c_166_n N_VGND_c_557_n 0.0177195f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_167_n N_VGND_c_557_n 0.012775f $X=0.622 $Y=0.825 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_212_n N_VGND_c_557_n 0.00474116f $X=0.712 $Y=1.16 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_166_n N_VGND_c_560_n 0.0175229f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_167_n N_VGND_c_560_n 0.00236869f $X=0.622 $Y=0.825 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_M1013_s N_VGND_c_564_n 0.00293425f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_166_n N_VGND_c_564_n 0.00980382f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_167_n N_VGND_c_564_n 0.0054368f $X=0.622 $Y=0.825 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_173_n N_A_213_47#_c_640_n 2.24658e-19 $X=1.625 $Y=1.395
+ $X2=0 $Y2=0
cc_206 N_A_27_47#_c_169_n N_A_213_47#_c_640_n 0.0479154f $X=2.86 $Y=1.16 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_167_n N_A_213_47#_c_643_n 0.00815106f $X=0.622 $Y=0.825
+ $X2=0 $Y2=0
cc_208 N_A_27_47#_c_169_n N_A_213_47#_c_643_n 0.0138439f $X=2.86 $Y=1.16 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_180_n N_A_213_47#_c_634_n 7.28392e-19 $X=2.475 $Y=1.395
+ $X2=0 $Y2=0
cc_210 N_A_27_47#_c_169_n N_A_213_47#_c_634_n 0.0795607f $X=2.86 $Y=1.16 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_170_n N_A_213_47#_c_634_n 0.00836703f $X=2.86 $Y=1.16 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_169_n N_A_213_47#_c_648_n 0.0135367f $X=2.86 $Y=1.16 $X2=0
+ $Y2=0
cc_213 N_A_c_287_n N_VPWR_c_358_n 9.84138e-19 $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_c_287_n N_VPWR_c_362_n 0.00429453f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_c_288_n N_VPWR_c_362_n 0.00429453f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_c_289_n N_VPWR_c_362_n 0.00429453f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_c_290_n N_VPWR_c_362_n 0.00429453f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_c_287_n N_VPWR_c_354_n 0.00621534f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A_c_288_n N_VPWR_c_354_n 0.00606499f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A_c_289_n N_VPWR_c_354_n 0.00606499f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A_c_290_n N_VPWR_c_354_n 0.00708599f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_c_287_n N_A_235_309#_c_446_n 0.00156101f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_c_287_n N_A_235_309#_c_450_n 0.0046027f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_c_287_n N_A_235_309#_c_455_n 0.0122062f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_c_288_n N_A_235_309#_c_455_n 0.013747f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A_c_289_n N_A_235_309#_c_430_n 0.0122476f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A_c_290_n N_A_235_309#_c_430_n 0.0137768f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_c_290_n N_A_235_309#_c_431_n 0.013169f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_c_285_n N_A_235_309#_c_431_n 0.00515666f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_230 A N_A_235_309#_c_431_n 0.0319592f $X=5.285 $Y=1.19 $X2=0 $Y2=0
cc_231 N_A_M1008_g N_Z_c_501_n 0.00992634f $X=4.385 $Y=0.56 $X2=0 $Y2=0
cc_232 N_A_M1009_g N_Z_c_501_n 0.0118443f $X=4.855 $Y=0.56 $X2=0 $Y2=0
cc_233 N_A_c_285_n N_Z_c_501_n 0.0115774f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_234 A N_Z_c_501_n 0.0815457f $X=5.285 $Y=1.19 $X2=0 $Y2=0
cc_235 N_A_c_289_n N_Z_c_503_n 0.0101048f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_c_285_n N_Z_c_503_n 0.0080139f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_237 A N_Z_c_503_n 0.0157686f $X=5.285 $Y=1.19 $X2=0 $Y2=0
cc_238 N_A_c_288_n N_Z_c_504_n 5.88772e-19 $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_c_289_n N_Z_c_504_n 0.0119866f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A_c_290_n N_Z_c_504_n 0.00940337f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A_c_285_n N_Z_c_504_n 0.00746666f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_242 A N_Z_c_504_n 0.031085f $X=5.285 $Y=1.19 $X2=0 $Y2=0
cc_243 N_A_c_281_n Z 0.011715f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_c_287_n Z 0.00120118f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A_c_282_n Z 0.012205f $X=3.915 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_c_288_n Z 0.00144916f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_M1008_g Z 0.00323572f $X=4.385 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A_c_289_n Z 2.10507e-19 $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_249 N_A_c_285_n Z 0.0408261f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_250 A Z 0.020034f $X=5.285 $Y=1.19 $X2=0 $Y2=0
cc_251 N_A_c_287_n Z 0.004285f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A_c_288_n Z 0.0137556f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_c_287_n N_Z_c_531_n 0.00862602f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A_c_288_n N_Z_c_531_n 0.00742548f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_c_289_n N_Z_c_531_n 5.51873e-19 $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_c_285_n N_Z_c_531_n 9.31598e-19 $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_257 N_A_c_281_n N_VGND_c_559_n 0.00276998f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A_c_281_n N_VGND_c_563_n 0.00357877f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_c_282_n N_VGND_c_563_n 0.00357877f $X=3.915 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_M1008_g N_VGND_c_563_n 0.00357877f $X=4.385 $Y=0.56 $X2=0 $Y2=0
cc_261 N_A_M1009_g N_VGND_c_563_n 0.00357877f $X=4.855 $Y=0.56 $X2=0 $Y2=0
cc_262 N_A_c_281_n N_VGND_c_564_n 0.00677297f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A_c_282_n N_VGND_c_564_n 0.00548399f $X=3.915 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A_M1008_g N_VGND_c_564_n 0.00548399f $X=4.385 $Y=0.56 $X2=0 $Y2=0
cc_265 N_A_M1009_g N_VGND_c_564_n 0.0064529f $X=4.855 $Y=0.56 $X2=0 $Y2=0
cc_266 N_A_c_281_n N_A_213_47#_c_637_n 0.0145888f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_c_282_n N_A_213_47#_c_637_n 0.00902754f $X=3.915 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_M1008_g N_A_213_47#_c_637_n 0.00903374f $X=4.385 $Y=0.56 $X2=0 $Y2=0
cc_269 N_A_M1009_g N_A_213_47#_c_637_n 0.00903374f $X=4.855 $Y=0.56 $X2=0 $Y2=0
cc_270 N_A_c_285_n N_A_213_47#_c_637_n 4.68623e-19 $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_271 N_VPWR_c_354_n N_A_235_309#_M1003_s 0.00429283f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_272 N_VPWR_c_354_n N_A_235_309#_M1011_s 0.00647849f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_354_n N_A_235_309#_M1016_s 0.00584403f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_354_n N_A_235_309#_M1012_d 0.00231272f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_354_n N_A_235_309#_M1017_d 0.00217523f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_355_n N_A_235_309#_c_432_n 0.0207729f $X=0.73 $Y=2.34 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_356_n N_A_235_309#_c_432_n 0.0146267f $X=1.605 $Y=2.72 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_357_n N_A_235_309#_c_432_n 0.0350594f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_354_n N_A_235_309#_c_432_n 0.00801045f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_280 N_VPWR_M1003_d N_A_235_309#_c_433_n 0.00357692f $X=1.625 $Y=1.545 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_357_n N_A_235_309#_c_433_n 0.0171295f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_357_n N_A_235_309#_c_444_n 0.0345089f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_358_n N_A_235_309#_c_444_n 0.0347423f $X=2.71 $Y=2.02 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_359_n N_A_235_309#_c_444_n 0.0118139f $X=2.545 $Y=2.72 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_354_n N_A_235_309#_c_444_n 0.00646998f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_286 N_VPWR_M1015_d N_A_235_309#_c_446_n 0.0036863f $X=2.565 $Y=1.545 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_358_n N_A_235_309#_c_446_n 0.0194148f $X=2.71 $Y=2.02 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_358_n N_A_235_309#_c_450_n 0.0243508f $X=2.71 $Y=2.02 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_362_n N_A_235_309#_c_455_n 0.0431443f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_354_n N_A_235_309#_c_455_n 0.0278172f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_358_n N_A_235_309#_c_482_n 0.0115776f $X=2.71 $Y=2.02 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_362_n N_A_235_309#_c_482_n 0.0119545f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_354_n N_A_235_309#_c_482_n 0.006547f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_c_362_n N_A_235_309#_c_430_n 0.0684239f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_354_n N_A_235_309#_c_430_n 0.0415073f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_362_n N_A_235_309#_c_487_n 0.0119545f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_354_n N_A_235_309#_c_487_n 0.006547f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_298 N_VPWR_c_354_n N_Z_M1005_s 0.00232895f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_299 N_VPWR_c_354_n N_Z_M1014_s 0.00232895f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_300 N_A_235_309#_c_455_n N_Z_M1005_s 0.00352848f $X=4.09 $Y=2.38 $X2=0 $Y2=0
cc_301 N_A_235_309#_c_430_n N_Z_M1014_s 0.00352392f $X=5.03 $Y=2.38 $X2=0 $Y2=0
cc_302 N_A_235_309#_M1012_d N_Z_c_503_n 0.00178587f $X=4.03 $Y=1.485 $X2=0 $Y2=0
cc_303 N_A_235_309#_c_492_p N_Z_c_503_n 0.0136682f $X=4.175 $Y=1.96 $X2=0 $Y2=0
cc_304 N_A_235_309#_c_492_p N_Z_c_504_n 0.0253827f $X=4.175 $Y=1.96 $X2=0 $Y2=0
cc_305 N_A_235_309#_c_430_n N_Z_c_504_n 0.0196128f $X=5.03 $Y=2.38 $X2=0 $Y2=0
cc_306 N_A_235_309#_c_431_n N_Z_c_504_n 0.0447996f $X=5.22 $Y=2.295 $X2=0 $Y2=0
cc_307 N_A_235_309#_c_446_n Z 0.00471239f $X=3.125 $Y=1.64 $X2=0 $Y2=0
cc_308 N_A_235_309#_c_446_n N_Z_c_531_n 0.00821099f $X=3.125 $Y=1.64 $X2=0 $Y2=0
cc_309 N_A_235_309#_c_450_n N_Z_c_531_n 0.0268778f $X=3.21 $Y=1.96 $X2=0 $Y2=0
cc_310 N_A_235_309#_c_455_n N_Z_c_531_n 0.0191829f $X=4.09 $Y=2.38 $X2=0 $Y2=0
cc_311 N_A_235_309#_c_492_p N_Z_c_531_n 0.0208308f $X=4.175 $Y=1.96 $X2=0 $Y2=0
cc_312 N_Z_M1001_s N_VGND_c_564_n 0.00256987f $X=3.52 $Y=0.235 $X2=0 $Y2=0
cc_313 N_Z_M1008_s N_VGND_c_564_n 0.00256987f $X=4.46 $Y=0.235 $X2=0 $Y2=0
cc_314 N_Z_c_501_n N_A_213_47#_M1002_d 0.00490548f $X=4.645 $Y=0.76 $X2=0 $Y2=0
cc_315 N_Z_c_501_n N_A_213_47#_M1009_d 0.00684154f $X=4.645 $Y=0.76 $X2=0 $Y2=0
cc_316 N_Z_M1001_s N_A_213_47#_c_637_n 0.00399738f $X=3.52 $Y=0.235 $X2=0 $Y2=0
cc_317 N_Z_M1008_s N_A_213_47#_c_637_n 0.00401386f $X=4.46 $Y=0.235 $X2=0 $Y2=0
cc_318 N_Z_c_501_n N_A_213_47#_c_637_n 0.0797406f $X=4.645 $Y=0.76 $X2=0 $Y2=0
cc_319 Z N_A_213_47#_c_637_n 0.0291055f $X=3.74 $Y=0.765 $X2=0 $Y2=0
cc_320 N_VGND_c_564_n N_A_213_47#_M1000_d 0.00560278f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_321 N_VGND_c_564_n N_A_213_47#_M1007_d 0.00316288f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_564_n N_A_213_47#_M1001_d 0.00210127f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_564_n N_A_213_47#_M1002_d 0.00255381f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_324 N_VGND_c_564_n N_A_213_47#_M1009_d 0.00266737f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_325 N_VGND_c_558_n N_A_213_47#_c_638_n 0.0171708f $X=1.69 $Y=0.36 $X2=0 $Y2=0
cc_326 N_VGND_c_561_n N_A_213_47#_c_638_n 0.0116627f $X=1.475 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_564_n N_A_213_47#_c_638_n 0.00644035f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_M1006_s N_A_213_47#_c_640_n 0.0038973f $X=1.555 $Y=0.235 $X2=0
+ $Y2=0
cc_329 N_VGND_c_558_n N_A_213_47#_c_640_n 0.0214497f $X=1.69 $Y=0.36 $X2=0 $Y2=0
cc_330 N_VGND_c_561_n N_A_213_47#_c_640_n 0.0023206f $X=1.475 $Y=0 $X2=0 $Y2=0
cc_331 N_VGND_c_562_n N_A_213_47#_c_640_n 0.0029785f $X=2.415 $Y=0 $X2=0 $Y2=0
cc_332 N_VGND_c_564_n N_A_213_47#_c_640_n 0.0113285f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_333 N_VGND_c_559_n N_A_213_47#_c_645_n 0.0172059f $X=2.63 $Y=0.36 $X2=0 $Y2=0
cc_334 N_VGND_c_562_n N_A_213_47#_c_645_n 0.011459f $X=2.415 $Y=0 $X2=0 $Y2=0
cc_335 N_VGND_c_564_n N_A_213_47#_c_645_n 0.00644035f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_336 N_VGND_M1010_s N_A_213_47#_c_634_n 0.00522868f $X=2.495 $Y=0.235 $X2=0
+ $Y2=0
cc_337 N_VGND_c_559_n N_A_213_47#_c_634_n 0.0250655f $X=2.63 $Y=0.36 $X2=0 $Y2=0
cc_338 N_VGND_c_562_n N_A_213_47#_c_634_n 0.0023206f $X=2.415 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_c_563_n N_A_213_47#_c_634_n 0.0031369f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_340 N_VGND_c_564_n N_A_213_47#_c_634_n 0.0110996f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_341 N_VGND_c_559_n N_A_213_47#_c_635_n 0.00158182f $X=2.63 $Y=0.36 $X2=0
+ $Y2=0
cc_342 N_VGND_c_559_n N_A_213_47#_c_636_n 0.0180544f $X=2.63 $Y=0.36 $X2=0 $Y2=0
cc_343 N_VGND_c_563_n N_A_213_47#_c_636_n 0.0231841f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_344 N_VGND_c_564_n N_A_213_47#_c_636_n 0.0128424f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_345 N_VGND_c_563_n N_A_213_47#_c_637_n 0.12028f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_564_n N_A_213_47#_c_637_n 0.0752499f $X=5.29 $Y=0 $X2=0 $Y2=0
