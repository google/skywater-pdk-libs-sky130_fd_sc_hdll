# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2i_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.720000 1.075000 4.025000 1.275000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.710000 0.995000 5.085000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.832500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.830000 1.325000 ;
        RECT 0.630000 0.725000 0.830000 0.995000 ;
    END
  END S
  PIN VGND
    ANTENNADIFFAREA  0.585000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.850000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.796250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 0.295000 5.425000 0.465000 ;
        RECT 2.965000 2.255000 5.425000 2.425000 ;
        RECT 5.200000 1.785000 5.425000 2.255000 ;
        RECT 5.255000 0.465000 5.425000 1.785000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.675000 ;
      RECT 0.085000  0.675000 0.260000 1.495000 ;
      RECT 0.085000  1.495000 1.545000 1.665000 ;
      RECT 0.085000  1.665000 0.260000 2.135000 ;
      RECT 0.085000  2.135000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.885000 0.545000 ;
      RECT 0.515000  2.255000 0.895000 2.635000 ;
      RECT 0.985000  1.835000 1.885000 2.005000 ;
      RECT 1.115000  0.575000 1.355000 0.935000 ;
      RECT 1.325000  1.155000 2.185000 1.325000 ;
      RECT 1.325000  1.325000 1.545000 1.495000 ;
      RECT 1.455000  2.255000 1.835000 2.635000 ;
      RECT 1.585000  0.085000 1.835000 0.885000 ;
      RECT 1.715000  1.495000 3.765000 1.665000 ;
      RECT 1.715000  1.665000 1.885000 1.835000 ;
      RECT 1.805000  1.075000 2.185000 1.155000 ;
      RECT 2.055000  0.295000 2.225000 0.735000 ;
      RECT 2.055000  0.735000 3.765000 0.905000 ;
      RECT 2.055000  2.135000 2.280000 2.465000 ;
      RECT 2.110000  1.835000 3.135000 1.915000 ;
      RECT 2.110000  1.915000 4.750000 2.005000 ;
      RECT 2.110000  2.005000 2.280000 2.135000 ;
      RECT 2.525000  0.085000 2.695000 0.545000 ;
      RECT 2.525000  2.175000 2.775000 2.635000 ;
      RECT 2.965000  2.005000 4.750000 2.085000 ;
      RECT 3.385000  0.655000 3.765000 0.735000 ;
      RECT 3.385000  1.665000 3.765000 1.715000 ;
      RECT 4.200000  0.655000 4.745000 0.825000 ;
      RECT 4.200000  0.825000 4.505000 0.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.170000  0.765000 1.340000 0.935000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.200000  0.765000 4.370000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 1.110000 0.735000 1.400000 0.780000 ;
      RECT 1.110000 0.780000 4.480000 0.920000 ;
      RECT 1.110000 0.920000 1.400000 0.965000 ;
      RECT 4.140000 0.735000 4.480000 0.780000 ;
      RECT 4.140000 0.920000 4.480000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2i_2
END LIBRARY
