* File: sky130_fd_sc_hdll__a22oi_4.pxi.spice
* Created: Thu Aug 27 18:54:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__A22OI_4%B2 N_B2_c_107_n N_B2_M1008_g N_B2_c_113_n
+ N_B2_M1002_g N_B2_c_108_n N_B2_M1010_g N_B2_c_114_n N_B2_M1013_g N_B2_c_109_n
+ N_B2_M1024_g N_B2_c_115_n N_B2_M1021_g N_B2_c_116_n N_B2_M1028_g N_B2_c_110_n
+ N_B2_M1030_g B2 N_B2_c_111_n N_B2_c_112_n B2 PM_SKY130_FD_SC_HDLL__A22OI_4%B2
x_PM_SKY130_FD_SC_HDLL__A22OI_4%B1 N_B1_c_190_n N_B1_M1015_g N_B1_c_196_n
+ N_B1_M1000_g N_B1_c_191_n N_B1_M1018_g N_B1_c_197_n N_B1_M1006_g N_B1_c_192_n
+ N_B1_M1026_g N_B1_c_198_n N_B1_M1009_g N_B1_c_193_n N_B1_M1027_g N_B1_c_199_n
+ N_B1_M1016_g B1 N_B1_c_194_n N_B1_c_195_n B1 PM_SKY130_FD_SC_HDLL__A22OI_4%B1
x_PM_SKY130_FD_SC_HDLL__A22OI_4%A1 N_A1_c_260_n N_A1_M1005_g N_A1_c_266_n
+ N_A1_M1004_g N_A1_c_261_n N_A1_M1012_g N_A1_c_267_n N_A1_M1007_g N_A1_c_262_n
+ N_A1_M1023_g N_A1_c_268_n N_A1_M1019_g N_A1_c_269_n N_A1_M1029_g N_A1_c_263_n
+ N_A1_M1031_g A1 N_A1_c_264_n N_A1_c_265_n A1 PM_SKY130_FD_SC_HDLL__A22OI_4%A1
x_PM_SKY130_FD_SC_HDLL__A22OI_4%A2 N_A2_c_322_n N_A2_M1001_g N_A2_c_328_n
+ N_A2_M1011_g N_A2_c_323_n N_A2_M1003_g N_A2_c_329_n N_A2_M1017_g N_A2_c_324_n
+ N_A2_M1014_g N_A2_c_330_n N_A2_M1022_g N_A2_c_331_n N_A2_M1025_g N_A2_c_325_n
+ N_A2_M1020_g A2 N_A2_c_326_n N_A2_c_327_n A2 PM_SKY130_FD_SC_HDLL__A22OI_4%A2
x_PM_SKY130_FD_SC_HDLL__A22OI_4%A_27_297# N_A_27_297#_M1002_d
+ N_A_27_297#_M1013_d N_A_27_297#_M1028_d N_A_27_297#_M1006_d
+ N_A_27_297#_M1016_d N_A_27_297#_M1007_s N_A_27_297#_M1029_s
+ N_A_27_297#_M1017_s N_A_27_297#_M1025_s N_A_27_297#_c_397_n
+ N_A_27_297#_c_398_n N_A_27_297#_c_413_n N_A_27_297#_c_461_p
+ N_A_27_297#_c_415_n N_A_27_297#_c_452_p N_A_27_297#_c_417_n
+ N_A_27_297#_c_457_p N_A_27_297#_c_419_n N_A_27_297#_c_399_n
+ N_A_27_297#_c_482_p N_A_27_297#_c_400_n N_A_27_297#_c_486_p
+ N_A_27_297#_c_401_n N_A_27_297#_c_487_p N_A_27_297#_c_402_n
+ N_A_27_297#_c_488_p N_A_27_297#_c_403_n N_A_27_297#_c_404_n
+ N_A_27_297#_c_489_p N_A_27_297#_c_483_p N_A_27_297#_c_484_p
+ N_A_27_297#_c_485_p N_A_27_297#_c_405_n N_A_27_297#_c_406_n
+ N_A_27_297#_c_407_n PM_SKY130_FD_SC_HDLL__A22OI_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A22OI_4%Y N_Y_M1015_s N_Y_M1026_s N_Y_M1005_s
+ N_Y_M1023_s N_Y_M1002_s N_Y_M1021_s N_Y_M1000_s N_Y_M1009_s N_Y_c_515_n
+ N_Y_c_540_n N_Y_c_513_n N_Y_c_514_n N_Y_c_517_n N_Y_c_518_n N_Y_c_519_n
+ N_Y_c_520_n N_Y_c_521_n Y Y PM_SKY130_FD_SC_HDLL__A22OI_4%Y
x_PM_SKY130_FD_SC_HDLL__A22OI_4%VPWR N_VPWR_M1004_d N_VPWR_M1019_d
+ N_VPWR_M1011_d N_VPWR_M1022_d N_VPWR_c_613_n N_VPWR_c_614_n N_VPWR_c_615_n
+ N_VPWR_c_616_n N_VPWR_c_617_n N_VPWR_c_618_n N_VPWR_c_619_n N_VPWR_c_620_n
+ N_VPWR_c_621_n N_VPWR_c_622_n N_VPWR_c_623_n N_VPWR_c_624_n VPWR
+ N_VPWR_c_625_n N_VPWR_c_612_n PM_SKY130_FD_SC_HDLL__A22OI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A22OI_4%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1010_s
+ N_A_27_47#_M1030_s N_A_27_47#_M1018_d N_A_27_47#_M1027_d N_A_27_47#_c_714_n
+ N_A_27_47#_c_715_n N_A_27_47#_c_716_n N_A_27_47#_c_729_n N_A_27_47#_c_717_n
+ N_A_27_47#_c_737_n N_A_27_47#_c_718_n N_A_27_47#_c_719_n N_A_27_47#_c_720_n
+ PM_SKY130_FD_SC_HDLL__A22OI_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__A22OI_4%VGND N_VGND_M1008_d N_VGND_M1024_d
+ N_VGND_M1001_s N_VGND_M1014_s N_VGND_c_786_n N_VGND_c_787_n N_VGND_c_788_n
+ N_VGND_c_789_n N_VGND_c_790_n N_VGND_c_791_n N_VGND_c_792_n N_VGND_c_793_n
+ N_VGND_c_794_n VGND N_VGND_c_795_n N_VGND_c_796_n N_VGND_c_797_n
+ N_VGND_c_798_n VGND PM_SKY130_FD_SC_HDLL__A22OI_4%VGND
x_PM_SKY130_FD_SC_HDLL__A22OI_4%A_883_47# N_A_883_47#_M1005_d
+ N_A_883_47#_M1012_d N_A_883_47#_M1031_d N_A_883_47#_M1003_d
+ N_A_883_47#_M1020_d N_A_883_47#_c_899_n N_A_883_47#_c_911_n
+ N_A_883_47#_c_900_n N_A_883_47#_c_901_n N_A_883_47#_c_919_n
+ N_A_883_47#_c_902_n N_A_883_47#_c_903_n N_A_883_47#_c_904_n
+ PM_SKY130_FD_SC_HDLL__A22OI_4%A_883_47#
cc_1 VNB N_B2_c_107_n 0.0219568f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B2_c_108_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_B2_c_109_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_4 VNB N_B2_c_110_n 0.0169251f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_B2_c_111_n 0.0179004f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.16
cc_6 VNB N_B2_c_112_n 0.0804963f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_7 VNB N_B1_c_190_n 0.0162503f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_B1_c_191_n 0.0168735f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_9 VNB N_B1_c_192_n 0.0169133f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_10 VNB N_B1_c_193_n 0.0223829f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_11 VNB N_B1_c_194_n 0.0886192f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.16
cc_12 VNB N_B1_c_195_n 0.0100559f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_13 VNB N_A1_c_260_n 0.0223829f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_A1_c_261_n 0.0169186f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_15 VNB N_A1_c_262_n 0.0173597f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_16 VNB N_A1_c_263_n 0.0171706f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_17 VNB N_A1_c_264_n 0.00333731f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.16
cc_18 VNB N_A1_c_265_n 0.0765141f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_19 VNB N_A2_c_322_n 0.0164927f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_20 VNB N_A2_c_323_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_21 VNB N_A2_c_324_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_22 VNB N_A2_c_325_n 0.0223965f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_23 VNB N_A2_c_326_n 0.0236945f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.16
cc_24 VNB N_A2_c_327_n 0.0801709f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_25 VNB N_Y_c_513_n 0.00106016f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.202
cc_26 VNB N_Y_c_514_n 0.00813346f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.175
cc_27 VNB N_VPWR_c_612_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_714_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_29 VNB N_A_27_47#_c_715_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_30 VNB N_A_27_47#_c_716_n 0.010462f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_31 VNB N_A_27_47#_c_717_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_718_n 0.00299398f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.202
cc_33 VNB N_A_27_47#_c_719_n 0.00262034f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.202
cc_34 VNB N_A_27_47#_c_720_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.202
cc_35 VNB N_VGND_c_786_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_36 VNB N_VGND_c_787_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_37 VNB N_VGND_c_788_n 0.00469188f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_38 VNB N_VGND_c_789_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.202
cc_39 VNB N_VGND_c_790_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_40 VNB N_VGND_c_791_n 0.115022f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.202
cc_41 VNB N_VGND_c_792_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_42 VNB N_VGND_c_793_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.16
cc_43 VNB N_VGND_c_794_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.16
cc_44 VNB N_VGND_c_795_n 0.0240576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_796_n 0.420295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_797_n 0.0218673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_798_n 0.00323927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_883_47#_c_899_n 0.0026606f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_49 VNB N_A_883_47#_c_900_n 0.00337803f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_50 VNB N_A_883_47#_c_901_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_51 VNB N_A_883_47#_c_902_n 0.0132268f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_52 VNB N_A_883_47#_c_903_n 0.0187437f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.202
cc_53 VNB N_A_883_47#_c_904_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=1.202
cc_54 VPB N_B2_c_113_n 0.0204632f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_55 VPB N_B2_c_114_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_56 VPB N_B2_c_115_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_57 VPB N_B2_c_116_n 0.015983f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_58 VPB N_B2_c_112_n 0.0500567f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_59 VPB N_B1_c_196_n 0.0158458f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_60 VPB N_B1_c_197_n 0.0158618f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_61 VPB N_B1_c_198_n 0.0158721f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_62 VPB N_B1_c_199_n 0.0202815f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_63 VPB N_B1_c_194_n 0.0541413f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.16
cc_64 VPB N_A1_c_266_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_65 VPB N_A1_c_267_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_66 VPB N_A1_c_268_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_67 VPB N_A1_c_269_n 0.0161064f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_68 VPB N_A1_c_265_n 0.0479065f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_69 VPB N_A2_c_328_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_70 VPB N_A2_c_329_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_71 VPB N_A2_c_330_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_72 VPB N_A2_c_331_n 0.0203443f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_73 VPB N_A2_c_327_n 0.048391f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_74 VPB N_A_27_297#_c_397_n 0.00753428f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_75 VPB N_A_27_297#_c_398_n 0.035724f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_76 VPB N_A_27_297#_c_399_n 0.00909917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_297#_c_400_n 0.00201926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_297#_c_401_n 0.00218917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_297#_c_402_n 0.00196267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_297#_c_403_n 0.00196267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_297#_c_404_n 0.00366598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_297#_c_405_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_297#_c_406_n 0.00469599f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_297#_c_407_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_Y_c_515_n 0.00477553f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.202
cc_86 VPB N_Y_c_513_n 0.00115826f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.202
cc_87 VPB N_Y_c_517_n 0.00196802f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.175
cc_88 VPB N_Y_c_518_n 0.00192868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_Y_c_519_n 0.0014926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_Y_c_520_n 3.11328e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_Y_c_521_n 0.00188656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB Y 0.00160976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_613_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.56
cc_94 VPB N_VPWR_c_614_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_95 VPB N_VPWR_c_615_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_96 VPB N_VPWR_c_616_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.202
cc_97 VPB N_VPWR_c_617_n 0.113457f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_98 VPB N_VPWR_c_618_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_99 VPB N_VPWR_c_619_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_100 VPB N_VPWR_c_620_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.202
cc_101 VPB N_VPWR_c_621_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.202
cc_102 VPB N_VPWR_c_622_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.16
cc_103 VPB N_VPWR_c_623_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_104 VPB N_VPWR_c_624_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.202
cc_105 VPB N_VPWR_c_625_n 0.0247905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_612_n 0.0525676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 N_B2_c_110_n N_B1_c_190_n 0.0167521f $X=1.93 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_108 N_B2_c_116_n N_B1_c_196_n 0.0214204f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_109 N_B2_c_111_n N_B1_c_194_n 0.00189067f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B2_c_112_n N_B1_c_194_n 0.0167521f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_111 N_B2_c_113_n N_A_27_297#_c_397_n 4.66918e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B2_c_113_n N_A_27_297#_c_398_n 0.0120287f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B2_c_114_n N_A_27_297#_c_398_n 6.66791e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B2_c_111_n N_A_27_297#_c_398_n 0.0271108f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_115 N_B2_c_112_n N_A_27_297#_c_398_n 3.18853e-19 $X=1.905 $Y=1.202 $X2=0
+ $Y2=0
cc_116 N_B2_c_113_n N_A_27_297#_c_413_n 0.0129846f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_117 N_B2_c_114_n N_A_27_297#_c_413_n 0.01161f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B2_c_115_n N_A_27_297#_c_415_n 0.01161f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B2_c_116_n N_A_27_297#_c_415_n 0.01161f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B2_c_116_n N_Y_c_515_n 0.0132696f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B2_c_111_n N_Y_c_515_n 0.0214433f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_122 N_B2_c_112_n N_Y_c_515_n 8.96166e-19 $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_123 N_B2_c_110_n N_Y_c_513_n 9.31031e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B2_c_111_n N_Y_c_513_n 0.0108693f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_125 N_B2_c_112_n N_Y_c_513_n 9.18042e-19 $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_126 N_B2_c_114_n N_Y_c_518_n 0.013205f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_127 N_B2_c_115_n N_Y_c_518_n 0.0132696f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B2_c_111_n N_Y_c_518_n 0.0487345f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_129 N_B2_c_112_n N_Y_c_518_n 0.00876269f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_130 N_B2_c_111_n N_Y_c_519_n 0.020385f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B2_c_112_n N_Y_c_519_n 0.00642616f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_132 N_B2_c_113_n Y 0.0012736f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_133 N_B2_c_111_n Y 0.0171234f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_134 N_B2_c_112_n Y 0.00552124f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_135 N_B2_c_113_n N_VPWR_c_617_n 0.00429425f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B2_c_114_n N_VPWR_c_617_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B2_c_115_n N_VPWR_c_617_n 0.00429453f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_138 N_B2_c_116_n N_VPWR_c_617_n 0.00429453f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B2_c_113_n N_VPWR_c_612_n 0.0069764f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B2_c_114_n N_VPWR_c_612_n 0.00606499f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B2_c_115_n N_VPWR_c_612_n 0.00606499f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B2_c_116_n N_VPWR_c_612_n 0.00609021f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B2_c_107_n N_A_27_47#_c_714_n 0.00686626f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B2_c_108_n N_A_27_47#_c_714_n 5.46296e-19 $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_145 N_B2_c_107_n N_A_27_47#_c_715_n 0.00901745f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B2_c_108_n N_A_27_47#_c_715_n 0.00901745f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_147 N_B2_c_111_n N_A_27_47#_c_715_n 0.0397461f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_148 N_B2_c_112_n N_A_27_47#_c_715_n 0.00345541f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_149 N_B2_c_107_n N_A_27_47#_c_716_n 0.00129539f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_150 N_B2_c_111_n N_A_27_47#_c_716_n 0.0278303f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_151 N_B2_c_107_n N_A_27_47#_c_729_n 5.24597e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B2_c_108_n N_A_27_47#_c_729_n 0.00651696f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B2_c_109_n N_A_27_47#_c_729_n 0.00693563f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B2_c_110_n N_A_27_47#_c_729_n 5.34196e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B2_c_109_n N_A_27_47#_c_717_n 0.00929182f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_156 N_B2_c_110_n N_A_27_47#_c_717_n 0.00650032f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_157 N_B2_c_111_n N_A_27_47#_c_717_n 0.0399344f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_158 N_B2_c_112_n N_A_27_47#_c_717_n 0.00468948f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_159 N_B2_c_110_n N_A_27_47#_c_737_n 0.00374999f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B2_c_109_n N_A_27_47#_c_718_n 5.13362e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B2_c_110_n N_A_27_47#_c_718_n 0.00748944f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B2_c_111_n N_A_27_47#_c_718_n 0.0137981f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_163 N_B2_c_108_n N_A_27_47#_c_720_n 0.00116636f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B2_c_109_n N_A_27_47#_c_720_n 0.00116636f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_165 N_B2_c_111_n N_A_27_47#_c_720_n 0.0306016f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_166 N_B2_c_112_n N_A_27_47#_c_720_n 0.00358305f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_167 N_B2_c_107_n N_VGND_c_786_n 0.00379224f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_168 N_B2_c_108_n N_VGND_c_786_n 0.00276126f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B2_c_108_n N_VGND_c_787_n 0.00423334f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B2_c_109_n N_VGND_c_787_n 0.00423334f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B2_c_109_n N_VGND_c_788_n 0.00385467f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B2_c_110_n N_VGND_c_788_n 0.00365101f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B2_c_110_n N_VGND_c_791_n 0.00395087f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B2_c_107_n N_VGND_c_796_n 0.00692024f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B2_c_108_n N_VGND_c_796_n 0.00597024f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B2_c_109_n N_VGND_c_796_n 0.00620835f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B2_c_110_n N_VGND_c_796_n 0.0058395f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B2_c_107_n N_VGND_c_797_n 0.00423334f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B1_c_194_n N_A1_c_264_n 2.11242e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_180 N_B1_c_195_n N_A1_c_264_n 0.0138294f $X=3.845 $Y=1.16 $X2=0 $Y2=0
cc_181 N_B1_c_194_n N_A1_c_265_n 0.00655684f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_182 N_B1_c_195_n N_A1_c_265_n 9.97586e-19 $X=3.845 $Y=1.16 $X2=0 $Y2=0
cc_183 N_B1_c_196_n N_A_27_297#_c_417_n 0.0115796f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_184 N_B1_c_197_n N_A_27_297#_c_417_n 0.01161f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B1_c_198_n N_A_27_297#_c_419_n 0.01161f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B1_c_199_n N_A_27_297#_c_419_n 0.0143578f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_187 N_B1_c_199_n N_A_27_297#_c_399_n 7.75197e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B1_c_194_n N_A_27_297#_c_399_n 0.00406365f $X=3.785 $Y=1.202 $X2=0
+ $Y2=0
cc_189 N_B1_c_195_n N_A_27_297#_c_399_n 0.0440535f $X=3.845 $Y=1.16 $X2=0 $Y2=0
cc_190 N_B1_c_196_n N_Y_c_515_n 0.0119811f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B1_c_194_n N_Y_c_515_n 4.83683e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_192 N_B1_c_190_n N_Y_c_540_n 0.00292615f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_193 N_B1_c_190_n N_Y_c_513_n 0.00300439f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_194 N_B1_c_196_n N_Y_c_513_n 0.00104479f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_195 N_B1_c_191_n N_Y_c_513_n 0.00297134f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B1_c_197_n N_Y_c_513_n 9.09762e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B1_c_194_n N_Y_c_513_n 0.035936f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_198 N_B1_c_195_n N_Y_c_513_n 0.0156971f $X=3.845 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B1_c_191_n N_Y_c_514_n 0.0120408f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_200 N_B1_c_192_n N_Y_c_514_n 0.0107547f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B1_c_193_n N_Y_c_514_n 0.0133144f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B1_c_194_n N_Y_c_514_n 0.0124123f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_203 N_B1_c_195_n N_Y_c_514_n 0.0964685f $X=3.845 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B1_c_197_n N_Y_c_517_n 0.014627f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B1_c_198_n N_Y_c_517_n 0.0132328f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B1_c_194_n N_Y_c_517_n 0.00885447f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_207 N_B1_c_195_n N_Y_c_517_n 0.0397352f $X=3.845 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B1_c_196_n N_Y_c_520_n 0.0037472f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B1_c_194_n N_Y_c_520_n 0.00139638f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_210 N_B1_c_199_n N_Y_c_521_n 6.32035e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B1_c_194_n N_Y_c_521_n 0.00663436f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_212 N_B1_c_195_n N_Y_c_521_n 0.020385f $X=3.845 $Y=1.16 $X2=0 $Y2=0
cc_213 N_B1_c_196_n N_VPWR_c_617_n 0.00429453f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B1_c_197_n N_VPWR_c_617_n 0.00429453f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_215 N_B1_c_198_n N_VPWR_c_617_n 0.00429453f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B1_c_199_n N_VPWR_c_617_n 0.00429453f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_217 N_B1_c_196_n N_VPWR_c_612_n 0.00609021f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B1_c_197_n N_VPWR_c_612_n 0.00606499f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B1_c_198_n N_VPWR_c_612_n 0.00606499f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_220 N_B1_c_199_n N_VPWR_c_612_n 0.00734734f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_221 N_B1_c_190_n N_A_27_47#_c_719_n 0.0130858f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B1_c_191_n N_A_27_47#_c_719_n 0.00931157f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_223 N_B1_c_192_n N_A_27_47#_c_719_n 0.00931157f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B1_c_193_n N_A_27_47#_c_719_n 0.00931157f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_225 N_B1_c_194_n N_A_27_47#_c_719_n 4.78495e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_226 N_B1_c_190_n N_VGND_c_791_n 0.00357877f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_227 N_B1_c_191_n N_VGND_c_791_n 0.00357877f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B1_c_192_n N_VGND_c_791_n 0.00357877f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B1_c_193_n N_VGND_c_791_n 0.00357877f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B1_c_190_n N_VGND_c_796_n 0.00538422f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B1_c_191_n N_VGND_c_796_n 0.00548399f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B1_c_192_n N_VGND_c_796_n 0.00548399f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B1_c_193_n N_VGND_c_796_n 0.00668309f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A1_c_263_n N_A2_c_322_n 0.0175316f $X=6.21 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_235 N_A1_c_269_n N_A2_c_328_n 0.00985632f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A1_c_264_n N_A2_c_326_n 0.0150082f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A1_c_265_n N_A2_c_326_n 8.87282e-19 $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_238 N_A1_c_264_n N_A2_c_327_n 2.42383e-19 $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A1_c_265_n N_A2_c_327_n 0.0175316f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_240 N_A1_c_266_n N_A_27_297#_c_400_n 0.0159606f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A1_c_267_n N_A_27_297#_c_400_n 0.0156273f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A1_c_264_n N_A_27_297#_c_400_n 0.0480109f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A1_c_265_n N_A_27_297#_c_400_n 0.00837544f $X=6.185 $Y=1.202 $X2=0
+ $Y2=0
cc_244 N_A1_c_268_n N_A_27_297#_c_401_n 0.0156273f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A1_c_269_n N_A_27_297#_c_401_n 0.0156202f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A1_c_264_n N_A_27_297#_c_401_n 0.0480109f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A1_c_265_n N_A_27_297#_c_401_n 0.00816971f $X=6.185 $Y=1.202 $X2=0
+ $Y2=0
cc_248 N_A1_c_264_n N_A_27_297#_c_405_n 0.0204509f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A1_c_265_n N_A_27_297#_c_405_n 0.00656533f $X=6.185 $Y=1.202 $X2=0
+ $Y2=0
cc_250 N_A1_c_260_n N_Y_c_514_n 0.0133144f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A1_c_261_n N_Y_c_514_n 0.0107547f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A1_c_262_n N_Y_c_514_n 0.0107547f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A1_c_264_n N_Y_c_514_n 0.0842481f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A1_c_265_n N_Y_c_514_n 0.0115423f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_255 N_A1_c_266_n N_VPWR_c_613_n 0.00300743f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A1_c_267_n N_VPWR_c_613_n 0.00300743f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A1_c_268_n N_VPWR_c_614_n 0.00300743f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A1_c_269_n N_VPWR_c_614_n 0.00300743f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A1_c_266_n N_VPWR_c_617_n 0.00702461f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A1_c_267_n N_VPWR_c_619_n 0.00702461f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A1_c_268_n N_VPWR_c_619_n 0.00702461f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A1_c_269_n N_VPWR_c_621_n 0.00702461f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A1_c_266_n N_VPWR_c_612_n 0.0136915f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A1_c_267_n N_VPWR_c_612_n 0.0124092f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A1_c_268_n N_VPWR_c_612_n 0.0124092f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A1_c_269_n N_VPWR_c_612_n 0.0124344f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A1_c_260_n N_VGND_c_791_n 0.00357877f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A1_c_261_n N_VGND_c_791_n 0.00357877f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A1_c_262_n N_VGND_c_791_n 0.00357877f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A1_c_263_n N_VGND_c_791_n 0.00357877f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A1_c_260_n N_VGND_c_796_n 0.00668309f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A1_c_261_n N_VGND_c_796_n 0.00548399f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A1_c_262_n N_VGND_c_796_n 0.00560377f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A1_c_263_n N_VGND_c_796_n 0.005504f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A1_c_260_n N_A_883_47#_c_899_n 0.00931157f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A1_c_261_n N_A_883_47#_c_899_n 0.00931157f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A1_c_262_n N_A_883_47#_c_899_n 0.00964761f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A1_c_263_n N_A_883_47#_c_899_n 0.0117007f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A1_c_264_n N_A_883_47#_c_899_n 0.0039487f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A1_c_263_n N_A_883_47#_c_900_n 6.06509e-19 $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A2_c_328_n N_A_27_297#_c_402_n 0.0156202f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_282 N_A2_c_329_n N_A_27_297#_c_402_n 0.0156273f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_283 N_A2_c_326_n N_A_27_297#_c_402_n 0.0487385f $X=7.89 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A2_c_327_n N_A_27_297#_c_402_n 0.00837544f $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_285 N_A2_c_330_n N_A_27_297#_c_403_n 0.0156273f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_286 N_A2_c_331_n N_A_27_297#_c_403_n 0.0158328f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_287 N_A2_c_326_n N_A_27_297#_c_403_n 0.0487385f $X=7.89 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A2_c_327_n N_A_27_297#_c_403_n 0.00816971f $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_289 N_A2_c_326_n N_A_27_297#_c_404_n 0.0214236f $X=7.89 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A2_c_326_n N_A_27_297#_c_406_n 0.0029993f $X=7.89 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A2_c_326_n N_A_27_297#_c_407_n 0.0204509f $X=7.89 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A2_c_327_n N_A_27_297#_c_407_n 0.00656533f $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_293 N_A2_c_328_n N_VPWR_c_615_n 0.00300743f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_294 N_A2_c_329_n N_VPWR_c_615_n 0.00300743f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_295 N_A2_c_330_n N_VPWR_c_616_n 0.00300743f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_296 N_A2_c_331_n N_VPWR_c_616_n 0.00300743f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_297 N_A2_c_328_n N_VPWR_c_621_n 0.00702461f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_298 N_A2_c_329_n N_VPWR_c_623_n 0.00702461f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_299 N_A2_c_330_n N_VPWR_c_623_n 0.00702461f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_300 N_A2_c_331_n N_VPWR_c_625_n 0.00702461f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A2_c_328_n N_VPWR_c_612_n 0.0124344f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A2_c_329_n N_VPWR_c_612_n 0.0124092f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A2_c_330_n N_VPWR_c_612_n 0.0124092f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_304 N_A2_c_331_n N_VPWR_c_612_n 0.0134501f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A2_c_322_n N_VGND_c_789_n 0.00378935f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A2_c_323_n N_VGND_c_789_n 0.00276126f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A2_c_324_n N_VGND_c_790_n 0.00385467f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A2_c_325_n N_VGND_c_790_n 0.00365402f $X=8.09 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A2_c_322_n N_VGND_c_791_n 0.00421816f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A2_c_323_n N_VGND_c_793_n 0.00423334f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A2_c_324_n N_VGND_c_793_n 0.00423334f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A2_c_325_n N_VGND_c_795_n 0.00396605f $X=8.09 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A2_c_322_n N_VGND_c_796_n 0.00600232f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A2_c_323_n N_VGND_c_796_n 0.00597024f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A2_c_324_n N_VGND_c_796_n 0.00620835f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A2_c_325_n N_VGND_c_796_n 0.00689094f $X=8.09 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A2_c_322_n N_A_883_47#_c_911_n 0.00282739f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A2_c_322_n N_A_883_47#_c_900_n 0.00513906f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A2_c_323_n N_A_883_47#_c_900_n 4.74935e-19 $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A2_c_326_n N_A_883_47#_c_900_n 0.0061524f $X=7.89 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A2_c_322_n N_A_883_47#_c_901_n 0.00901745f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A2_c_323_n N_A_883_47#_c_901_n 0.00895898f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A2_c_326_n N_A_883_47#_c_901_n 0.0398926f $X=7.89 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A2_c_327_n N_A_883_47#_c_901_n 0.00345541f $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_325 N_A2_c_322_n N_A_883_47#_c_919_n 5.24597e-19 $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A2_c_323_n N_A_883_47#_c_919_n 0.00651696f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A2_c_324_n N_A_883_47#_c_919_n 0.00693563f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A2_c_325_n N_A_883_47#_c_919_n 5.34196e-19 $X=8.09 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A2_c_324_n N_A_883_47#_c_902_n 0.00929182f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A2_c_325_n N_A_883_47#_c_902_n 0.00936658f $X=8.09 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A2_c_326_n N_A_883_47#_c_902_n 0.071856f $X=7.89 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A2_c_327_n N_A_883_47#_c_902_n 0.00468948f $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_333 N_A2_c_324_n N_A_883_47#_c_903_n 5.69266e-19 $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A2_c_325_n N_A_883_47#_c_903_n 0.00857123f $X=8.09 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A2_c_323_n N_A_883_47#_c_904_n 0.00116636f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A2_c_324_n N_A_883_47#_c_904_n 0.00116636f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A2_c_326_n N_A_883_47#_c_904_n 0.0307014f $X=7.89 $Y=1.16 $X2=0 $Y2=0
cc_338 N_A2_c_327_n N_A_883_47#_c_904_n 0.00358305f $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_339 N_A_27_297#_c_413_n N_Y_M1002_s 0.00345323f $X=1.075 $Y=2.38 $X2=0 $Y2=0
cc_340 N_A_27_297#_c_415_n N_Y_M1021_s 0.00352392f $X=2.015 $Y=2.38 $X2=0 $Y2=0
cc_341 N_A_27_297#_c_417_n N_Y_M1000_s 0.00352392f $X=2.955 $Y=2.38 $X2=0 $Y2=0
cc_342 N_A_27_297#_c_419_n N_Y_M1009_s 0.00352392f $X=3.895 $Y=2.38 $X2=0 $Y2=0
cc_343 N_A_27_297#_M1028_d N_Y_c_515_n 0.00187422f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_344 N_A_27_297#_c_415_n N_Y_c_515_n 0.00387236f $X=2.015 $Y=2.38 $X2=0 $Y2=0
cc_345 N_A_27_297#_c_452_p N_Y_c_515_n 0.0143571f $X=2.14 $Y=1.96 $X2=0 $Y2=0
cc_346 N_A_27_297#_c_417_n N_Y_c_515_n 0.00235803f $X=2.955 $Y=2.38 $X2=0 $Y2=0
cc_347 N_A_27_297#_c_399_n N_Y_c_514_n 0.00728694f $X=4.28 $Y=1.625 $X2=0 $Y2=0
cc_348 N_A_27_297#_M1006_d N_Y_c_517_n 0.00187422f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_349 N_A_27_297#_c_417_n N_Y_c_517_n 0.00387236f $X=2.955 $Y=2.38 $X2=0 $Y2=0
cc_350 N_A_27_297#_c_457_p N_Y_c_517_n 0.0143571f $X=3.08 $Y=1.96 $X2=0 $Y2=0
cc_351 N_A_27_297#_c_419_n N_Y_c_517_n 0.00387236f $X=3.895 $Y=2.38 $X2=0 $Y2=0
cc_352 N_A_27_297#_M1013_d N_Y_c_518_n 0.00187422f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_353 N_A_27_297#_c_413_n N_Y_c_518_n 0.00387236f $X=1.075 $Y=2.38 $X2=0 $Y2=0
cc_354 N_A_27_297#_c_461_p N_Y_c_518_n 0.0143571f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_355 N_A_27_297#_c_415_n N_Y_c_518_n 0.00387236f $X=2.015 $Y=2.38 $X2=0 $Y2=0
cc_356 N_A_27_297#_c_415_n N_Y_c_519_n 0.0134104f $X=2.015 $Y=2.38 $X2=0 $Y2=0
cc_357 N_A_27_297#_c_417_n N_Y_c_520_n 0.0150725f $X=2.955 $Y=2.38 $X2=0 $Y2=0
cc_358 N_A_27_297#_c_419_n N_Y_c_521_n 0.0134104f $X=3.895 $Y=2.38 $X2=0 $Y2=0
cc_359 N_A_27_297#_c_399_n N_Y_c_521_n 0.00226124f $X=4.28 $Y=1.625 $X2=0 $Y2=0
cc_360 N_A_27_297#_c_398_n Y 0.0423323f $X=0.26 $Y=1.64 $X2=0 $Y2=0
cc_361 N_A_27_297#_c_413_n Y 0.0131056f $X=1.075 $Y=2.38 $X2=0 $Y2=0
cc_362 N_A_27_297#_c_400_n N_VPWR_M1004_d 0.00187091f $X=5.355 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_363 N_A_27_297#_c_401_n N_VPWR_M1019_d 0.00187091f $X=6.295 $Y=1.54 $X2=0
+ $Y2=0
cc_364 N_A_27_297#_c_402_n N_VPWR_M1011_d 0.00187091f $X=7.235 $Y=1.54 $X2=0
+ $Y2=0
cc_365 N_A_27_297#_c_403_n N_VPWR_M1022_d 0.00187091f $X=8.175 $Y=1.54 $X2=0
+ $Y2=0
cc_366 N_A_27_297#_c_400_n N_VPWR_c_613_n 0.0143191f $X=5.355 $Y=1.54 $X2=0
+ $Y2=0
cc_367 N_A_27_297#_c_401_n N_VPWR_c_614_n 0.0143191f $X=6.295 $Y=1.54 $X2=0
+ $Y2=0
cc_368 N_A_27_297#_c_402_n N_VPWR_c_615_n 0.0143191f $X=7.235 $Y=1.54 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_403_n N_VPWR_c_616_n 0.0143191f $X=8.175 $Y=1.54 $X2=0
+ $Y2=0
cc_370 N_A_27_297#_c_397_n N_VPWR_c_617_n 0.0215579f $X=0.257 $Y=2.295 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_413_n N_VPWR_c_617_n 0.0367458f $X=1.075 $Y=2.38 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_415_n N_VPWR_c_617_n 0.0386815f $X=2.015 $Y=2.38 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_417_n N_VPWR_c_617_n 0.0386815f $X=2.955 $Y=2.38 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_c_419_n N_VPWR_c_617_n 0.0386815f $X=3.895 $Y=2.38 $X2=0
+ $Y2=0
cc_375 N_A_27_297#_c_482_p N_VPWR_c_617_n 0.0515688f $X=4.28 $Y=2.295 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_c_483_p N_VPWR_c_617_n 0.0149886f $X=1.2 $Y=2.38 $X2=0 $Y2=0
cc_377 N_A_27_297#_c_484_p N_VPWR_c_617_n 0.0149886f $X=2.14 $Y=2.38 $X2=0 $Y2=0
cc_378 N_A_27_297#_c_485_p N_VPWR_c_617_n 0.0149886f $X=3.08 $Y=2.38 $X2=0 $Y2=0
cc_379 N_A_27_297#_c_486_p N_VPWR_c_619_n 0.0149311f $X=5.48 $Y=2.3 $X2=0 $Y2=0
cc_380 N_A_27_297#_c_487_p N_VPWR_c_621_n 0.0149311f $X=6.42 $Y=2.3 $X2=0 $Y2=0
cc_381 N_A_27_297#_c_488_p N_VPWR_c_623_n 0.0149311f $X=7.36 $Y=2.3 $X2=0 $Y2=0
cc_382 N_A_27_297#_c_489_p N_VPWR_c_625_n 0.0161853f $X=8.3 $Y=2.3 $X2=0 $Y2=0
cc_383 N_A_27_297#_M1002_d N_VPWR_c_612_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_M1013_d N_VPWR_c_612_n 0.00231264f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_385 N_A_27_297#_M1028_d N_VPWR_c_612_n 0.00231264f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_386 N_A_27_297#_M1006_d N_VPWR_c_612_n 0.00231264f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_M1016_d N_VPWR_c_612_n 0.00722341f $X=3.875 $Y=1.485 $X2=0
+ $Y2=0
cc_388 N_A_27_297#_M1007_s N_VPWR_c_612_n 0.00370124f $X=5.335 $Y=1.485 $X2=0
+ $Y2=0
cc_389 N_A_27_297#_M1029_s N_VPWR_c_612_n 0.00370124f $X=6.275 $Y=1.485 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_M1017_s N_VPWR_c_612_n 0.00370124f $X=7.215 $Y=1.485 $X2=0
+ $Y2=0
cc_391 N_A_27_297#_M1025_s N_VPWR_c_612_n 0.00462075f $X=8.155 $Y=1.485 $X2=0
+ $Y2=0
cc_392 N_A_27_297#_c_397_n N_VPWR_c_612_n 0.0127375f $X=0.257 $Y=2.295 $X2=0
+ $Y2=0
cc_393 N_A_27_297#_c_413_n N_VPWR_c_612_n 0.0225861f $X=1.075 $Y=2.38 $X2=0
+ $Y2=0
cc_394 N_A_27_297#_c_415_n N_VPWR_c_612_n 0.0239144f $X=2.015 $Y=2.38 $X2=0
+ $Y2=0
cc_395 N_A_27_297#_c_417_n N_VPWR_c_612_n 0.0239144f $X=2.955 $Y=2.38 $X2=0
+ $Y2=0
cc_396 N_A_27_297#_c_419_n N_VPWR_c_612_n 0.0239144f $X=3.895 $Y=2.38 $X2=0
+ $Y2=0
cc_397 N_A_27_297#_c_482_p N_VPWR_c_612_n 0.0296541f $X=4.28 $Y=2.295 $X2=0
+ $Y2=0
cc_398 N_A_27_297#_c_486_p N_VPWR_c_612_n 0.00955092f $X=5.48 $Y=2.3 $X2=0 $Y2=0
cc_399 N_A_27_297#_c_487_p N_VPWR_c_612_n 0.00955092f $X=6.42 $Y=2.3 $X2=0 $Y2=0
cc_400 N_A_27_297#_c_488_p N_VPWR_c_612_n 0.00955092f $X=7.36 $Y=2.3 $X2=0 $Y2=0
cc_401 N_A_27_297#_c_489_p N_VPWR_c_612_n 0.00955092f $X=8.3 $Y=2.3 $X2=0 $Y2=0
cc_402 N_A_27_297#_c_483_p N_VPWR_c_612_n 0.00962421f $X=1.2 $Y=2.38 $X2=0 $Y2=0
cc_403 N_A_27_297#_c_484_p N_VPWR_c_612_n 0.00962421f $X=2.14 $Y=2.38 $X2=0
+ $Y2=0
cc_404 N_A_27_297#_c_485_p N_VPWR_c_612_n 0.00962421f $X=3.08 $Y=2.38 $X2=0
+ $Y2=0
cc_405 N_A_27_297#_c_406_n N_A_883_47#_c_900_n 0.00719897f $X=6.42 $Y=1.62 $X2=0
+ $Y2=0
cc_406 N_Y_M1002_s N_VPWR_c_612_n 0.00232895f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_407 N_Y_M1021_s N_VPWR_c_612_n 0.00232895f $X=1.525 $Y=1.485 $X2=0 $Y2=0
cc_408 N_Y_M1000_s N_VPWR_c_612_n 0.00232895f $X=2.465 $Y=1.485 $X2=0 $Y2=0
cc_409 N_Y_M1009_s N_VPWR_c_612_n 0.00232895f $X=3.405 $Y=1.485 $X2=0 $Y2=0
cc_410 N_Y_c_514_n N_A_27_47#_M1018_d 0.00409698f $X=5.95 $Y=0.73 $X2=0 $Y2=0
cc_411 N_Y_c_514_n N_A_27_47#_M1027_d 0.00672859f $X=5.95 $Y=0.73 $X2=0 $Y2=0
cc_412 N_Y_c_515_n N_A_27_47#_c_718_n 0.00491589f $X=2.395 $Y=1.535 $X2=0 $Y2=0
cc_413 N_Y_c_513_n N_A_27_47#_c_718_n 0.00159171f $X=2.545 $Y=1.445 $X2=0 $Y2=0
cc_414 N_Y_M1015_s N_A_27_47#_c_719_n 0.00399909f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_415 N_Y_M1026_s N_A_27_47#_c_719_n 0.00400389f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_416 N_Y_c_540_n N_A_27_47#_c_719_n 0.0183182f $X=2.545 $Y=0.885 $X2=0 $Y2=0
cc_417 N_Y_c_514_n N_A_27_47#_c_719_n 0.08118f $X=5.95 $Y=0.73 $X2=0 $Y2=0
cc_418 N_Y_c_514_n N_VGND_c_791_n 0.00348529f $X=5.95 $Y=0.73 $X2=0 $Y2=0
cc_419 N_Y_M1015_s N_VGND_c_796_n 0.00256987f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_420 N_Y_M1026_s N_VGND_c_796_n 0.00256987f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_421 N_Y_M1005_s N_VGND_c_796_n 0.00256987f $X=4.825 $Y=0.235 $X2=0 $Y2=0
cc_422 N_Y_M1023_s N_VGND_c_796_n 0.00297142f $X=5.765 $Y=0.235 $X2=0 $Y2=0
cc_423 N_Y_c_514_n N_VGND_c_796_n 0.0116681f $X=5.95 $Y=0.73 $X2=0 $Y2=0
cc_424 N_Y_c_514_n N_A_883_47#_M1005_d 0.0069299f $X=5.95 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_425 N_Y_c_514_n N_A_883_47#_M1012_d 0.00406311f $X=5.95 $Y=0.73 $X2=0 $Y2=0
cc_426 N_Y_M1005_s N_A_883_47#_c_899_n 0.00400389f $X=4.825 $Y=0.235 $X2=0 $Y2=0
cc_427 N_Y_M1023_s N_A_883_47#_c_899_n 0.00507817f $X=5.765 $Y=0.235 $X2=0 $Y2=0
cc_428 N_Y_c_514_n N_A_883_47#_c_899_n 0.0960567f $X=5.95 $Y=0.73 $X2=0 $Y2=0
cc_429 N_A_27_47#_c_715_n N_VGND_M1008_d 0.00251047f $X=0.985 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_430 N_A_27_47#_c_717_n N_VGND_M1024_d 0.00348805f $X=1.925 $Y=0.815 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_c_714_n N_VGND_c_786_n 0.0181628f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_432 N_A_27_47#_c_715_n N_VGND_c_786_n 0.0127273f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_c_715_n N_VGND_c_787_n 0.00198695f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_729_n N_VGND_c_787_n 0.0223596f $X=1.2 $Y=0.39 $X2=0 $Y2=0
cc_435 N_A_27_47#_c_717_n N_VGND_c_787_n 0.00266636f $X=1.925 $Y=0.815 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_729_n N_VGND_c_788_n 0.0183628f $X=1.2 $Y=0.39 $X2=0 $Y2=0
cc_437 N_A_27_47#_c_717_n N_VGND_c_788_n 0.0131987f $X=1.925 $Y=0.815 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_c_737_n N_VGND_c_788_n 0.0172916f $X=2.075 $Y=0.475 $X2=0
+ $Y2=0
cc_439 N_A_27_47#_c_718_n N_VGND_c_788_n 0.00582645f $X=2.075 $Y=0.725 $X2=0
+ $Y2=0
cc_440 N_A_27_47#_c_717_n N_VGND_c_791_n 0.00199443f $X=1.925 $Y=0.815 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_c_737_n N_VGND_c_791_n 0.0186086f $X=2.075 $Y=0.475 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_719_n N_VGND_c_791_n 0.112077f $X=4.02 $Y=0.39 $X2=0 $Y2=0
cc_443 N_A_27_47#_M1008_s N_VGND_c_796_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_M1010_s N_VGND_c_796_n 0.0025535f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_M1030_s N_VGND_c_796_n 0.00215206f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_M1018_d N_VGND_c_796_n 0.00255381f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_M1027_d N_VGND_c_796_n 0.00250339f $X=3.835 $Y=0.235 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_714_n N_VGND_c_796_n 0.0124119f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_715_n N_VGND_c_796_n 0.00972452f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_729_n N_VGND_c_796_n 0.0141302f $X=1.2 $Y=0.39 $X2=0 $Y2=0
cc_451 N_A_27_47#_c_717_n N_VGND_c_796_n 0.0100158f $X=1.925 $Y=0.815 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_737_n N_VGND_c_796_n 0.0111017f $X=2.075 $Y=0.475 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_c_719_n N_VGND_c_796_n 0.0703895f $X=4.02 $Y=0.39 $X2=0 $Y2=0
cc_454 N_A_27_47#_c_714_n N_VGND_c_797_n 0.0209752f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_455 N_A_27_47#_c_715_n N_VGND_c_797_n 0.00266636f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_719_n N_A_883_47#_c_899_n 0.0188708f $X=4.02 $Y=0.39 $X2=0
+ $Y2=0
cc_457 N_VGND_c_796_n N_A_883_47#_M1005_d 0.00209344f $X=8.51 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_458 N_VGND_c_796_n N_A_883_47#_M1012_d 0.00255381f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_459 N_VGND_c_796_n N_A_883_47#_M1031_d 0.00215206f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_460 N_VGND_c_796_n N_A_883_47#_M1003_d 0.0025535f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_796_n N_A_883_47#_M1020_d 0.00209319f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_462 N_VGND_c_791_n N_A_883_47#_c_899_n 0.112077f $X=6.805 $Y=0 $X2=0 $Y2=0
cc_463 N_VGND_c_796_n N_A_883_47#_c_899_n 0.0703895f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_464 N_VGND_c_789_n N_A_883_47#_c_911_n 0.0141571f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_465 N_VGND_c_791_n N_A_883_47#_c_911_n 0.0152108f $X=6.805 $Y=0 $X2=0 $Y2=0
cc_466 N_VGND_c_796_n N_A_883_47#_c_911_n 0.00940698f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_467 N_VGND_c_789_n N_A_883_47#_c_900_n 0.00471242f $X=6.89 $Y=0.39 $X2=0
+ $Y2=0
cc_468 N_VGND_M1001_s N_A_883_47#_c_901_n 0.00251047f $X=6.705 $Y=0.235 $X2=0
+ $Y2=0
cc_469 N_VGND_c_789_n N_A_883_47#_c_901_n 0.0127273f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_470 N_VGND_c_791_n N_A_883_47#_c_901_n 0.00266636f $X=6.805 $Y=0 $X2=0 $Y2=0
cc_471 N_VGND_c_793_n N_A_883_47#_c_901_n 0.00198695f $X=7.745 $Y=0 $X2=0 $Y2=0
cc_472 N_VGND_c_796_n N_A_883_47#_c_901_n 0.00972452f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_790_n N_A_883_47#_c_919_n 0.0183628f $X=7.83 $Y=0.39 $X2=0 $Y2=0
cc_474 N_VGND_c_793_n N_A_883_47#_c_919_n 0.0223596f $X=7.745 $Y=0 $X2=0 $Y2=0
cc_475 N_VGND_c_796_n N_A_883_47#_c_919_n 0.0141302f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_476 N_VGND_M1014_s N_A_883_47#_c_902_n 0.00348805f $X=7.645 $Y=0.235 $X2=0
+ $Y2=0
cc_477 N_VGND_c_790_n N_A_883_47#_c_902_n 0.0131987f $X=7.83 $Y=0.39 $X2=0 $Y2=0
cc_478 N_VGND_c_793_n N_A_883_47#_c_902_n 0.00266636f $X=7.745 $Y=0 $X2=0 $Y2=0
cc_479 N_VGND_c_795_n N_A_883_47#_c_902_n 0.00199443f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_480 N_VGND_c_796_n N_A_883_47#_c_902_n 0.0100158f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_481 N_VGND_c_790_n N_A_883_47#_c_903_n 0.0223967f $X=7.83 $Y=0.39 $X2=0 $Y2=0
cc_482 N_VGND_c_795_n N_A_883_47#_c_903_n 0.024373f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_483 N_VGND_c_796_n N_A_883_47#_c_903_n 0.0141066f $X=8.51 $Y=0 $X2=0 $Y2=0
