* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_120_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=1.275e+12p ps=8.55e+06u
M1001 a_396_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=4.225e+11p pd=3.9e+06u as=3.8675e+11p ps=3.79e+06u
M1002 Y a_120_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.1e+11p pd=2.62e+06u as=0p ps=0u
M1003 VPWR B1 a_492_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 a_120_297# A2_N a_122_47# VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u
M1005 a_396_47# a_120_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1006 a_122_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_492_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A2_N a_120_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B2 a_396_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
